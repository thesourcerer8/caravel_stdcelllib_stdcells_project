VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ASYNC3
  CLASS CORE ;
  FOREIGN ASYNC3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 1.370 0.655 1.510 0.845 ;
        RECT 3.215 0.655 3.505 0.730 ;
        RECT 1.370 0.515 3.505 0.655 ;
        RECT 3.215 0.440 3.505 0.515 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.060 3.025 1.135 ;
        RECT 8.495 1.060 8.785 1.135 ;
        RECT 2.735 0.920 8.785 1.060 ;
        RECT 2.735 0.845 3.025 0.920 ;
        RECT 8.495 0.845 8.785 0.920 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.189000 ;
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 10.415 2.195 10.705 2.485 ;
        RECT 10.490 0.730 10.630 2.195 ;
        RECT 7.055 0.655 7.345 0.730 ;
        RECT 10.415 0.655 10.705 0.730 ;
        RECT 7.055 0.515 10.705 0.655 ;
        RECT 7.055 0.440 7.345 0.515 ;
        RECT 10.415 0.440 10.705 0.515 ;
    END
  END C
  PIN CN
    ANTENNAGATEAREA 0.189000 ;
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 1.775 1.995 2.065 2.070 ;
        RECT 9.935 1.995 10.225 2.070 ;
        RECT 1.775 1.855 10.225 1.995 ;
        RECT 1.775 1.780 2.065 1.855 ;
        RECT 9.935 1.780 10.225 1.855 ;
        RECT 10.010 1.135 10.150 1.780 ;
        RECT 9.935 0.845 10.225 1.135 ;
    END
  END CN
  PIN VGND
    ANTENNADIFFAREA 0.914200 ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 8.975 2.735 9.265 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.747200 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 11.520 3.415 ;
        RECT 0.155 3.090 11.365 3.245 ;
        RECT 4.635 2.715 4.965 3.090 ;
        RECT 8.955 2.715 9.285 3.090 ;
      LAYER mcon ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 9.035 2.795 9.205 2.965 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 11.520 3.330 ;
      LAYER li1 ;
        RECT 3.675 2.580 4.005 2.910 ;
        RECT 6.315 2.580 6.645 2.910 ;
        RECT 0.795 2.260 1.125 2.505 ;
        RECT 0.795 2.175 1.105 2.260 ;
        RECT 1.755 2.175 2.085 2.505 ;
        RECT 7.515 2.260 7.845 2.505 ;
        RECT 10.395 2.260 10.725 2.505 ;
        RECT 7.535 2.175 7.845 2.260 ;
        RECT 10.415 2.175 10.725 2.260 ;
        RECT 1.275 2.005 1.585 2.090 ;
        RECT 1.275 1.760 1.605 2.005 ;
        RECT 1.355 1.155 1.525 1.760 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 1.835 0.750 2.005 2.175 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 2.795 1.155 2.965 1.760 ;
        RECT 4.235 1.210 4.405 1.760 ;
        RECT 3.275 1.155 4.405 1.210 ;
        RECT 7.115 1.155 7.285 1.760 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 3.275 1.040 4.485 1.155 ;
        RECT 0.795 0.655 1.105 0.750 ;
        RECT 0.795 0.420 1.125 0.655 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.275 0.500 3.445 1.040 ;
        RECT 4.155 0.920 4.485 1.040 ;
        RECT 7.035 0.920 7.365 1.155 ;
        RECT 4.175 0.825 4.465 0.920 ;
        RECT 7.035 0.825 7.345 0.920 ;
        RECT 3.675 0.420 4.005 0.750 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 6.315 0.420 6.645 0.750 ;
        RECT 7.115 0.500 7.285 0.825 ;
        RECT 7.595 0.750 7.765 1.615 ;
        RECT 8.555 1.155 8.725 1.760 ;
        RECT 8.475 0.920 8.805 1.155 ;
        RECT 8.475 0.825 8.785 0.920 ;
        RECT 9.915 0.825 10.245 1.155 ;
        RECT 7.515 0.420 7.845 0.750 ;
        RECT 8.955 0.420 9.285 0.750 ;
        RECT 10.415 0.655 10.725 0.750 ;
        RECT 10.395 0.420 10.725 0.655 ;
        RECT 4.715 0.240 4.885 0.420 ;
        RECT 9.035 0.240 9.205 0.420 ;
        RECT 0.155 0.085 11.365 0.240 ;
        RECT 0.000 -0.085 11.520 0.085 ;
      LAYER mcon ;
        RECT 3.755 2.660 3.925 2.830 ;
        RECT 6.395 2.660 6.565 2.830 ;
        RECT 0.875 2.255 1.045 2.425 ;
        RECT 7.595 2.255 7.765 2.425 ;
        RECT 10.475 2.255 10.645 2.425 ;
        RECT 1.835 1.840 2.005 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 9.995 1.840 10.165 2.010 ;
        RECT 7.595 1.445 7.765 1.615 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 0.875 0.500 1.045 0.670 ;
        RECT 3.755 0.500 3.925 0.670 ;
        RECT 6.395 0.500 6.565 0.670 ;
        RECT 8.555 0.905 8.725 1.075 ;
        RECT 9.995 0.905 10.165 1.075 ;
        RECT 10.475 0.500 10.645 0.670 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
      LAYER met1 ;
        RECT 3.695 2.815 3.985 2.890 ;
        RECT 6.335 2.815 6.625 2.890 ;
        RECT 3.695 2.675 6.625 2.815 ;
        RECT 3.695 2.600 3.985 2.675 ;
        RECT 6.335 2.600 6.625 2.675 ;
        RECT 0.815 2.410 1.105 2.485 ;
        RECT 7.535 2.410 7.825 2.485 ;
        RECT 0.815 2.270 7.825 2.410 ;
        RECT 0.815 2.195 1.105 2.270 ;
        RECT 7.535 2.195 7.825 2.270 ;
        RECT 7.535 1.600 7.825 1.675 ;
        RECT 0.890 1.460 7.825 1.600 ;
        RECT 0.890 0.730 1.030 1.460 ;
        RECT 7.535 1.385 7.825 1.460 ;
        RECT 0.815 0.440 1.105 0.730 ;
        RECT 3.695 0.655 3.985 0.730 ;
        RECT 6.335 0.655 6.625 0.730 ;
        RECT 3.695 0.515 6.625 0.655 ;
        RECT 3.695 0.440 3.985 0.515 ;
        RECT 6.335 0.440 6.625 0.515 ;
  END
END ASYNC3
END LIBRARY

