magic
tech sky130A
magscale 1 2
timestamp 1624918199
<< obsli1 >>
rect 1152 2092 58848 57293
<< obsm1 >>
rect 16 1417 59888 57325
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< obsm2 >>
rect 22 59144 156 59200
rect 324 59144 636 59200
rect 804 59144 1116 59200
rect 1284 59144 1692 59200
rect 1860 59144 2172 59200
rect 2340 59144 2748 59200
rect 2916 59144 3228 59200
rect 3396 59144 3804 59200
rect 3972 59144 4284 59200
rect 4452 59144 4860 59200
rect 5028 59144 5340 59200
rect 5508 59144 5916 59200
rect 6084 59144 6396 59200
rect 6564 59144 6972 59200
rect 7140 59144 7452 59200
rect 7620 59144 8028 59200
rect 8196 59144 8508 59200
rect 8676 59144 9084 59200
rect 9252 59144 9564 59200
rect 9732 59144 10140 59200
rect 10308 59144 10620 59200
rect 10788 59144 11196 59200
rect 11364 59144 11676 59200
rect 11844 59144 12252 59200
rect 12420 59144 12732 59200
rect 12900 59144 13308 59200
rect 13476 59144 13788 59200
rect 13956 59144 14364 59200
rect 14532 59144 14844 59200
rect 15012 59144 15324 59200
rect 15492 59144 15900 59200
rect 16068 59144 16380 59200
rect 16548 59144 16956 59200
rect 17124 59144 17436 59200
rect 17604 59144 18012 59200
rect 18180 59144 18492 59200
rect 18660 59144 19068 59200
rect 19236 59144 19548 59200
rect 19716 59144 20124 59200
rect 20292 59144 20604 59200
rect 20772 59144 21180 59200
rect 21348 59144 21660 59200
rect 21828 59144 22236 59200
rect 22404 59144 22716 59200
rect 22884 59144 23292 59200
rect 23460 59144 23772 59200
rect 23940 59144 24348 59200
rect 24516 59144 24828 59200
rect 24996 59144 25404 59200
rect 25572 59144 25884 59200
rect 26052 59144 26460 59200
rect 26628 59144 26940 59200
rect 27108 59144 27516 59200
rect 27684 59144 27996 59200
rect 28164 59144 28572 59200
rect 28740 59144 29052 59200
rect 29220 59144 29628 59200
rect 29796 59144 30108 59200
rect 30276 59144 30588 59200
rect 30756 59144 31164 59200
rect 31332 59144 31644 59200
rect 31812 59144 32220 59200
rect 32388 59144 32700 59200
rect 32868 59144 33276 59200
rect 33444 59144 33756 59200
rect 33924 59144 34332 59200
rect 34500 59144 34812 59200
rect 34980 59144 35388 59200
rect 35556 59144 35868 59200
rect 36036 59144 36444 59200
rect 36612 59144 36924 59200
rect 37092 59144 37500 59200
rect 37668 59144 37980 59200
rect 38148 59144 38556 59200
rect 38724 59144 39036 59200
rect 39204 59144 39612 59200
rect 39780 59144 40092 59200
rect 40260 59144 40668 59200
rect 40836 59144 41148 59200
rect 41316 59144 41724 59200
rect 41892 59144 42204 59200
rect 42372 59144 42780 59200
rect 42948 59144 43260 59200
rect 43428 59144 43836 59200
rect 44004 59144 44316 59200
rect 44484 59144 44892 59200
rect 45060 59144 45372 59200
rect 45540 59144 45852 59200
rect 46020 59144 46428 59200
rect 46596 59144 46908 59200
rect 47076 59144 47484 59200
rect 47652 59144 47964 59200
rect 48132 59144 48540 59200
rect 48708 59144 49020 59200
rect 49188 59144 49596 59200
rect 49764 59144 50076 59200
rect 50244 59144 50652 59200
rect 50820 59144 51132 59200
rect 51300 59144 51708 59200
rect 51876 59144 52188 59200
rect 52356 59144 52764 59200
rect 52932 59144 53244 59200
rect 53412 59144 53820 59200
rect 53988 59144 54300 59200
rect 54468 59144 54876 59200
rect 55044 59144 55356 59200
rect 55524 59144 55932 59200
rect 56100 59144 56412 59200
rect 56580 59144 56988 59200
rect 57156 59144 57468 59200
rect 57636 59144 58044 59200
rect 58212 59144 58524 59200
rect 58692 59144 59100 59200
rect 59268 59144 59580 59200
rect 59748 59144 59882 59200
rect 22 856 59882 59144
rect 420 800 444 856
rect 900 800 924 856
rect 1284 800 1308 856
rect 1764 800 1788 856
rect 2244 800 2268 856
rect 2628 800 2652 856
rect 3108 800 3132 856
rect 3588 800 3612 856
rect 3972 800 3996 856
rect 4452 800 4476 856
rect 4836 800 4860 856
rect 5316 800 5340 856
rect 5796 800 5820 856
rect 6180 800 6204 856
rect 6660 800 6684 856
rect 7140 800 7164 856
rect 7524 800 7548 856
rect 8004 800 8028 856
rect 8388 800 8412 856
rect 8868 800 8892 856
rect 9348 800 9372 856
rect 9732 800 9756 856
rect 10212 800 10236 856
rect 10692 800 10716 856
rect 11076 800 11100 856
rect 11556 800 11580 856
rect 11940 800 11964 856
rect 12420 800 12444 856
rect 12900 800 12924 856
rect 13284 800 13308 856
rect 13764 800 13788 856
rect 14244 800 14268 856
rect 14628 800 14652 856
rect 15108 800 15132 856
rect 15588 800 15612 856
rect 15972 800 15996 856
rect 16452 800 16476 856
rect 16836 800 16860 856
rect 17316 800 17340 856
rect 17796 800 17820 856
rect 18180 800 18204 856
rect 18660 800 18684 856
rect 19140 800 19164 856
rect 19524 800 19548 856
rect 20004 800 20028 856
rect 20388 800 20412 856
rect 20868 800 20892 856
rect 21348 800 21372 856
rect 21732 800 21756 856
rect 22212 800 22236 856
rect 22692 800 22716 856
rect 23076 800 23100 856
rect 23556 800 23580 856
rect 23940 800 23964 856
rect 24420 800 24444 856
rect 24900 800 24924 856
rect 25284 800 25308 856
rect 25764 800 25788 856
rect 26244 800 26268 856
rect 26628 800 26652 856
rect 27108 800 27132 856
rect 27588 800 27612 856
rect 27972 800 27996 856
rect 28452 800 28476 856
rect 28836 800 28860 856
rect 29316 800 29340 856
rect 29796 800 29820 856
rect 30180 800 30204 856
rect 30660 800 30684 856
rect 31140 800 31164 856
rect 31524 800 31548 856
rect 32004 800 32028 856
rect 32388 800 32412 856
rect 32868 800 32892 856
rect 33348 800 33372 856
rect 33732 800 33756 856
rect 34212 800 34236 856
rect 34692 800 34716 856
rect 35076 800 35100 856
rect 35556 800 35580 856
rect 35940 800 35964 856
rect 36420 800 36444 856
rect 36900 800 36924 856
rect 37284 800 37308 856
rect 37764 800 37788 856
rect 38244 800 38268 856
rect 38628 800 38652 856
rect 39108 800 39132 856
rect 39588 800 39612 856
rect 39972 800 39996 856
rect 40452 800 40476 856
rect 40836 800 40860 856
rect 41316 800 41340 856
rect 41796 800 41820 856
rect 42180 800 42204 856
rect 42660 800 42684 856
rect 43140 800 43164 856
rect 43524 800 43548 856
rect 44004 800 44028 856
rect 44388 800 44412 856
rect 44868 800 44892 856
rect 45348 800 45372 856
rect 45732 800 45756 856
rect 46212 800 46236 856
rect 46692 800 46716 856
rect 47076 800 47100 856
rect 47556 800 47580 856
rect 47940 800 47964 856
rect 48420 800 48444 856
rect 48900 800 48924 856
rect 49284 800 49308 856
rect 49764 800 49788 856
rect 50244 800 50268 856
rect 50628 800 50652 856
rect 51108 800 51132 856
rect 51588 800 51612 856
rect 51972 800 51996 856
rect 52452 800 52476 856
rect 52836 800 52860 856
rect 53316 800 53340 856
rect 53796 800 53820 856
rect 54180 800 54204 856
rect 54660 800 54684 856
rect 55140 800 55164 856
rect 55524 800 55548 856
rect 56004 800 56028 856
rect 56388 800 56412 856
rect 56868 800 56892 856
rect 57348 800 57372 856
rect 57732 800 57756 856
rect 58212 800 58236 856
rect 58692 800 58716 856
rect 59076 800 59100 856
rect 59556 800 59580 856
<< obsm3 >>
rect 4256 2631 50656 57309
<< metal4 >>
rect 4256 2616 4576 57324
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 2616 19936 57324
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 2616 35296 57324
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 2616 50656 57324
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 13172 0 13228 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 499 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 500 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 501 nsew signal output
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 502 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 503 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 504 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 505 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 506 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 507 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 508 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 509 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 510 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 511 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 512 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 513 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 514 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 515 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 516 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 517 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 518 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 519 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 520 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 521 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 522 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 523 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 524 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 525 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 526 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 527 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 528 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 529 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 530 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 531 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 532 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 533 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 534 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 535 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 536 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 537 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 538 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 539 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 540 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 541 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 542 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 543 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 544 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 545 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 546 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 547 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 548 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 549 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 550 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 551 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 552 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 553 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 554 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 555 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 556 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 557 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 558 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 559 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 560 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 561 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 562 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 563 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 564 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 565 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 566 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 567 nsew signal output
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 568 nsew signal output
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 569 nsew signal output
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 570 nsew signal output
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 571 nsew signal output
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 572 nsew signal output
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 573 nsew signal output
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 574 nsew signal output
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 575 nsew signal output
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 576 nsew signal output
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 577 nsew signal output
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 578 nsew signal output
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 579 nsew signal output
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 580 nsew signal output
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 581 nsew signal output
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 582 nsew signal output
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 583 nsew signal output
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 584 nsew signal output
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 585 nsew signal output
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 586 nsew signal output
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 587 nsew signal output
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 588 nsew signal output
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 589 nsew signal output
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 590 nsew signal output
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 591 nsew signal output
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 592 nsew signal output
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 593 nsew signal output
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 594 nsew signal output
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 595 nsew signal output
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 596 nsew signal output
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 597 nsew signal output
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 598 nsew signal output
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 599 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 600 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 601 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 602 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 603 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 604 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 606 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 607 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 608 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 609 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 610 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 611 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 612 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 613 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 614 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 615 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 616 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 618 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 619 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 620 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 2177346
string GDS_START 251226
<< end >>

