VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 0.580 3.060 0.870 3.090 ;
        RECT 0.580 2.890 0.640 3.060 ;
        RECT 0.810 2.890 0.870 3.060 ;
        RECT 0.580 2.830 0.870 2.890 ;
        RECT 3.220 3.060 3.510 3.090 ;
        RECT 3.220 2.890 3.280 3.060 ;
        RECT 3.450 2.890 3.510 3.060 ;
        RECT 3.220 2.830 3.510 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.220 0.360 3.510 0.420 ;
        RECT 3.220 0.240 3.280 0.360 ;
        RECT 3.450 0.240 3.510 0.360 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.150 4.950 2.440 ;
        RECT 4.730 0.690 4.870 2.150 ;
        RECT 4.660 0.400 4.950 0.690 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.560 3.060 0.890 3.140 ;
        RECT 0.560 2.890 0.640 3.060 ;
        RECT 0.810 2.890 0.890 3.060 ;
        RECT 0.560 2.810 0.890 2.890 ;
        RECT 3.200 3.060 3.530 3.140 ;
        RECT 3.200 2.890 3.280 3.060 ;
        RECT 3.450 2.890 3.530 3.060 ;
        RECT 3.200 2.810 3.530 2.890 ;
        RECT 1.760 2.380 2.090 2.460 ;
        RECT 1.760 2.230 1.840 2.380 ;
        RECT 1.780 2.210 1.840 2.230 ;
        RECT 2.010 2.210 2.090 2.380 ;
        RECT 4.640 2.380 4.970 2.460 ;
        RECT 4.640 2.230 4.720 2.380 ;
        RECT 1.780 2.130 2.090 2.210 ;
        RECT 4.660 2.210 4.720 2.230 ;
        RECT 4.890 2.210 4.970 2.380 ;
        RECT 4.660 2.130 4.970 2.210 ;
        RECT 1.280 1.980 1.610 2.060 ;
        RECT 1.280 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 2.720 1.980 3.050 2.060 ;
        RECT 2.720 1.810 2.800 1.980 ;
        RECT 2.970 1.810 3.050 1.980 ;
        RECT 2.720 1.730 3.050 1.810 ;
        RECT 4.160 1.980 4.490 2.060 ;
        RECT 4.160 1.810 4.240 1.980 ;
        RECT 4.410 1.810 4.490 1.980 ;
        RECT 4.160 1.730 4.490 1.810 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.880 1.360 1.030 ;
        RECT 1.300 0.860 1.360 0.880 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.300 0.780 1.610 0.860 ;
        RECT 2.720 1.030 3.050 1.110 ;
        RECT 2.720 0.860 2.800 1.030 ;
        RECT 2.970 0.860 3.050 1.030 ;
        RECT 2.720 0.780 3.050 0.860 ;
        RECT 4.160 1.030 4.490 1.110 ;
        RECT 4.160 0.860 4.240 1.030 ;
        RECT 4.410 0.860 4.490 1.030 ;
        RECT 4.160 0.780 4.490 0.860 ;
        RECT 0.800 0.630 1.130 0.710 ;
        RECT 0.800 0.460 0.880 0.630 ;
        RECT 1.050 0.460 1.130 0.630 ;
        RECT 4.660 0.630 4.970 0.710 ;
        RECT 4.660 0.610 4.720 0.630 ;
        RECT 0.800 0.380 1.130 0.460 ;
        RECT 4.640 0.460 4.720 0.610 ;
        RECT 4.890 0.460 4.970 0.630 ;
        RECT 3.200 0.360 3.530 0.440 ;
        RECT 4.640 0.380 4.970 0.460 ;
        RECT 3.200 0.190 3.280 0.360 ;
        RECT 3.450 0.190 3.530 0.360 ;
        RECT 3.200 0.110 3.530 0.190 ;
      LAYER met1 ;
        RECT 1.780 2.380 2.070 2.440 ;
        RECT 1.780 2.370 1.840 2.380 ;
        RECT 0.890 2.230 1.840 2.370 ;
        RECT 0.890 0.690 1.030 2.230 ;
        RECT 1.780 2.210 1.840 2.230 ;
        RECT 2.010 2.370 2.070 2.380 ;
        RECT 2.010 2.230 4.390 2.370 ;
        RECT 2.010 2.210 2.070 2.230 ;
        RECT 1.780 2.150 2.070 2.210 ;
        RECT 4.250 2.040 4.390 2.230 ;
        RECT 4.180 1.980 4.470 2.040 ;
        RECT 4.180 1.810 4.240 1.980 ;
        RECT 4.410 1.810 4.470 1.980 ;
        RECT 4.180 1.750 4.470 1.810 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 4.180 1.030 4.470 1.090 ;
        RECT 4.180 0.860 4.240 1.030 ;
        RECT 4.410 0.860 4.470 1.030 ;
        RECT 4.180 0.800 4.470 0.860 ;
        RECT 0.820 0.630 1.110 0.690 ;
        RECT 0.820 0.460 0.880 0.630 ;
        RECT 1.050 0.460 1.110 0.630 ;
        RECT 0.820 0.400 1.110 0.460 ;
  END
END AND2X1
END LIBRARY

