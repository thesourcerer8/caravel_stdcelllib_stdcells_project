magic
tech sky130A
timestamp 1624066178
<< nwell >>
rect 0 179 720 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
<< ndiff >>
rect 82 67 111 73
rect 82 66 88 67
rect 58 50 88 66
rect 105 66 111 67
rect 370 67 399 73
rect 370 66 376 67
rect 105 50 137 66
rect 58 24 137 50
rect 152 49 281 66
rect 152 32 184 49
rect 201 32 281 49
rect 152 24 281 32
rect 296 50 376 66
rect 393 66 399 67
rect 610 67 639 73
rect 610 66 616 67
rect 393 50 425 66
rect 296 24 425 50
rect 440 49 569 66
rect 440 32 472 49
rect 489 32 569 49
rect 440 24 569 32
rect 584 50 616 66
rect 633 66 639 67
rect 633 50 663 66
rect 584 24 663 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 88 243
rect 105 226 137 243
rect 58 225 137 226
rect 152 301 281 309
rect 152 284 184 301
rect 201 284 281 301
rect 152 225 281 284
rect 296 243 425 309
rect 296 226 376 243
rect 393 226 425 243
rect 296 225 425 226
rect 440 301 569 309
rect 440 284 472 301
rect 489 284 569 301
rect 440 225 569 284
rect 584 243 663 309
rect 584 226 616 243
rect 633 226 663 243
rect 584 225 663 226
rect 82 220 111 225
rect 370 220 399 225
rect 610 220 639 225
<< ndiffc >>
rect 88 50 105 67
rect 184 32 201 49
rect 376 50 393 67
rect 472 32 489 49
rect 616 50 633 67
<< pdiffc >>
rect 88 226 105 243
rect 184 284 201 301
rect 376 226 393 243
rect 472 284 489 301
rect 616 226 633 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
<< locali >>
rect 176 301 209 309
rect 176 284 184 301
rect 201 284 209 301
rect 176 276 209 284
rect 464 301 497 309
rect 464 284 472 301
rect 489 284 497 301
rect 464 276 497 284
rect 80 243 113 251
rect 80 226 88 243
rect 105 226 113 243
rect 80 218 113 226
rect 368 243 401 251
rect 368 226 376 243
rect 393 226 401 243
rect 608 243 641 251
rect 608 226 616 243
rect 633 226 641 243
rect 368 218 399 226
rect 610 218 641 226
rect 130 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 416 108 449 116
rect 416 92 424 108
rect 272 83 305 91
rect 418 91 424 92
rect 441 91 449 108
rect 418 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 80 67 111 75
rect 80 50 88 67
rect 105 66 111 67
rect 368 67 401 75
rect 105 50 113 66
rect 80 42 113 50
rect 176 49 209 57
rect 176 32 184 49
rect 201 32 209 49
rect 368 50 376 67
rect 393 50 401 67
rect 610 67 641 75
rect 610 66 616 67
rect 368 42 401 50
rect 464 49 497 57
rect 176 27 209 32
rect 176 24 184 27
rect 201 24 209 27
rect 464 32 472 49
rect 489 32 497 49
rect 608 50 616 66
rect 633 50 641 67
rect 608 42 641 50
rect 464 27 497 32
rect 464 24 472 27
rect 489 24 497 27
<< viali >>
rect 184 284 201 301
rect 472 284 489 301
rect 88 226 105 243
rect 376 226 393 243
rect 616 226 633 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 88 50 105 67
rect 376 50 393 67
rect 184 10 201 27
rect 616 50 633 67
rect 472 10 489 27
<< metal1 >>
rect 0 309 720 357
rect 178 301 207 309
rect 178 284 184 301
rect 201 284 207 301
rect 178 278 207 284
rect 466 301 495 309
rect 466 284 472 301
rect 489 284 495 301
rect 466 278 495 284
rect 82 243 111 249
rect 82 226 88 243
rect 105 241 111 243
rect 370 243 399 249
rect 370 241 376 243
rect 105 227 376 241
rect 105 226 111 227
rect 82 220 111 226
rect 370 226 376 227
rect 393 241 399 243
rect 610 243 639 249
rect 610 241 616 243
rect 393 227 616 241
rect 393 226 399 227
rect 370 220 399 226
rect 610 226 616 227
rect 633 226 639 243
rect 610 220 639 226
rect 89 73 103 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 200 159 201
rect 274 201 303 207
rect 274 200 280 201
rect 153 186 280 200
rect 153 184 159 186
rect 130 178 159 184
rect 274 184 280 186
rect 297 200 303 201
rect 418 201 447 207
rect 418 200 424 201
rect 297 186 424 200
rect 297 184 303 186
rect 274 178 303 184
rect 418 184 424 186
rect 441 200 447 201
rect 562 201 591 207
rect 562 200 568 201
rect 441 186 568 200
rect 441 184 447 186
rect 418 178 447 184
rect 562 184 568 186
rect 585 184 591 201
rect 562 178 591 184
rect 137 114 151 178
rect 281 114 295 178
rect 425 114 439 178
rect 569 114 583 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 274 108 303 114
rect 274 91 280 108
rect 297 91 303 108
rect 274 85 303 91
rect 418 108 447 114
rect 418 91 424 108
rect 441 91 447 108
rect 418 85 447 91
rect 562 108 591 114
rect 562 91 568 108
rect 585 91 591 108
rect 562 85 591 91
rect 617 73 631 220
rect 82 67 111 73
rect 82 50 88 67
rect 105 50 111 67
rect 82 44 111 50
rect 370 67 399 73
rect 370 50 376 67
rect 393 66 399 67
rect 610 67 639 73
rect 610 66 616 67
rect 393 52 616 66
rect 393 50 399 52
rect 370 44 399 50
rect 610 50 616 52
rect 633 50 639 67
rect 610 44 639 50
rect 178 27 207 33
rect 178 24 184 27
rect 0 10 184 24
rect 201 24 207 27
rect 466 27 495 33
rect 466 24 472 27
rect 201 10 472 24
rect 489 24 495 27
rect 489 10 720 24
rect 0 -24 720 10
<< labels >>
rlabel metal1 0 309 720 357 0 VDD
port 1 se
rlabel metal1 0 -24 720 24 0 GND
port 2 se
rlabel metal1 370 44 399 52 0 Y
port 3 se
rlabel metal1 610 44 639 52 0 Y
port 4 se
rlabel metal1 370 52 639 66 0 Y
port 5 se
rlabel metal1 82 44 111 73 0 Y
port 6 se
rlabel metal1 370 66 399 73 0 Y
port 7 se
rlabel metal1 610 66 639 73 0 Y
port 8 se
rlabel metal1 89 73 103 220 0 Y
port 9 se
rlabel metal1 617 73 631 220 0 Y
port 10 se
rlabel metal1 82 220 111 227 0 Y
port 11 se
rlabel metal1 370 220 399 227 0 Y
port 12 se
rlabel metal1 610 220 639 227 0 Y
port 13 se
rlabel metal1 82 227 639 241 0 Y
port 14 se
rlabel metal1 82 241 111 249 0 Y
port 15 se
rlabel metal1 370 241 399 249 0 Y
port 16 se
rlabel metal1 610 241 639 249 0 Y
port 17 se
rlabel metal1 130 85 159 114 0 A
port 18 se
rlabel metal1 274 85 303 114 0 A
port 19 se
rlabel metal1 418 85 447 114 0 A
port 20 se
rlabel metal1 562 85 591 114 0 A
port 21 se
rlabel metal1 137 114 151 178 0 A
port 22 se
rlabel metal1 281 114 295 178 0 A
port 23 se
rlabel metal1 425 114 439 178 0 A
port 24 se
rlabel metal1 569 114 583 178 0 A
port 25 se
rlabel metal1 130 178 159 186 0 A
port 26 se
rlabel metal1 274 178 303 186 0 A
port 27 se
rlabel metal1 418 178 447 186 0 A
port 28 se
rlabel metal1 562 178 591 186 0 A
port 29 se
rlabel metal1 130 186 591 200 0 A
port 30 se
rlabel metal1 130 200 159 207 0 A
port 31 se
rlabel metal1 274 200 303 207 0 A
port 32 se
rlabel metal1 418 200 447 207 0 A
port 33 se
rlabel metal1 562 200 591 207 0 A
port 34 se
<< properties >>
string FIXED_BBOX 0 0 720 333
<< end >>
