magic
tech sky130A
magscale 1 2
timestamp 1636962374
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2592 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
rect 1713 48 1743 132
rect 2001 48 2031 132
rect 2289 48 2319 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
rect 1713 450 1743 618
rect 2001 450 2031 618
rect 2289 450 2319 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 355 134 413 146
rect 355 132 367 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 643 134 701 146
rect 643 132 655 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 100 655 132
rect 689 132 701 134
rect 931 134 989 146
rect 931 132 943 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 977 100 1137 132
rect 879 48 1137 100
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1507 134 1565 146
rect 1507 132 1519 134
rect 1265 100 1425 132
rect 1167 48 1425 100
rect 1455 100 1519 132
rect 1553 132 1565 134
rect 1795 134 1853 146
rect 1795 132 1807 134
rect 1553 100 1713 132
rect 1455 48 1713 100
rect 1743 100 1807 132
rect 1841 132 1853 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1841 100 2001 132
rect 1743 48 2001 100
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2371 134 2429 146
rect 2371 132 2383 134
rect 2129 100 2289 132
rect 2031 48 2289 100
rect 2319 100 2383 132
rect 2417 132 2429 134
rect 2417 100 2477 132
rect 2319 48 2477 100
<< pdiff >>
rect 115 593 273 618
rect 115 559 127 593
rect 161 559 273 593
rect 115 450 273 559
rect 303 485 561 618
rect 303 451 367 485
rect 401 451 561 485
rect 303 450 561 451
rect 591 593 849 618
rect 591 559 655 593
rect 689 559 849 593
rect 591 450 849 559
rect 879 485 1137 618
rect 879 451 943 485
rect 977 451 1137 485
rect 879 450 1137 451
rect 1167 593 1425 618
rect 1167 559 1231 593
rect 1265 559 1425 593
rect 1167 450 1425 559
rect 1455 485 1713 618
rect 1455 451 1519 485
rect 1553 451 1713 485
rect 1455 450 1713 451
rect 1743 593 2001 618
rect 1743 559 1807 593
rect 1841 559 2001 593
rect 1743 450 2001 559
rect 2031 485 2289 618
rect 2031 451 2095 485
rect 2129 451 2289 485
rect 2031 450 2289 451
rect 2319 593 2477 618
rect 2319 559 2383 593
rect 2417 559 2477 593
rect 2319 450 2477 559
rect 355 439 413 450
rect 931 439 989 450
rect 1507 439 1565 450
rect 2083 439 2141 450
<< ndiffc >>
rect 127 100 161 134
rect 367 100 401 134
rect 655 100 689 134
rect 943 100 977 134
rect 1231 100 1265 134
rect 1519 100 1553 134
rect 1807 100 1841 134
rect 2095 100 2129 134
rect 2383 100 2417 134
<< pdiffc >>
rect 127 559 161 593
rect 367 451 401 485
rect 655 559 689 593
rect 943 451 977 485
rect 1231 559 1265 593
rect 1519 451 1553 485
rect 1807 559 1841 593
rect 2095 451 2129 485
rect 2383 559 2417 593
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 2001 618 2031 644
rect 2289 618 2319 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 2001 418 2031 450
rect 2289 418 2319 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 181 2337 215
rect 2271 165 2337 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 2001 132 2031 165
rect 2289 132 2319 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
rect 1713 22 1743 48
rect 2001 22 2031 48
rect 2289 22 2319 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 2287 368 2321 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 2287 181 2321 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2592 683
rect 31 643 2561 649
rect 31 618 605 643
rect 739 618 2561 643
rect 111 593 177 618
rect 111 559 127 593
rect 161 559 177 593
rect 111 543 177 559
rect 639 593 705 609
rect 639 559 655 593
rect 689 559 705 593
rect 639 543 705 559
rect 1215 593 1281 618
rect 1215 559 1231 593
rect 1265 559 1281 593
rect 1215 543 1281 559
rect 1791 593 1857 618
rect 1791 559 1807 593
rect 1841 559 1857 593
rect 1791 543 1857 559
rect 2367 593 2433 618
rect 2367 559 2383 593
rect 2417 559 2433 593
rect 2367 543 2433 559
rect 351 485 417 501
rect 351 452 367 485
rect 355 451 367 452
rect 401 451 417 485
rect 355 435 417 451
rect 927 485 993 501
rect 927 451 943 485
rect 977 451 993 485
rect 1503 485 1569 501
rect 1503 452 1519 485
rect 927 435 993 451
rect 1507 451 1519 452
rect 1553 451 1569 485
rect 2079 485 2145 501
rect 2079 452 2095 485
rect 1507 435 1569 451
rect 2083 451 2095 452
rect 2129 451 2145 485
rect 2083 435 2145 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 893 418
rect 831 368 847 402
rect 881 401 893 402
rect 1119 402 1185 418
rect 881 368 897 401
rect 831 352 897 368
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 559 231 593 352
rect 1135 231 1169 352
rect 1711 231 1745 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 184 609 215
rect 831 215 897 231
rect 593 181 605 184
rect 543 165 605 181
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 184 1185 215
rect 1407 215 1473 231
rect 1169 181 1181 184
rect 1119 165 1181 181
rect 1407 181 1423 215
rect 1457 184 1473 215
rect 1695 215 1761 231
rect 1457 181 1469 184
rect 1407 165 1469 181
rect 1695 181 1711 215
rect 1745 184 1761 215
rect 1983 215 2049 231
rect 1745 181 1757 184
rect 1695 165 1757 181
rect 1983 181 1999 215
rect 2033 184 2049 215
rect 2033 181 2045 184
rect 1983 165 2045 181
rect 2095 150 2129 262
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 184 2337 215
rect 2321 181 2333 184
rect 2271 165 2333 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 355 134 417 150
rect 355 131 367 134
rect 111 84 177 100
rect 351 100 367 131
rect 401 100 417 134
rect 351 84 417 100
rect 639 134 705 150
rect 639 100 655 134
rect 689 100 705 134
rect 931 134 993 150
rect 931 131 943 134
rect 639 84 705 100
rect 927 100 943 131
rect 977 100 993 134
rect 927 84 993 100
rect 1215 134 1281 150
rect 1215 100 1231 134
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 1503 134 1569 150
rect 1503 100 1519 134
rect 1553 100 1569 134
rect 1503 84 1569 100
rect 1791 134 1857 150
rect 1791 100 1807 134
rect 1841 100 1857 134
rect 1791 84 1857 100
rect 2079 134 2145 150
rect 2079 100 2095 134
rect 2129 100 2145 134
rect 2079 84 2145 100
rect 2367 134 2433 150
rect 2367 100 2383 134
rect 2417 100 2433 134
rect 2367 84 2433 100
rect 31 17 2561 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2592 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 127 559 161 593
rect 655 559 689 593
rect 1231 559 1265 593
rect 1807 559 1841 593
rect 2383 559 2417 593
rect 367 451 401 485
rect 943 451 977 485
rect 1519 451 1553 485
rect 2095 451 2129 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 2287 368 2321 402
rect 2095 262 2129 296
rect 271 181 305 215
rect 847 181 881 215
rect 1423 181 1457 215
rect 1999 181 2033 215
rect 2287 181 2321 215
rect 127 100 161 134
rect 367 100 401 134
rect 655 100 689 134
rect 943 100 977 134
rect 1231 100 1265 134
rect 1519 100 1553 134
rect 1807 100 1841 134
rect 2383 100 2417 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2592 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2592 683
rect 0 618 2592 649
rect 115 593 173 618
rect 115 559 127 593
rect 161 559 173 593
rect 643 593 701 618
rect 115 547 173 559
rect 274 535 590 563
rect 643 559 655 593
rect 689 559 701 593
rect 1219 593 1277 618
rect 643 547 701 559
rect 274 414 302 535
rect 355 485 413 497
rect 355 451 367 485
rect 401 451 413 485
rect 355 439 413 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 274 227 302 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 370 212 398 439
rect 562 414 590 535
rect 850 535 1166 563
rect 1219 559 1231 593
rect 1265 559 1277 593
rect 1795 593 1853 618
rect 1219 547 1277 559
rect 850 414 878 535
rect 931 485 989 497
rect 931 451 943 485
rect 977 451 989 485
rect 931 439 989 451
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 850 227 878 356
rect 835 215 893 227
rect 835 212 847 215
rect 370 184 847 212
rect 370 146 398 184
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 946 212 974 439
rect 1138 414 1166 535
rect 1426 535 1742 563
rect 1795 559 1807 593
rect 1841 559 1853 593
rect 1795 547 1853 559
rect 2371 593 2429 618
rect 2371 559 2383 593
rect 2417 559 2429 593
rect 2371 547 2429 559
rect 1426 414 1454 535
rect 1507 485 1565 497
rect 1507 451 1519 485
rect 1553 451 1565 485
rect 1507 439 1565 451
rect 1123 402 1181 414
rect 1123 368 1135 402
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 1411 402 1469 414
rect 1411 368 1423 402
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1426 227 1454 356
rect 1411 215 1469 227
rect 1411 212 1423 215
rect 946 184 1423 212
rect 946 146 974 184
rect 1411 181 1423 184
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 1522 212 1550 439
rect 1714 414 1742 535
rect 2083 485 2141 497
rect 2083 451 2095 485
rect 2129 451 2141 485
rect 2083 439 2141 451
rect 1699 402 1757 414
rect 1699 368 1711 402
rect 1745 368 1757 402
rect 1699 356 1757 368
rect 1987 402 2045 414
rect 1987 368 1999 402
rect 2033 368 2045 402
rect 1987 356 2045 368
rect 2002 227 2030 356
rect 2098 308 2126 439
rect 2275 402 2333 414
rect 2275 368 2287 402
rect 2321 368 2333 402
rect 2275 356 2333 368
rect 2083 296 2141 308
rect 2083 262 2095 296
rect 2129 262 2141 296
rect 2083 250 2141 262
rect 2290 227 2318 356
rect 1987 215 2045 227
rect 1987 212 1999 215
rect 1522 184 1999 212
rect 1522 146 1550 184
rect 1987 181 1999 184
rect 2033 212 2045 215
rect 2275 215 2333 227
rect 2275 212 2287 215
rect 2033 184 2287 212
rect 2033 181 2045 184
rect 1987 169 2045 181
rect 2275 181 2287 184
rect 2321 181 2333 215
rect 2275 169 2333 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 355 134 413 146
rect 355 100 367 134
rect 401 100 413 134
rect 355 88 413 100
rect 643 134 701 146
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 931 134 989 146
rect 931 100 943 134
rect 977 100 989 134
rect 931 88 989 100
rect 1219 134 1277 146
rect 1219 100 1231 134
rect 1265 100 1277 134
rect 1219 88 1277 100
rect 1507 134 1565 146
rect 1507 100 1519 134
rect 1553 100 1565 134
rect 1507 88 1565 100
rect 1795 134 1853 146
rect 1795 100 1807 134
rect 1841 100 1853 134
rect 1795 88 1853 100
rect 2371 134 2429 146
rect 2371 100 2383 134
rect 2417 100 2429 134
rect 2371 88 2429 100
rect 130 48 158 88
rect 658 48 686 88
rect 1234 48 1262 88
rect 1810 48 1838 88
rect 2386 48 2414 88
rect 0 17 2592 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2592 17
rect 0 -48 2592 -17
<< labels >>
rlabel metal1 0 618 2592 714 0 VPWR
port 2 se
rlabel metal1 0 618 2592 714 0 VPWR
port 2 se
rlabel metal1 0 -48 2592 48 0 VGND
port 1 se
rlabel metal1 0 -48 2592 48 0 VGND
port 1 se
rlabel metal1 2083 250 2141 308 0 Y
port 3 se
rlabel metal1 2098 308 2126 439 0 Y
port 3 se
rlabel metal1 2083 439 2141 497 0 Y
port 3 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel metal1 547 356 605 414 0 A
port 0 se
rlabel metal1 274 414 302 535 0 A
port 0 se
rlabel metal1 562 414 590 535 0 A
port 0 se
rlabel metal1 274 535 590 563 0 A
port 0 se
rlabel locali 0 -17 2592 17 4 VGND
port 1 se ground default abutment
rlabel locali 31 17 2561 48 4 VGND
port 1 se ground default abutment
rlabel locali 0 649 2592 683 4 VPWR
port 2 se power default abutment
rlabel metal1 31 618 2561 649 4 VGND
port 1 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2592 666
<< end >>
