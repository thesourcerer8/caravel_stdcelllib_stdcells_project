MACRO OR2X1
 CLASS CORE ;
 FOREIGN OR2X1 0 0 ;
 SIZE 5.76 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN vdd
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;
    END
  END vdd

  PIN gnd
   DIRECTION INOUT ;
   USE GROUND ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
    END
  END gnd

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 4.65500000 0.44000000 4.94500000 0.73000000 ;
        RECT 4.73000000 0.73000000 4.87000000 2.19500000 ;
        RECT 4.65500000 2.19500000 4.94500000 2.48500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
        RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
        RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
    END
  END B


  OBS
    LAYER locali ;
      RECT ( 0 3.42 ) ( 5.76 3.57 ) ;
      RECT ( 0 3.25 ) ( 0.16 3.42 ) ;
      RECT ( 0.33 3.25 ) ( 0.64 3.42 ) ;
      RECT ( 0.81 3.25 ) ( 1.12 3.42 ) ;
      RECT ( 1.29 3.25 ) ( 1.6 3.42 ) ;
      RECT ( 1.77 3.25 ) ( 2.08 3.42 ) ;
      RECT ( 2.25 3.25 ) ( 2.56 3.42 ) ;
      RECT ( 2.73 3.25 ) ( 3.04 3.42 ) ;
      RECT ( 3.21 3.25 ) ( 3.52 3.42 ) ;
      RECT ( 3.69 3.25 ) ( 4 3.42 ) ;
      RECT ( 4.17 3.25 ) ( 4.48 3.42 ) ;
      RECT ( 4.65 3.25 ) ( 4.96 3.42 ) ;
      RECT ( 5.13 3.25 ) ( 5.44 3.42 ) ;
      RECT ( 5.61 3.25 ) ( 5.76 3.42 ) ;
      RECT ( 0 3.09 ) ( 5.76 3.25 ) ;
      RECT ( 3.2 2.99 ) ( 3.53 3.09 ) ;
      RECT ( 3.2 2.82 ) ( 3.28 2.99 ) ;
      RECT ( 3.45 2.82 ) ( 3.53 2.99 ) ;
      RECT ( 3.2 2.74 ) ( 3.53 2.82 ) ;
      RECT ( 0.8 2.43 ) ( 1.13 2.51 ) ;
      RECT ( 0.8 2.26 ) ( 0.88 2.43 ) ;
      RECT ( 1.05 2.26 ) ( 1.13 2.43 ) ;
      RECT ( 4.64 2.43 ) ( 4.97 2.51 ) ;
      RECT ( 4.64 2.26 ) ( 4.72 2.43 ) ;
      RECT ( 4.89 2.26 ) ( 4.97 2.43 ) ;
      RECT ( 0.8 2.18 ) ( 1.11 2.26 ) ;
      RECT ( 4.64 2.18 ) ( 4.97 2.26 ) ;
      RECT ( 1.28 2.01 ) ( 1.61 2.09 ) ;
      RECT ( 1.28 1.84 ) ( 1.36 2.01 ) ;
      RECT ( 1.53 1.84 ) ( 1.61 2.01 ) ;
      RECT ( 1.28 1.76 ) ( 1.61 1.84 ) ;
      RECT ( 2.72 2.01 ) ( 3.05 2.09 ) ;
      RECT ( 2.72 1.84 ) ( 2.8 2.01 ) ;
      RECT ( 2.97 1.84 ) ( 3.05 2.01 ) ;
      RECT ( 2.72 1.76 ) ( 3.05 1.84 ) ;
      RECT ( 4.16 2.01 ) ( 4.47 2.09 ) ;
      RECT ( 4.16 1.84 ) ( 4.24 2.01 ) ;
      RECT ( 4.41 1.84 ) ( 4.49 2.01 ) ;
      RECT ( 4.16 1.76 ) ( 4.49 1.84 ) ;
      RECT ( 1.28 1.08 ) ( 1.61 1.16 ) ;
      RECT ( 1.28 0.91 ) ( 1.36 1.08 ) ;
      RECT ( 1.53 0.91 ) ( 1.61 1.08 ) ;
      RECT ( 2.72 1.08 ) ( 3.05 1.16 ) ;
      RECT ( 2.72 0.92 ) ( 2.8 1.08 ) ;
      RECT ( 1.28 0.83 ) ( 1.61 0.91 ) ;
      RECT ( 2.74 0.91 ) ( 2.8 0.92 ) ;
      RECT ( 2.97 0.91 ) ( 3.05 1.08 ) ;
      RECT ( 2.74 0.83 ) ( 3.05 0.91 ) ;
      RECT ( 4.16 1.08 ) ( 4.49 1.16 ) ;
      RECT ( 4.16 0.91 ) ( 4.24 1.08 ) ;
      RECT ( 4.41 0.92 ) ( 4.49 1.08 ) ;
      RECT ( 4.41 0.91 ) ( 4.47 0.92 ) ;
      RECT ( 4.16 0.83 ) ( 4.47 0.91 ) ;
      RECT ( 2.24 0.67 ) ( 2.57 0.75 ) ;
      RECT ( 0.56 0.51 ) ( 0.89 0.59 ) ;
      RECT ( 0.56 0.34 ) ( 0.64 0.51 ) ;
      RECT ( 0.81 0.34 ) ( 0.89 0.51 ) ;
      RECT ( 2.24 0.5 ) ( 2.32 0.67 ) ;
      RECT ( 2.49 0.5 ) ( 2.57 0.67 ) ;
      RECT ( 4.64 0.67 ) ( 4.97 0.75 ) ;
      RECT ( 2.24 0.42 ) ( 2.57 0.5 ) ;
      RECT ( 3.2 0.51 ) ( 3.53 0.59 ) ;
      RECT ( 0.56 0.26 ) ( 0.89 0.34 ) ;
      RECT ( 3.2 0.34 ) ( 3.28 0.51 ) ;
      RECT ( 3.45 0.34 ) ( 3.53 0.51 ) ;
      RECT ( 4.64 0.5 ) ( 4.72 0.67 ) ;
      RECT ( 4.89 0.5 ) ( 4.97 0.67 ) ;
      RECT ( 4.64 0.42 ) ( 4.97 0.5 ) ;
      RECT ( 3.2 0.24 ) ( 3.53 0.34 ) ;
      RECT ( 0 0.09 ) ( 0.39 0.24 ) ;
      RECT ( 1.06 0.09 ) ( 5.76 0.24 ) ;
      RECT ( 0 -0.09 ) ( 0.16 0.09 ) ;
      RECT ( 0.33 -0.09 ) ( 0.64 0.09 ) ;
      RECT ( 0.81 -0.09 ) ( 1.12 0.09 ) ;
      RECT ( 1.29 -0.09 ) ( 1.6 0.09 ) ;
      RECT ( 1.77 -0.09 ) ( 2.08 0.09 ) ;
      RECT ( 2.25 -0.09 ) ( 2.56 0.09 ) ;
      RECT ( 2.73 -0.09 ) ( 3.04 0.09 ) ;
      RECT ( 3.21 -0.09 ) ( 3.52 0.09 ) ;
      RECT ( 3.69 -0.09 ) ( 4 0.09 ) ;
      RECT ( 4.17 -0.09 ) ( 4.48 0.09 ) ;
      RECT ( 4.65 -0.09 ) ( 4.96 0.09 ) ;
      RECT ( 5.13 -0.09 ) ( 5.44 0.09 ) ;
      RECT ( 5.61 -0.09 ) ( 5.76 0.09 ) ;
      RECT ( 0 -0.24 ) ( 5.76 -0.09 ) ;
    LAYER metal1 ;
      RECT ( 0 3.42 ) ( 5.76 3.57 ) ;
      RECT ( 0 3.25 ) ( 0.16 3.42 ) ;
      RECT ( 0.33 3.25 ) ( 0.64 3.42 ) ;
      RECT ( 0.81 3.25 ) ( 1.12 3.42 ) ;
      RECT ( 1.29 3.25 ) ( 1.6 3.42 ) ;
      RECT ( 1.77 3.25 ) ( 2.08 3.42 ) ;
      RECT ( 2.25 3.25 ) ( 2.56 3.42 ) ;
      RECT ( 2.73 3.25 ) ( 3.04 3.42 ) ;
      RECT ( 3.21 3.25 ) ( 3.52 3.42 ) ;
      RECT ( 3.69 3.25 ) ( 4 3.42 ) ;
      RECT ( 4.17 3.25 ) ( 4.48 3.42 ) ;
      RECT ( 4.65 3.25 ) ( 4.96 3.42 ) ;
      RECT ( 5.13 3.25 ) ( 5.44 3.42 ) ;
      RECT ( 5.61 3.25 ) ( 5.76 3.42 ) ;
      RECT ( 0 2.99 ) ( 5.76 3.25 ) ;
      RECT ( 0 2.82 ) ( 3.28 2.99 ) ;
      RECT ( 3.45 2.82 ) ( 5.76 2.99 ) ;
      RECT ( 0 2.43 ) ( 5.76 2.82 ) ;
      RECT ( 0 2.26 ) ( 0.88 2.43 ) ;
      RECT ( 1.05 2.26 ) ( 4.72 2.43 ) ;
      RECT ( 4.89 2.26 ) ( 5.76 2.43 ) ;
      RECT ( 0 2.01 ) ( 5.76 2.26 ) ;
      RECT ( 0 1.84 ) ( 1.36 2.01 ) ;
      RECT ( 1.53 1.84 ) ( 2.8 2.01 ) ;
      RECT ( 2.97 1.84 ) ( 4.24 2.01 ) ;
      RECT ( 4.41 1.84 ) ( 5.76 2.01 ) ;
      RECT ( 0 1.08 ) ( 5.76 1.84 ) ;
      RECT ( 0 0.91 ) ( 1.36 1.08 ) ;
      RECT ( 1.53 0.91 ) ( 2.8 1.08 ) ;
      RECT ( 2.97 0.91 ) ( 4.24 1.08 ) ;
      RECT ( 4.41 0.91 ) ( 5.76 1.08 ) ;
      RECT ( 0 0.67 ) ( 5.76 0.91 ) ;
      RECT ( 0 0.51 ) ( 2.32 0.67 ) ;
      RECT ( 0 0.34 ) ( 0.64 0.51 ) ;
      RECT ( 0.81 0.5 ) ( 2.32 0.51 ) ;
      RECT ( 2.49 0.5 ) ( 4.72 0.67 ) ;
      RECT ( 4.89 0.5 ) ( 5.76 0.67 ) ;
      RECT ( 0.81 0.34 ) ( 5.76 0.5 ) ;
      RECT ( 0 0.09 ) ( 5.76 0.34 ) ;
      RECT ( 0 -0.09 ) ( 0.16 0.09 ) ;
      RECT ( 0.33 -0.09 ) ( 0.64 0.09 ) ;
      RECT ( 0.81 -0.09 ) ( 1.12 0.09 ) ;
      RECT ( 1.29 -0.09 ) ( 1.6 0.09 ) ;
      RECT ( 1.77 -0.09 ) ( 2.08 0.09 ) ;
      RECT ( 2.25 -0.09 ) ( 2.56 0.09 ) ;
      RECT ( 2.73 -0.09 ) ( 3.04 0.09 ) ;
      RECT ( 3.21 -0.09 ) ( 3.52 0.09 ) ;
      RECT ( 3.69 -0.09 ) ( 4 0.09 ) ;
      RECT ( 4.17 -0.09 ) ( 4.48 0.09 ) ;
      RECT ( 4.65 -0.09 ) ( 4.96 0.09 ) ;
      RECT ( 5.13 -0.09 ) ( 5.44 0.09 ) ;
      RECT ( 5.61 -0.09 ) ( 5.76 0.09 ) ;
      RECT ( 0 -0.24 ) ( 5.76 -0.09 ) ;

  end
END OR2X1
