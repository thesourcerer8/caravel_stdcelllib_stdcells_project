MACRO BUFX4
 CLASS CORE ;
 FOREIGN BUFX4 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.69500000 0.39500000 3.98500000 0.47000000 ;
        RECT 3.69500000 0.47000000 4.87000000 0.61000000 ;
        RECT 3.69500000 0.61000000 3.98500000 0.68500000 ;
        RECT 3.21500000 2.15000000 3.50500000 2.22500000 ;
        RECT 3.69500000 2.15000000 3.98500000 2.22500000 ;
        RECT 4.73000000 0.61000000 4.87000000 2.22500000 ;
        RECT 3.21500000 2.22500000 4.87000000 2.36500000 ;
        RECT 3.21500000 2.36500000 3.50500000 2.44000000 ;
        RECT 3.69500000 2.36500000 3.98500000 2.44000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.29500000 1.74500000 1.58500000 2.03500000 ;
    END
  END A


END BUFX4
