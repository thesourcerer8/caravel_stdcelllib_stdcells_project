VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.370 0.870 2.440 ;
        RECT 3.220 2.370 3.510 2.440 ;
        RECT 0.580 2.230 3.510 2.370 ;
        RECT 0.580 2.150 0.870 2.230 ;
        RECT 3.220 2.150 3.510 2.230 ;
        RECT 6.100 2.150 6.390 2.440 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 6.170 0.690 6.310 2.150 ;
        RECT 0.580 0.610 0.870 0.690 ;
        RECT 3.220 0.610 3.510 0.690 ;
        RECT 6.100 0.610 6.390 0.690 ;
        RECT 0.580 0.470 6.390 0.610 ;
        RECT 0.580 0.400 0.870 0.470 ;
        RECT 3.220 0.400 3.510 0.470 ;
        RECT 6.100 0.400 6.390 0.470 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.960 1.590 2.040 ;
        RECT 2.740 1.960 3.030 2.040 ;
        RECT 4.180 1.960 4.470 2.040 ;
        RECT 5.620 1.960 5.910 2.040 ;
        RECT 1.300 1.820 5.910 1.960 ;
        RECT 1.300 1.750 1.590 1.820 ;
        RECT 2.740 1.750 3.030 1.820 ;
        RECT 4.180 1.750 4.470 1.820 ;
        RECT 5.620 1.750 5.910 1.820 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 5.690 1.090 5.830 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
        RECT 2.740 0.800 3.030 1.090 ;
        RECT 4.180 0.800 4.470 1.090 ;
        RECT 5.620 0.800 5.910 1.090 ;
    END
  END A
END INVX8
END LIBRARY

