MACRO LOFTY
 CLASS CORE ;
 FOREIGN LOFTY 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 21.60000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 21.60000000 0.24000000 ;
    END
  END GND

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.01500000 0.39500000 2.30500000 0.68500000 ;
        RECT 2.09000000 0.68500000 2.23000000 2.28500000 ;
        RECT 2.01500000 2.28500000 2.54500000 2.57500000 ;
    END
  END Q

  PIN ASEL_P
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 5.61500000 0.80000000 5.90500000 1.09000000 ;
        RECT 5.69000000 1.09000000 5.83000000 1.74500000 ;
        RECT 5.61500000 1.74500000 5.90500000 2.03500000 ;
    END
  END ASEL_P

  PIN USEXOR_N
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 15.69500000 0.53000000 15.98500000 0.60500000 ;
        RECT 20.01500000 0.53000000 20.30500000 0.60500000 ;
        RECT 15.69500000 0.60500000 20.30500000 0.74500000 ;
        RECT 15.69500000 0.74500000 15.98500000 0.82000000 ;
        RECT 20.01500000 0.74500000 20.30500000 0.82000000 ;
    END
  END USEXOR_N

  PIN USEMUX_N
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.81500000 0.39500000 1.10500000 0.68500000 ;
        RECT 1.29500000 0.80000000 1.58500000 1.09000000 ;
        RECT 1.37000000 1.09000000 1.51000000 1.74500000 ;
        RECT 1.29500000 1.74500000 1.58500000 1.88000000 ;
        RECT 1.29500000 1.88000000 1.82500000 2.03500000 ;
        RECT 1.53500000 2.03500000 1.82500000 2.17000000 ;
        RECT 0.89000000 0.68500000 1.03000000 2.22500000 ;
        RECT 1.53500000 2.17000000 1.75000000 2.22500000 ;
        RECT 0.89000000 2.22500000 1.75000000 2.36500000 ;
    END
  END USEMUX_N

  PIN USEXOR_P
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 8.49500000 1.74500000 8.78500000 2.03500000 ;
       LAYER metal2 ;
        RECT 17.13500000 1.74500000 17.42500000 2.03500000 ;
    END
  END USEXOR_P

  PIN ASEL_N
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7.05500000 0.80000000 7.34500000 1.09000000 ;
        RECT 7.13000000 1.09000000 7.27000000 1.34000000 ;
        RECT 7.05500000 1.34000000 7.34500000 1.63000000 ;
    END
  END ASEL_N

  PIN BSEL_N
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 18.57500000 1.34000000 18.86500000 2.03500000 ;
    END
  END BSEL_N

  PIN BSEL_P
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 14.25500000 1.34000000 14.54500000 1.63000000 ;
    END
  END BSEL_P

  PIN MUXSEL_P
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 10.65500000 1.74500000 10.94500000 1.82000000 ;
        RECT 10.65500000 1.82000000 11.11000000 2.01500000 ;
        RECT 11.85500000 1.74500000 12.14500000 2.01500000 ;
        RECT 11.61500000 2.01500000 12.14500000 2.03500000 ;
        RECT 10.41500000 2.01500000 11.11000000 2.03500000 ;
        RECT 10.41500000 2.03500000 10.70500000 2.09000000 ;
        RECT 10.97000000 2.03500000 11.11000000 2.09000000 ;
        RECT 11.61500000 2.03500000 11.90500000 2.09000000 ;
        RECT 10.97000000 2.09000000 11.90500000 2.23000000 ;
        RECT 9.05000000 2.09000000 10.70500000 2.23000000 ;
        RECT 10.41500000 2.23000000 10.70500000 2.30500000 ;
        RECT 11.61500000 2.23000000 11.90500000 2.30500000 ;
        RECT 7.53500000 2.28500000 7.82500000 2.36000000 ;
        RECT 9.05000000 2.23000000 9.19000000 2.36000000 ;
        RECT 7.53500000 2.36000000 9.19000000 2.50000000 ;
        RECT 7.53500000 2.50000000 7.82500000 2.57500000 ;
    END
  END MUXSEL_P

  PIN USEMUX_P
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.73500000 0.80000000 3.02500000 1.09000000 ;
        RECT 3.21500000 1.20500000 3.50500000 1.49500000 ;
        RECT 2.81000000 1.09000000 2.95000000 1.74500000 ;
        RECT 2.73500000 1.74500000 3.02500000 1.88000000 ;
        RECT 2.49500000 1.88000000 3.02500000 2.03500000 ;
        RECT 2.49500000 2.03500000 2.78500000 2.17000000 ;
        RECT 2.57000000 2.17000000 2.78500000 2.22500000 ;
        RECT 3.29000000 1.49500000 3.43000000 2.22500000 ;
        RECT 2.57000000 2.22500000 3.43000000 2.36500000 ;
    END
  END USEMUX_P

  PIN MUXSEL_N
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 10.65500000 1.74500000 10.94500000 1.82000000 ;
        RECT 10.65500000 1.82000000 11.11000000 2.01500000 ;
        RECT 11.85500000 1.74500000 12.14500000 2.01500000 ;
        RECT 11.61500000 2.01500000 12.14500000 2.03500000 ;
        RECT 10.41500000 2.01500000 11.11000000 2.03500000 ;
        RECT 10.41500000 2.03500000 10.70500000 2.09000000 ;
        RECT 10.97000000 2.03500000 11.11000000 2.09000000 ;
        RECT 11.61500000 2.03500000 11.90500000 2.09000000 ;
        RECT 10.97000000 2.09000000 11.90500000 2.23000000 ;
        RECT 9.05000000 2.09000000 10.70500000 2.23000000 ;
        RECT 10.41500000 2.23000000 10.70500000 2.30500000 ;
        RECT 11.61500000 2.23000000 11.90500000 2.30500000 ;
        RECT 7.53500000 2.28500000 7.82500000 2.36000000 ;
        RECT 9.05000000 2.23000000 9.19000000 2.36000000 ;
        RECT 7.53500000 2.36000000 9.19000000 2.50000000 ;
        RECT 7.53500000 2.50000000 7.82500000 2.57500000 ;
    END
  END MUXSEL_N


END LOFTY
