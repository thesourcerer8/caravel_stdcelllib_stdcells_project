magic
tech sky130A
magscale 1 2
timestamp 1636809582
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1440 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 643 134 701 146
rect 643 132 655 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 48 561 132
rect 591 100 655 132
rect 689 132 701 134
rect 931 134 989 146
rect 931 132 943 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 977 100 1137 132
rect 879 48 1137 100
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1265 100 1325 132
rect 1167 48 1325 100
<< pdiff >>
rect 115 593 273 618
rect 115 559 127 593
rect 161 559 273 593
rect 115 450 273 559
rect 303 450 561 618
rect 591 485 849 618
rect 591 451 655 485
rect 689 451 849 485
rect 591 450 849 451
rect 879 593 1137 618
rect 879 559 943 593
rect 977 559 1137 593
rect 879 450 1137 559
rect 1167 485 1325 618
rect 1167 451 1231 485
rect 1265 451 1325 485
rect 1167 450 1325 451
rect 643 439 701 450
rect 1219 439 1277 450
<< ndiffc >>
rect 127 100 161 134
rect 655 100 689 134
rect 943 100 977 134
rect 1231 100 1265 134
<< pdiffc >>
rect 127 559 161 593
rect 655 451 689 485
rect 943 559 977 593
rect 1231 451 1265 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
<< locali >>
rect 0 649 943 683
rect 977 649 1440 683
rect 31 643 1409 649
rect 31 618 893 643
rect 1027 618 1409 643
rect 111 593 177 618
rect 111 559 127 593
rect 161 559 177 593
rect 111 543 177 559
rect 927 593 993 609
rect 927 559 943 593
rect 977 559 993 593
rect 927 543 993 559
rect 639 485 705 501
rect 639 452 655 485
rect 643 451 655 452
rect 689 451 705 485
rect 1215 485 1281 501
rect 1215 452 1231 485
rect 643 435 705 451
rect 1219 451 1231 452
rect 1265 451 1281 485
rect 1219 435 1281 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 847 231 881 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 184 609 215
rect 831 215 897 231
rect 593 181 605 184
rect 543 165 605 181
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 184 1185 215
rect 1169 181 1181 184
rect 1119 165 1181 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 639 134 705 150
rect 639 100 655 134
rect 689 100 705 134
rect 931 134 993 150
rect 931 131 943 134
rect 639 84 705 100
rect 927 100 943 131
rect 977 100 993 134
rect 927 84 993 100
rect 1215 134 1281 150
rect 1215 100 1231 134
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 943 48 977 84
rect 31 17 1409 48
rect 0 -17 943 17
rect 977 -17 1440 17
<< viali >>
rect 943 649 977 683
rect 127 559 161 593
rect 943 559 977 593
rect 655 451 689 485
rect 1231 451 1265 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 271 181 305 215
rect 559 181 593 215
rect 1135 181 1169 215
rect 127 100 161 134
rect 655 100 689 134
rect 1231 100 1265 134
rect 943 -17 977 17
<< metal1 >>
rect 0 683 1440 714
rect 0 649 943 683
rect 977 649 1440 683
rect 0 618 1440 649
rect 115 593 173 618
rect 115 559 127 593
rect 161 559 173 593
rect 115 547 173 559
rect 931 593 989 618
rect 931 559 943 593
rect 977 559 989 593
rect 931 547 989 559
rect 643 485 701 497
rect 643 451 655 485
rect 689 451 701 485
rect 1219 485 1277 497
rect 1219 482 1231 485
rect 643 439 701 451
rect 850 454 1231 482
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 274 227 302 356
rect 562 227 590 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 658 212 686 439
rect 850 414 878 454
rect 1219 451 1231 454
rect 1265 451 1277 485
rect 1219 439 1277 451
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 1123 402 1181 414
rect 1123 368 1135 402
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 1138 227 1166 356
rect 1123 215 1181 227
rect 1123 212 1135 215
rect 658 184 1135 212
rect 658 146 686 184
rect 1123 181 1135 184
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 1234 146 1262 439
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 643 134 701 146
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 1219 134 1277 146
rect 1219 100 1231 134
rect 1265 100 1277 134
rect 1219 88 1277 100
rect 130 48 158 88
rect 0 17 1440 48
rect 0 -17 943 17
rect 977 -17 1440 17
rect 0 -48 1440 -17
<< labels >>
rlabel metal1 0 618 1440 714 0 VPWR
port 5 se
rlabel metal1 0 618 1440 714 0 VPWR
port 5 se
rlabel metal1 0 -48 1440 48 0 VGND
port 4 se
rlabel metal1 0 -48 1440 48 0 VGND
port 4 se
rlabel metal1 1219 88 1277 146 0 C
port 2 se
rlabel metal1 835 356 893 414 0 C
port 2 se
rlabel metal1 1234 146 1262 439 0 C
port 2 se
rlabel metal1 850 414 878 454 0 C
port 2 se
rlabel metal1 1219 439 1277 454 0 C
port 2 se
rlabel metal1 850 454 1277 482 0 C
port 2 se
rlabel metal1 1219 482 1277 497 0 C
port 2 se
rlabel metal1 643 88 701 146 0 CN
port 3 se
rlabel metal1 658 146 686 184 0 CN
port 3 se
rlabel metal1 1123 169 1181 184 0 CN
port 3 se
rlabel metal1 658 184 1181 212 0 CN
port 3 se
rlabel metal1 1123 212 1181 227 0 CN
port 3 se
rlabel metal1 1138 227 1166 356 0 CN
port 3 se
rlabel metal1 1123 356 1181 414 0 CN
port 3 se
rlabel metal1 658 212 686 439 0 CN
port 3 se
rlabel metal1 643 439 701 497 0 CN
port 3 se
rlabel metal1 547 169 605 227 0 B
port 1 se
rlabel metal1 562 227 590 356 0 B
port 1 se
rlabel metal1 547 356 605 414 0 B
port 1 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel locali 0 -17 1440 17 4 VGND
port 4 se ground default abutment
rlabel locali 31 17 1409 48 4 VGND
port 4 se ground default abutment
rlabel locali 0 649 1440 683 4 VPWR
port 5 se power default abutment
rlabel metal1 31 618 1409 649 4 VGND
port 4 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1440 666
<< end >>
