VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.995 1.585 2.070 ;
        RECT 2.735 1.995 3.025 2.070 ;
        RECT 1.295 1.855 3.025 1.995 ;
        RECT 1.295 1.780 1.585 1.855 ;
        RECT 2.735 1.780 3.025 1.855 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 2.735 0.845 3.025 1.135 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 0.562100 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 1.775 2.735 2.065 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.155 3.090 4.165 3.245 ;
        RECT 1.755 2.715 2.085 3.090 ;
      LAYER mcon ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 1.835 2.795 2.005 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 2.063300 ;
    PORT
      LAYER met1 ;
        RECT 0.815 2.410 1.105 2.485 ;
        RECT 3.215 2.410 3.505 2.485 ;
        RECT 0.815 2.270 3.505 2.410 ;
        RECT 0.815 2.195 1.105 2.270 ;
        RECT 3.215 2.195 3.505 2.270 ;
        RECT 0.890 0.730 1.030 2.195 ;
        RECT 3.290 0.730 3.430 2.195 ;
        RECT 0.815 0.440 1.105 0.730 ;
        RECT 3.215 0.440 3.505 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 4.320 3.330 ;
      LAYER li1 ;
        RECT 0.795 2.260 1.125 2.505 ;
        RECT 0.795 2.175 1.105 2.260 ;
        RECT 3.195 2.175 3.525 2.505 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 2.005 3.025 2.090 ;
        RECT 2.715 1.760 3.045 2.005 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.295 0.825 1.605 0.920 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 2.715 0.825 3.025 0.920 ;
        RECT 0.795 0.420 1.125 0.750 ;
        RECT 1.775 0.655 2.085 0.750 ;
        RECT 1.755 0.420 2.085 0.655 ;
        RECT 3.195 0.420 3.525 0.750 ;
        RECT 0.155 0.085 4.165 0.240 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.875 2.255 1.045 2.425 ;
        RECT 3.275 2.255 3.445 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 0.875 0.500 1.045 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
  END
END INVX4
END LIBRARY

