MACRO CLKBUF1
 CLASS CORE ;
 FOREIGN CLKBUF1 0 0 ;
 SIZE 12.96 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 12.96000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 12.96000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 12.96000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 12.96000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 10.41500000 1.25000000 10.70500000 1.54000000 ;
        RECT 10.49000000 1.54000000 10.63000000 2.19500000 ;
        RECT 10.41500000 2.19500000 10.70500000 2.48500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
        RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
        RECT 1.37000000 2.07000000 1.51000000 2.67500000 ;
        RECT 2.81000000 2.07000000 2.95000000 2.67500000 ;
        RECT 1.37000000 2.67500000 2.95000000 2.81500000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 8.55500000 0.90500000 8.72500000 1.07500000 ;
     RECT 9.99500000 0.90500000 10.16500000 1.07500000 ;
     RECT 11.43500000 0.90500000 11.60500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 8.55500000 1.84000000 8.72500000 2.01000000 ;
     RECT 9.99500000 1.84000000 10.16500000 2.01000000 ;
     RECT 11.43500000 1.84000000 11.60500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 1.83500000 2.25500000 2.00500000 2.42500000 ;
     RECT 4.71500000 2.25500000 4.88500000 2.42500000 ;
     RECT 7.59500000 2.25500000 7.76500000 2.42500000 ;
     RECT 10.47500000 2.25500000 10.64500000 2.42500000 ;
     RECT 0.63500000 2.79500000 0.80500000 2.96500000 ;
     RECT 3.27500000 2.79500000 3.44500000 2.96500000 ;
     RECT 6.15500000 2.79500000 6.32500000 2.96500000 ;
     RECT 9.03500000 2.79500000 9.20500000 2.96500000 ;
     RECT 11.91500000 2.79500000 12.08500000 2.96500000 ;

    LAYER ndiffc ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 1.83500000 0.50000000 2.00500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;
     RECT 4.71500000 0.50000000 4.88500000 0.67000000 ;
     RECT 6.15500000 0.50000000 6.32500000 0.67000000 ;
     RECT 7.59500000 0.50000000 7.76500000 0.67000000 ;
     RECT 9.03500000 0.50000000 9.20500000 0.67000000 ;
     RECT 10.47500000 0.50000000 10.64500000 0.67000000 ;
     RECT 11.91500000 0.50000000 12.08500000 0.67000000 ;

    LAYER li1 ;
     RECT 0.00000000 -0.24000000 12.96000000 0.24000000 ;
     RECT 0.55500000 0.42000000 0.88500000 0.75000000 ;
     RECT 1.75500000 0.42000000 2.08500000 0.75000000 ;
     RECT 3.19500000 0.42000000 3.52500000 0.75000000 ;
     RECT 4.63500000 0.42000000 4.96500000 0.75000000 ;
     RECT 6.07500000 0.42000000 6.40500000 0.75000000 ;
     RECT 7.51500000 0.42000000 7.84500000 0.75000000 ;
     RECT 8.95500000 0.42000000 9.28500000 0.75000000 ;
     RECT 11.83500000 0.42000000 12.16500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 4.15500000 0.82500000 4.48500000 1.15500000 ;
     RECT 7.03500000 0.82500000 7.36500000 1.15500000 ;
     RECT 9.91500000 0.82500000 10.24500000 1.15500000 ;
     RECT 11.35500000 0.82500000 11.68500000 1.15500000 ;
     RECT 10.39500000 0.42000000 10.72500000 0.75000000 ;
     RECT 10.47500000 0.75000000 10.64500000 1.48000000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 2.79500000 1.15500000 2.96500000 1.76000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 4.15500000 1.76000000 4.48500000 2.09000000 ;
     RECT 5.59500000 0.82500000 5.92500000 1.15500000 ;
     RECT 5.67500000 1.15500000 5.84500000 1.76000000 ;
     RECT 5.59500000 1.76000000 5.92500000 2.09000000 ;
     RECT 7.03500000 1.76000000 7.36500000 2.09000000 ;
     RECT 8.47500000 0.82500000 8.80500000 1.15500000 ;
     RECT 8.55500000 1.15500000 8.72500000 1.76000000 ;
     RECT 8.47500000 1.76000000 8.80500000 2.09000000 ;
     RECT 9.91500000 1.76000000 10.24500000 2.09000000 ;
     RECT 11.35500000 1.76000000 11.68500000 2.09000000 ;
     RECT 1.75500000 2.17500000 2.08500000 2.50500000 ;
     RECT 4.63500000 2.17500000 4.96500000 2.50500000 ;
     RECT 7.51500000 2.17500000 7.84500000 2.50500000 ;
     RECT 10.39500000 2.17500000 10.72500000 2.50500000 ;
     RECT 0.55500000 2.71500000 0.88500000 3.04500000 ;
     RECT 3.19500000 2.71500000 3.52500000 3.04500000 ;
     RECT 6.07500000 2.71500000 6.40500000 3.04500000 ;
     RECT 8.95500000 2.71500000 9.28500000 3.04500000 ;
     RECT 11.83500000 2.71500000 12.16500000 3.04500000 ;
     RECT 0.00000000 3.09000000 12.96000000 3.57000000 ;

    LAYER viali ;
     RECT 6.15500000 -0.08500000 6.32500000 0.08500000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 1.83500000 0.50000000 2.00500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;
     RECT 4.71500000 0.50000000 4.88500000 0.67000000 ;
     RECT 6.15500000 0.50000000 6.32500000 0.67000000 ;
     RECT 7.59500000 0.50000000 7.76500000 0.67000000 ;
     RECT 9.03500000 0.50000000 9.20500000 0.67000000 ;
     RECT 11.91500000 0.50000000 12.08500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 9.99500000 0.90500000 10.16500000 1.07500000 ;
     RECT 11.43500000 0.90500000 11.60500000 1.07500000 ;
     RECT 10.47500000 1.31000000 10.64500000 1.48000000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 8.55500000 1.84000000 8.72500000 2.01000000 ;
     RECT 9.99500000 1.84000000 10.16500000 2.01000000 ;
     RECT 11.43500000 1.84000000 11.60500000 2.01000000 ;
     RECT 1.83500000 2.25500000 2.00500000 2.42500000 ;
     RECT 4.71500000 2.25500000 4.88500000 2.42500000 ;
     RECT 7.59500000 2.25500000 7.76500000 2.42500000 ;
     RECT 10.47500000 2.25500000 10.64500000 2.42500000 ;
     RECT 0.63500000 2.79500000 0.80500000 2.96500000 ;
     RECT 3.27500000 2.79500000 3.44500000 2.96500000 ;
     RECT 6.15500000 2.79500000 6.32500000 2.96500000 ;
     RECT 9.03500000 2.79500000 9.20500000 2.96500000 ;
     RECT 11.91500000 2.79500000 12.08500000 2.96500000 ;
     RECT 6.15500000 3.24500000 6.32500000 3.41500000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 12.96000000 0.24000000 ;
     RECT 0.65000000 0.24000000 0.79000000 0.44000000 ;
     RECT 3.29000000 0.24000000 3.43000000 0.44000000 ;
     RECT 6.17000000 0.24000000 6.31000000 0.44000000 ;
     RECT 9.05000000 0.24000000 9.19000000 0.44000000 ;
     RECT 11.93000000 0.24000000 12.07000000 0.44000000 ;
     RECT 0.57500000 0.44000000 0.86500000 0.73000000 ;
     RECT 3.21500000 0.44000000 3.50500000 0.73000000 ;
     RECT 6.09500000 0.44000000 6.38500000 0.73000000 ;
     RECT 8.97500000 0.44000000 9.26500000 0.73000000 ;
     RECT 11.85500000 0.44000000 12.14500000 0.73000000 ;
     RECT 7.53500000 0.44000000 7.82500000 0.73000000 ;
     RECT 7.61000000 0.73000000 7.75000000 0.92000000 ;
     RECT 9.93500000 0.84500000 10.22500000 0.92000000 ;
     RECT 11.37500000 0.84500000 11.66500000 0.92000000 ;
     RECT 7.61000000 0.92000000 11.66500000 1.06000000 ;
     RECT 9.93500000 1.06000000 10.22500000 1.13500000 ;
     RECT 11.37500000 1.06000000 11.66500000 1.13500000 ;
     RECT 10.01000000 1.13500000 10.15000000 1.78000000 ;
     RECT 11.45000000 1.13500000 11.59000000 1.78000000 ;
     RECT 9.93500000 1.78000000 10.22500000 2.07000000 ;
     RECT 11.37500000 1.78000000 11.66500000 2.07000000 ;
     RECT 7.61000000 1.06000000 7.75000000 2.19500000 ;
     RECT 7.53500000 2.19500000 7.82500000 2.48500000 ;
     RECT 10.41500000 1.25000000 10.70500000 1.54000000 ;
     RECT 10.49000000 1.54000000 10.63000000 2.19500000 ;
     RECT 10.41500000 2.19500000 10.70500000 2.48500000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
     RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
     RECT 1.37000000 2.07000000 1.51000000 2.67500000 ;
     RECT 2.81000000 2.07000000 2.95000000 2.67500000 ;
     RECT 1.37000000 2.67500000 2.95000000 2.81500000 ;
     RECT 1.77500000 0.44000000 2.06500000 0.73000000 ;
     RECT 1.85000000 0.73000000 1.99000000 0.92000000 ;
     RECT 4.17500000 0.84500000 4.46500000 0.92000000 ;
     RECT 1.85000000 0.92000000 4.46500000 1.06000000 ;
     RECT 4.17500000 1.06000000 4.46500000 1.13500000 ;
     RECT 4.25000000 1.13500000 4.39000000 1.78000000 ;
     RECT 4.17500000 1.78000000 4.46500000 2.07000000 ;
     RECT 5.61500000 1.78000000 5.90500000 2.07000000 ;
     RECT 1.85000000 1.06000000 1.99000000 2.19500000 ;
     RECT 1.77500000 2.19500000 2.06500000 2.48500000 ;
     RECT 4.25000000 2.07000000 4.39000000 2.67500000 ;
     RECT 5.69000000 2.07000000 5.83000000 2.67500000 ;
     RECT 4.25000000 2.67500000 5.83000000 2.81500000 ;
     RECT 4.65500000 0.44000000 4.94500000 0.73000000 ;
     RECT 4.73000000 0.73000000 4.87000000 0.92000000 ;
     RECT 7.05500000 0.84500000 7.34500000 0.92000000 ;
     RECT 4.73000000 0.92000000 7.34500000 1.06000000 ;
     RECT 7.05500000 1.06000000 7.34500000 1.13500000 ;
     RECT 7.13000000 1.13500000 7.27000000 1.78000000 ;
     RECT 7.05500000 1.78000000 7.34500000 2.07000000 ;
     RECT 8.49500000 1.78000000 8.78500000 2.07000000 ;
     RECT 4.73000000 1.06000000 4.87000000 2.19500000 ;
     RECT 4.65500000 2.19500000 4.94500000 2.48500000 ;
     RECT 7.13000000 2.07000000 7.27000000 2.67500000 ;
     RECT 8.57000000 2.07000000 8.71000000 2.67500000 ;
     RECT 7.13000000 2.67500000 8.71000000 2.81500000 ;
     RECT 0.57500000 2.73500000 0.86500000 3.09000000 ;
     RECT 3.21500000 2.73500000 3.50500000 3.09000000 ;
     RECT 6.09500000 2.73500000 6.38500000 3.09000000 ;
     RECT 8.97500000 2.73500000 9.26500000 3.09000000 ;
     RECT 11.85500000 2.73500000 12.14500000 3.09000000 ;
     RECT 0.00000000 3.09000000 12.96000000 3.57000000 ;

 END
END CLKBUF1
