magic
tech sky130A
magscale 1 2
timestamp 1624953866
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 864 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 643 134 701 146
rect 643 132 655 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 102 561 132
rect 303 68 367 102
rect 401 68 561 102
rect 303 48 561 68
rect 591 100 655 132
rect 689 132 701 134
rect 689 100 749 132
rect 591 48 749 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 598 561 618
rect 303 564 367 598
rect 401 564 561 598
rect 303 450 561 564
rect 591 485 749 618
rect 591 451 655 485
rect 689 451 749 485
rect 591 450 749 451
rect 115 439 173 450
rect 643 439 701 450
<< ndiffc >>
rect 127 100 161 134
rect 367 68 401 102
rect 655 100 689 134
<< pdiffc >>
rect 127 451 161 485
rect 367 564 401 598
rect 655 451 689 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 273 418 303 450
rect 561 418 591 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 273 132 303 165
rect 561 132 591 165
rect 273 22 303 48
rect 561 22 591 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 271 181 305 215
rect 559 181 593 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 31 618 833 649
rect 351 598 417 618
rect 351 564 367 598
rect 401 564 417 598
rect 351 548 417 564
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 639 485 705 501
rect 639 451 655 485
rect 689 451 705 485
rect 639 435 705 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 605 418
rect 543 368 559 402
rect 593 401 605 402
rect 593 368 609 401
rect 543 352 609 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 184 609 215
rect 593 181 605 184
rect 543 165 605 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 639 134 705 150
rect 111 84 177 100
rect 351 102 417 118
rect 351 68 367 102
rect 401 68 417 102
rect 639 100 655 134
rect 689 100 705 134
rect 639 84 705 100
rect 351 48 417 68
rect 31 17 833 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 367 564 401 598
rect 127 451 161 485
rect 655 451 689 485
rect 271 368 305 402
rect 559 368 593 402
rect 271 181 305 215
rect 559 181 593 215
rect 127 100 161 134
rect 367 68 401 102
rect 655 100 689 134
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 714
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 618 864 649
rect 355 598 413 618
rect 355 564 367 598
rect 401 564 413 598
rect 355 552 413 564
rect 115 485 173 497
rect 115 451 127 485
rect 161 482 173 485
rect 643 485 701 497
rect 643 482 655 485
rect 161 454 655 482
rect 161 451 173 454
rect 115 439 173 451
rect 643 451 655 454
rect 689 451 701 485
rect 643 439 701 451
rect 130 146 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 399 317 402
rect 547 402 605 414
rect 547 399 559 402
rect 305 371 559 399
rect 305 368 317 371
rect 259 356 317 368
rect 547 368 559 371
rect 593 368 605 402
rect 547 356 605 368
rect 274 227 302 356
rect 562 227 590 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 658 146 686 439
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 643 134 701 146
rect 115 88 173 100
rect 355 102 413 114
rect 355 68 367 102
rect 401 68 413 102
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 355 48 413 68
rect 0 17 864 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -48 864 -17
<< labels >>
rlabel metal1 0 618 864 714 0 VPWR
port 2 se
rlabel metal1 0 618 864 714 0 VPWR
port 2 se
rlabel metal1 0 -48 864 48 0 VGND
port 1 se
rlabel metal1 0 -48 864 48 0 VGND
port 1 se
rlabel metal1 115 88 173 146 0 Y
port 3 se
rlabel metal1 643 88 701 146 0 Y
port 3 se
rlabel metal1 130 146 158 439 0 Y
port 3 se
rlabel metal1 658 146 686 439 0 Y
port 3 se
rlabel metal1 115 439 173 454 0 Y
port 3 se
rlabel metal1 643 439 701 454 0 Y
port 3 se
rlabel metal1 115 454 701 482 0 Y
port 3 se
rlabel metal1 115 482 173 497 0 Y
port 3 se
rlabel metal1 643 482 701 497 0 Y
port 3 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 547 169 605 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 562 227 590 356 0 A
port 0 se
rlabel metal1 259 356 317 371 0 A
port 0 se
rlabel metal1 547 356 605 371 0 A
port 0 se
rlabel metal1 259 371 605 399 0 A
port 0 se
rlabel metal1 259 399 317 414 0 A
port 0 se
rlabel metal1 547 399 605 414 0 A
port 0 se
rlabel locali 0 -17 864 17 4 VGND
port 1 se ground default abutment
rlabel locali 31 17 833 48 4 VGND
port 1 se ground default abutment
rlabel locali 0 649 864 683 4 VPWR
port 2 se power default abutment
rlabel locali 31 618 833 649 4 VGND
port 1 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 864 666
<< end >>
