magic
tech sky130A
magscale 1 2
timestamp 1624887581
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1152 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 739 134 797 146
rect 739 132 751 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 102 561 132
rect 303 68 367 102
rect 401 68 561 102
rect 303 48 561 68
rect 591 100 751 132
rect 785 132 797 134
rect 785 100 849 132
rect 591 48 849 100
rect 879 102 1037 132
rect 879 68 943 102
rect 977 68 1037 102
rect 879 48 1037 68
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 598 561 618
rect 303 564 367 598
rect 401 564 561 598
rect 303 450 561 564
rect 591 485 849 618
rect 591 451 751 485
rect 785 451 849 485
rect 591 450 849 451
rect 879 598 1037 618
rect 879 564 943 598
rect 977 564 1037 598
rect 879 450 1037 564
rect 115 439 173 450
rect 739 439 797 450
<< ndiffc >>
rect 127 100 161 134
rect 367 68 401 102
rect 751 100 785 134
rect 943 68 977 102
<< pdiffc >>
rect 127 451 161 485
rect 367 564 401 598
rect 751 451 785 485
rect 943 564 977 598
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 31 618 1121 649
rect 351 598 417 618
rect 351 564 367 598
rect 401 564 417 598
rect 351 548 417 564
rect 927 598 993 618
rect 927 564 943 598
rect 977 564 993 598
rect 927 548 993 564
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 735 485 801 501
rect 735 451 751 485
rect 785 451 801 485
rect 735 435 801 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 835 402 897 418
rect 835 401 847 402
rect 543 352 609 368
rect 831 368 847 401
rect 881 368 897 402
rect 831 352 897 368
rect 271 231 305 262
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 831 215 897 231
rect 831 184 847 215
rect 543 165 609 181
rect 835 181 847 184
rect 881 181 897 215
rect 835 165 897 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 735 134 801 150
rect 111 84 177 100
rect 351 102 417 118
rect 351 68 367 102
rect 401 68 417 102
rect 735 100 751 134
rect 785 100 801 134
rect 735 84 801 100
rect 927 102 993 118
rect 351 48 417 68
rect 927 68 943 102
rect 977 68 993 102
rect 927 48 993 68
rect 31 17 1121 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 367 564 401 598
rect 943 564 977 598
rect 127 451 161 485
rect 751 451 785 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 271 262 305 296
rect 559 181 593 215
rect 847 181 881 215
rect 127 100 161 134
rect 367 68 401 102
rect 751 100 785 134
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 714
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 618 1152 649
rect 355 598 413 618
rect 355 564 367 598
rect 401 564 413 598
rect 355 552 413 564
rect 931 598 989 618
rect 931 564 943 598
rect 977 564 989 598
rect 931 552 989 564
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 115 439 173 451
rect 739 485 797 497
rect 739 451 751 485
rect 785 482 797 485
rect 785 454 974 482
rect 785 451 797 454
rect 739 439 797 451
rect 130 212 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 274 308 302 356
rect 259 296 317 308
rect 259 262 271 296
rect 305 262 317 296
rect 259 250 317 262
rect 562 227 590 356
rect 850 227 878 356
rect 547 215 605 227
rect 547 212 559 215
rect 130 184 559 212
rect 130 146 158 184
rect 547 181 559 184
rect 593 212 605 215
rect 835 215 893 227
rect 835 212 847 215
rect 593 184 847 212
rect 593 181 605 184
rect 547 169 605 181
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 739 134 797 146
rect 115 88 173 100
rect 355 102 413 114
rect 355 68 367 102
rect 401 68 413 102
rect 739 100 751 134
rect 785 131 797 134
rect 946 131 974 454
rect 785 103 974 131
rect 785 100 797 103
rect 739 88 797 100
rect 355 48 413 68
rect 0 17 1152 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -48 1152 -17
<< labels >>
rlabel metal1 0 618 1152 714 0 VDD
port 1 se
rlabel metal1 0 618 1152 714 0 VDD
port 2 se
rlabel metal1 0 -48 1152 48 0 GND
port 3 se
rlabel metal1 0 -48 1152 48 0 GND
port 4 se
rlabel metal1 739 88 797 103 0 Y
port 5 se
rlabel metal1 739 103 974 131 0 Y
port 6 se
rlabel metal1 739 131 797 146 0 Y
port 7 se
rlabel metal1 739 439 797 454 0 Y
port 8 se
rlabel metal1 946 131 974 454 0 Y
port 9 se
rlabel metal1 739 454 974 482 0 Y
port 10 se
rlabel metal1 739 482 797 497 0 Y
port 11 se
rlabel metal1 259 250 317 308 0 A
port 12 se
rlabel metal1 274 308 302 356 0 A
port 13 se
rlabel metal1 259 356 317 414 0 A
port 14 se
rlabel locali 0 -17 1152 17 4 GND
port 3 se
rlabel locali 31 17 1121 48 4 GND
port 3 se
rlabel locali 0 649 1152 683 4 VDD
port 1 se
rlabel locali 31 618 1121 649 4 VDD
port 1 se
<< properties >>
string FIXED_BBOX 0 0 1152 666
<< end >>
