VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.780 3.010 2.070 3.090 ;
        RECT 7.540 3.070 7.600 3.090 ;
        RECT 7.770 3.070 7.830 3.090 ;
        RECT 7.540 3.010 7.830 3.070 ;
        RECT 1.780 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.070 3.010 ;
        RECT 1.780 2.780 2.070 2.840 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.270 2.070 0.330 ;
        RECT 1.780 0.240 1.840 0.270 ;
        RECT 2.010 0.240 2.070 0.270 ;
        RECT 7.540 0.270 7.830 0.330 ;
        RECT 7.540 0.240 7.600 0.270 ;
        RECT 7.770 0.240 7.830 0.270 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.140 2.410 5.430 2.490 ;
        RECT 5.140 2.270 6.310 2.410 ;
        RECT 5.140 2.200 5.430 2.270 ;
        RECT 5.140 0.660 5.430 0.730 ;
        RECT 6.170 0.660 6.310 2.270 ;
        RECT 5.140 0.520 6.310 0.660 ;
        RECT 5.140 0.440 5.430 0.520 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 5.620 2.000 5.910 2.070 ;
        RECT 4.250 1.860 5.910 2.000 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 4.250 1.140 4.390 1.860 ;
        RECT 5.620 1.780 5.910 1.860 ;
        RECT 1.300 1.060 1.590 1.140 ;
        RECT 4.180 1.060 4.470 1.140 ;
        RECT 1.300 0.920 4.470 1.060 ;
        RECT 1.300 0.850 1.590 0.920 ;
        RECT 4.180 0.850 4.470 0.920 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.810 2.680 8.710 2.820 ;
        RECT 2.810 2.070 2.950 2.680 ;
        RECT 8.570 2.070 8.710 2.680 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 8.500 1.780 8.790 2.070 ;
        RECT 8.570 1.140 8.710 1.780 ;
        RECT 8.500 0.850 8.790 1.140 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 1.760 3.010 2.090 3.090 ;
        RECT 1.760 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.090 3.010 ;
        RECT 1.760 2.760 2.090 2.840 ;
        RECT 7.520 3.070 7.600 3.090 ;
        RECT 7.770 3.070 7.850 3.090 ;
        RECT 7.520 3.010 7.850 3.070 ;
        RECT 7.520 2.840 7.600 3.010 ;
        RECT 7.770 2.840 7.850 3.010 ;
        RECT 7.520 2.760 7.850 2.840 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 5.120 2.430 5.450 2.510 ;
        RECT 5.120 2.260 5.200 2.430 ;
        RECT 5.370 2.260 5.450 2.430 ;
        RECT 8.960 2.430 9.290 2.510 ;
        RECT 8.960 2.260 9.040 2.430 ;
        RECT 9.210 2.260 9.290 2.430 ;
        RECT 5.120 2.180 5.430 2.260 ;
        RECT 8.980 2.180 9.290 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 3.450 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 2.800 1.160 2.970 1.760 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.920 5.680 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 5.620 0.910 5.680 0.920 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.620 0.830 5.930 0.910 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.370 1.080 ;
        RECT 7.040 0.830 7.370 0.910 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 8.480 0.910 8.560 1.080 ;
        RECT 8.730 0.910 8.810 1.080 ;
        RECT 8.480 0.830 8.810 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 5.120 0.670 5.450 0.750 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 1.760 0.490 2.090 0.570 ;
        RECT 1.760 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.090 0.490 ;
        RECT 5.120 0.500 5.200 0.670 ;
        RECT 5.370 0.500 5.450 0.670 ;
        RECT 8.980 0.670 9.290 0.750 ;
        RECT 8.980 0.660 9.040 0.670 ;
        RECT 5.120 0.420 5.450 0.500 ;
        RECT 7.520 0.490 7.850 0.570 ;
        RECT 1.760 0.270 2.090 0.320 ;
        RECT 1.760 0.240 1.840 0.270 ;
        RECT 2.010 0.240 2.090 0.270 ;
        RECT 7.520 0.320 7.600 0.490 ;
        RECT 7.770 0.320 7.850 0.490 ;
        RECT 8.960 0.500 9.040 0.660 ;
        RECT 9.210 0.500 9.290 0.670 ;
        RECT 8.960 0.420 9.290 0.500 ;
        RECT 7.520 0.270 7.850 0.320 ;
        RECT 7.520 0.240 7.600 0.270 ;
        RECT 7.770 0.240 7.850 0.270 ;
      LAYER met1 ;
        RECT 0.580 2.430 0.870 2.490 ;
        RECT 0.580 2.260 0.640 2.430 ;
        RECT 0.810 2.410 0.870 2.430 ;
        RECT 8.980 2.430 9.270 2.490 ;
        RECT 0.810 2.270 1.990 2.410 ;
        RECT 0.810 2.260 0.870 2.270 ;
        RECT 0.580 2.200 0.870 2.260 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 1.850 1.600 1.990 2.270 ;
        RECT 8.980 2.260 9.040 2.430 ;
        RECT 9.210 2.260 9.270 2.430 ;
        RECT 8.980 2.200 9.270 2.260 ;
        RECT 3.220 2.010 3.510 2.070 ;
        RECT 3.220 1.840 3.280 2.010 ;
        RECT 3.450 1.840 3.510 2.010 ;
        RECT 3.220 1.780 3.510 1.840 ;
        RECT 7.060 2.010 7.350 2.070 ;
        RECT 7.060 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.350 2.010 ;
        RECT 7.060 1.780 7.350 1.840 ;
        RECT 3.290 1.600 3.430 1.780 ;
        RECT 1.850 1.460 3.430 1.600 ;
        RECT 7.130 1.140 7.270 1.780 ;
        RECT 5.620 1.080 5.910 1.140 ;
        RECT 5.620 1.060 5.680 1.080 ;
        RECT 4.730 0.920 5.680 1.060 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.660 0.870 0.670 ;
        RECT 4.730 0.660 4.870 0.920 ;
        RECT 5.620 0.910 5.680 0.920 ;
        RECT 5.850 0.910 5.910 1.080 ;
        RECT 5.620 0.850 5.910 0.910 ;
        RECT 7.060 1.080 7.350 1.140 ;
        RECT 7.060 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.350 1.080 ;
        RECT 7.060 0.850 7.350 0.910 ;
        RECT 0.810 0.520 4.870 0.660 ;
        RECT 7.130 0.660 7.270 0.850 ;
        RECT 9.050 0.730 9.190 2.200 ;
        RECT 8.980 0.670 9.270 0.730 ;
        RECT 8.980 0.660 9.040 0.670 ;
        RECT 7.130 0.520 9.040 0.660 ;
        RECT 0.810 0.500 0.870 0.520 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 8.980 0.500 9.040 0.520 ;
        RECT 9.210 0.500 9.270 0.670 ;
        RECT 8.980 0.440 9.270 0.500 ;
  END
END XOR2X1
END LIBRARY

