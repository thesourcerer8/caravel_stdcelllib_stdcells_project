magic
tech sky130A
timestamp 1624702890
<< nwell >>
rect 0 179 1296 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
rect 857 24 872 66
rect 1001 24 1016 66
rect 1145 24 1160 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
rect 857 225 872 309
rect 1001 225 1016 309
rect 1145 225 1160 309
<< ndiff >>
rect 178 67 207 73
rect 178 66 184 67
rect 58 51 137 66
rect 58 34 64 51
rect 81 34 137 51
rect 58 24 137 34
rect 152 50 184 66
rect 201 66 207 67
rect 466 67 495 73
rect 466 66 472 67
rect 201 50 281 66
rect 152 24 281 50
rect 296 51 425 66
rect 296 34 328 51
rect 345 34 425 51
rect 296 24 425 34
rect 440 50 472 66
rect 489 66 495 67
rect 754 67 783 73
rect 754 66 760 67
rect 489 50 569 66
rect 440 24 569 50
rect 584 51 713 66
rect 584 34 616 51
rect 633 34 713 51
rect 584 24 713 34
rect 728 50 760 66
rect 777 66 783 67
rect 1042 67 1071 73
rect 1042 66 1048 67
rect 777 50 857 66
rect 728 24 857 50
rect 872 51 1001 66
rect 872 34 904 51
rect 921 34 1001 51
rect 872 24 1001 34
rect 1016 50 1048 66
rect 1065 66 1071 67
rect 1065 50 1145 66
rect 1016 24 1145 50
rect 1160 51 1239 66
rect 1160 34 1192 51
rect 1209 34 1239 51
rect 1160 24 1239 34
<< pdiff >>
rect 58 299 137 309
rect 58 282 64 299
rect 81 282 137 299
rect 58 225 137 282
rect 152 243 281 309
rect 152 226 184 243
rect 201 226 281 243
rect 152 225 281 226
rect 296 299 425 309
rect 296 282 328 299
rect 345 282 425 299
rect 296 225 425 282
rect 440 243 569 309
rect 440 226 472 243
rect 489 226 569 243
rect 440 225 569 226
rect 584 299 713 309
rect 584 282 616 299
rect 633 282 713 299
rect 584 225 713 282
rect 728 243 857 309
rect 728 226 760 243
rect 777 226 857 243
rect 728 225 857 226
rect 872 299 1001 309
rect 872 282 904 299
rect 921 282 1001 299
rect 872 225 1001 282
rect 1016 243 1145 309
rect 1016 226 1048 243
rect 1065 226 1145 243
rect 1016 225 1145 226
rect 1160 299 1239 309
rect 1160 282 1192 299
rect 1209 282 1239 299
rect 1160 225 1239 282
rect 178 220 207 225
rect 466 220 495 225
rect 754 220 783 225
rect 1042 220 1071 225
<< ndiffc >>
rect 64 34 81 51
rect 184 50 201 67
rect 328 34 345 51
rect 472 50 489 67
rect 616 34 633 51
rect 760 50 777 67
rect 904 34 921 51
rect 1048 50 1065 67
rect 1192 34 1209 51
<< pdiffc >>
rect 64 282 81 299
rect 184 226 201 243
rect 328 282 345 299
rect 472 226 489 243
rect 616 282 633 299
rect 760 226 777 243
rect 904 282 921 299
rect 1048 226 1065 243
rect 1192 282 1209 299
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 713 309 728 322
rect 857 309 872 322
rect 1001 309 1016 322
rect 1145 309 1160 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 713 209 728 225
rect 857 209 872 225
rect 1001 209 1016 225
rect 1145 209 1160 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 848 201 881 209
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 992 201 1025 209
rect 992 184 1000 201
rect 1017 184 1025 201
rect 992 176 1025 184
rect 1136 201 1169 209
rect 1136 184 1144 201
rect 1161 184 1169 201
rect 1136 176 1169 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 992 108 1025 116
rect 992 91 1000 108
rect 1017 91 1025 108
rect 992 83 1025 91
rect 1136 108 1169 116
rect 1136 91 1144 108
rect 1161 91 1169 108
rect 1136 83 1169 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 713 66 728 83
rect 857 66 872 83
rect 1001 66 1016 83
rect 1145 66 1160 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
rect 857 11 872 24
rect 1001 11 1016 24
rect 1145 11 1160 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 856 184 873 201
rect 1000 184 1017 201
rect 1144 184 1161 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
rect 856 91 873 108
rect 1000 91 1017 108
rect 1144 91 1161 108
<< locali >>
rect 0 342 1296 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 736 342
rect 753 325 784 342
rect 801 325 832 342
rect 849 325 880 342
rect 897 325 928 342
rect 945 325 976 342
rect 993 325 1024 342
rect 1041 325 1072 342
rect 1089 325 1120 342
rect 1137 325 1168 342
rect 1185 325 1216 342
rect 1233 325 1264 342
rect 1281 325 1296 342
rect 0 309 1296 325
rect 56 299 89 309
rect 56 282 64 299
rect 81 282 89 299
rect 56 274 89 282
rect 320 299 353 309
rect 320 282 328 299
rect 345 282 353 299
rect 320 274 353 282
rect 608 299 641 309
rect 608 282 616 299
rect 633 282 641 299
rect 608 274 641 282
rect 896 299 929 309
rect 896 282 904 299
rect 921 282 929 299
rect 896 274 929 282
rect 1184 299 1217 309
rect 1184 282 1192 299
rect 1209 282 1217 299
rect 1184 274 1217 282
rect 176 243 209 251
rect 176 226 184 243
rect 201 226 209 243
rect 464 243 497 251
rect 464 226 472 243
rect 489 226 497 243
rect 178 218 209 226
rect 466 218 497 226
rect 752 243 785 251
rect 752 226 760 243
rect 777 226 785 243
rect 1040 243 1073 251
rect 1040 226 1048 243
rect 1065 226 1073 243
rect 752 218 785 226
rect 1042 218 1073 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 735 209
rect 848 201 881 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 992 201 1025 209
rect 992 184 1000 201
rect 1017 184 1025 201
rect 992 176 1025 184
rect 1136 201 1169 209
rect 1136 184 1144 201
rect 1161 184 1169 201
rect 1136 176 1169 184
rect 280 116 297 176
rect 568 116 585 176
rect 856 116 873 176
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 92 449 108
rect 560 108 593 116
rect 441 91 447 92
rect 416 83 447 91
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 92 737 108
rect 848 108 881 116
rect 729 91 735 92
rect 704 83 735 91
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 992 108 1025 116
rect 992 91 1000 108
rect 1017 92 1025 108
rect 1017 91 1023 92
rect 992 83 1023 91
rect 1048 75 1065 131
rect 1136 108 1169 116
rect 1136 91 1144 108
rect 1161 91 1169 108
rect 1136 83 1169 91
rect 178 67 209 75
rect 178 66 184 67
rect 56 51 89 59
rect 56 34 64 51
rect 81 34 89 51
rect 176 50 184 66
rect 201 50 209 67
rect 464 67 497 75
rect 176 42 209 50
rect 320 51 353 59
rect 56 24 89 34
rect 320 34 328 51
rect 345 34 353 51
rect 464 50 472 67
rect 489 50 497 67
rect 752 67 785 75
rect 464 42 497 50
rect 608 51 641 59
rect 320 24 353 34
rect 608 34 616 51
rect 633 34 641 51
rect 752 50 760 67
rect 777 50 785 67
rect 1040 67 1073 75
rect 752 42 785 50
rect 896 51 929 59
rect 608 24 641 34
rect 896 34 904 51
rect 921 34 929 51
rect 1040 50 1048 67
rect 1065 50 1073 67
rect 1040 42 1073 50
rect 1184 51 1217 59
rect 896 24 929 34
rect 1184 34 1192 51
rect 1209 34 1217 51
rect 1184 24 1217 34
rect 0 9 1296 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 736 9
rect 753 -9 784 9
rect 801 -9 832 9
rect 849 -9 880 9
rect 897 -9 928 9
rect 945 -9 976 9
rect 993 -9 1024 9
rect 1041 -9 1072 9
rect 1089 -9 1120 9
rect 1137 -9 1168 9
rect 1185 -9 1216 9
rect 1233 -9 1264 9
rect 1281 -9 1296 9
rect 0 -24 1296 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 448 325 465 342
rect 496 325 513 342
rect 544 325 561 342
rect 592 325 609 342
rect 640 325 657 342
rect 688 325 705 342
rect 736 325 753 342
rect 784 325 801 342
rect 832 325 849 342
rect 880 325 897 342
rect 928 325 945 342
rect 976 325 993 342
rect 1024 325 1041 342
rect 1072 325 1089 342
rect 1120 325 1137 342
rect 1168 325 1185 342
rect 1216 325 1233 342
rect 1264 325 1281 342
rect 64 282 81 299
rect 328 282 345 299
rect 616 282 633 299
rect 904 282 921 299
rect 1192 282 1209 299
rect 184 226 201 243
rect 472 226 489 243
rect 760 226 777 243
rect 1048 226 1065 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 856 184 873 201
rect 1000 184 1017 201
rect 1144 184 1161 201
rect 1048 131 1065 148
rect 136 91 153 108
rect 424 91 441 108
rect 712 91 729 108
rect 1000 91 1017 108
rect 1144 91 1161 108
rect 64 34 81 51
rect 184 50 201 67
rect 328 34 345 51
rect 472 50 489 67
rect 616 34 633 51
rect 760 50 777 67
rect 904 34 921 51
rect 1192 34 1209 51
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
rect 448 -9 465 9
rect 496 -9 513 9
rect 544 -9 561 9
rect 592 -9 609 9
rect 640 -9 657 9
rect 688 -9 705 9
rect 736 -9 753 9
rect 784 -9 801 9
rect 832 -9 849 9
rect 880 -9 897 9
rect 928 -9 945 9
rect 976 -9 993 9
rect 1024 -9 1041 9
rect 1072 -9 1089 9
rect 1120 -9 1137 9
rect 1168 -9 1185 9
rect 1216 -9 1233 9
rect 1264 -9 1281 9
<< metal1 >>
rect 0 342 1296 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 592 342
rect 609 325 640 342
rect 657 325 688 342
rect 705 325 736 342
rect 753 325 784 342
rect 801 325 832 342
rect 849 325 880 342
rect 897 325 928 342
rect 945 325 976 342
rect 993 325 1024 342
rect 1041 325 1072 342
rect 1089 325 1120 342
rect 1137 325 1168 342
rect 1185 325 1216 342
rect 1233 325 1264 342
rect 1281 325 1296 342
rect 0 309 1296 325
rect 58 299 87 309
rect 58 282 64 299
rect 81 282 87 299
rect 322 299 351 309
rect 322 282 328 299
rect 345 282 351 299
rect 610 299 639 309
rect 610 282 616 299
rect 633 282 639 299
rect 898 299 927 309
rect 898 282 904 299
rect 921 282 927 299
rect 58 276 87 282
rect 137 268 295 282
rect 322 276 351 282
rect 137 207 151 268
rect 178 243 207 249
rect 178 226 184 243
rect 201 226 207 243
rect 178 220 207 226
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 137 114 151 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 185 106 199 220
rect 281 207 295 268
rect 425 268 583 282
rect 610 276 639 282
rect 425 207 439 268
rect 466 243 495 249
rect 466 226 472 243
rect 489 226 495 243
rect 466 220 495 226
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 425 114 439 178
rect 418 108 447 114
rect 418 106 424 108
rect 185 92 424 106
rect 185 73 199 92
rect 418 91 424 92
rect 441 91 447 108
rect 418 85 447 91
rect 473 106 487 220
rect 569 207 583 268
rect 713 268 871 282
rect 898 276 927 282
rect 1186 299 1215 309
rect 1186 282 1192 299
rect 1209 282 1215 299
rect 1186 276 1215 282
rect 713 207 727 268
rect 754 243 783 249
rect 754 226 760 243
rect 777 226 783 243
rect 754 220 783 226
rect 562 201 591 207
rect 562 184 568 201
rect 585 184 591 201
rect 562 178 591 184
rect 706 201 735 207
rect 706 184 712 201
rect 729 184 735 201
rect 706 178 735 184
rect 713 114 727 178
rect 706 108 735 114
rect 706 106 712 108
rect 473 92 712 106
rect 473 73 487 92
rect 706 91 712 92
rect 729 91 735 108
rect 706 85 735 91
rect 761 106 775 220
rect 857 207 871 268
rect 1042 243 1071 249
rect 1042 226 1048 243
rect 1065 226 1071 243
rect 1042 220 1071 226
rect 850 201 879 207
rect 850 184 856 201
rect 873 184 879 201
rect 850 178 879 184
rect 994 201 1023 207
rect 994 184 1000 201
rect 1017 184 1023 201
rect 994 178 1023 184
rect 1001 114 1015 178
rect 1049 154 1063 220
rect 1138 201 1167 207
rect 1138 184 1144 201
rect 1161 184 1167 201
rect 1138 178 1167 184
rect 1042 148 1071 154
rect 1042 131 1048 148
rect 1065 131 1071 148
rect 1042 125 1071 131
rect 1145 114 1159 178
rect 994 108 1023 114
rect 994 106 1000 108
rect 761 92 1000 106
rect 761 73 775 92
rect 994 91 1000 92
rect 1017 106 1023 108
rect 1138 108 1167 114
rect 1138 106 1144 108
rect 1017 92 1144 106
rect 1017 91 1023 92
rect 994 85 1023 91
rect 1138 91 1144 92
rect 1161 91 1167 108
rect 1138 85 1167 91
rect 178 67 207 73
rect 58 51 87 57
rect 58 34 64 51
rect 81 34 87 51
rect 178 50 184 67
rect 201 50 207 67
rect 466 67 495 73
rect 178 44 207 50
rect 322 51 351 57
rect 58 24 87 34
rect 322 34 328 51
rect 345 34 351 51
rect 466 50 472 67
rect 489 50 495 67
rect 754 67 783 73
rect 466 44 495 50
rect 610 51 639 57
rect 322 24 351 34
rect 610 34 616 51
rect 633 34 639 51
rect 754 50 760 67
rect 777 50 783 67
rect 754 44 783 50
rect 898 51 927 57
rect 610 24 639 34
rect 898 34 904 51
rect 921 34 927 51
rect 898 24 927 34
rect 1186 51 1215 57
rect 1186 34 1192 51
rect 1209 34 1215 51
rect 1186 24 1215 34
rect 0 9 1296 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 592 9
rect 609 -9 640 9
rect 657 -9 688 9
rect 705 -9 736 9
rect 753 -9 784 9
rect 801 -9 832 9
rect 849 -9 880 9
rect 897 -9 928 9
rect 945 -9 976 9
rect 993 -9 1024 9
rect 1041 -9 1072 9
rect 1089 -9 1120 9
rect 1137 -9 1168 9
rect 1185 -9 1216 9
rect 1233 -9 1264 9
rect 1281 -9 1296 9
rect 0 -24 1296 -9
<< labels >>
rlabel locali 0 309 1296 357 0 VDD
port 1 se
rlabel metal1 0 309 1296 357 0 VDD
port 2 se
rlabel locali 0 -24 1296 24 0 GND
port 3 se
rlabel metal1 0 -24 1296 24 0 GND
port 4 se
rlabel metal1 1042 125 1071 154 0 Y
port 5 se
rlabel metal1 1049 154 1063 220 0 Y
port 6 se
rlabel metal1 1042 220 1071 249 0 Y
port 7 se
rlabel metal1 130 85 159 114 0 A
port 8 se
rlabel metal1 137 114 151 178 0 A
port 9 se
rlabel metal1 130 178 159 207 0 A
port 10 se
rlabel metal1 274 178 303 207 0 A
port 11 se
rlabel metal1 137 207 151 268 0 A
port 12 se
rlabel metal1 281 207 295 268 0 A
port 13 se
rlabel metal1 137 268 295 282 0 A
port 14 se
<< properties >>
string FIXED_BBOX 0 0 1296 333
<< end >>
