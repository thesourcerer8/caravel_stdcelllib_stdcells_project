VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.310 1.580 0.360 ;
        RECT 0.080 0.290 0.090 0.310 ;
        RECT 0.200 0.290 0.210 0.310 ;
        RECT 0.060 0.280 0.090 0.290 ;
        RECT 0.180 0.280 0.210 0.290 ;
        RECT 0.320 0.290 0.330 0.310 ;
        RECT 0.490 0.290 0.500 0.310 ;
        RECT 0.750 0.290 0.760 0.310 ;
        RECT 0.800 0.300 0.810 0.310 ;
        RECT 1.210 0.290 1.220 0.310 ;
        RECT 0.320 0.280 0.350 0.290 ;
        RECT 0.470 0.280 0.500 0.290 ;
        RECT 0.560 0.280 0.590 0.290 ;
        RECT 0.610 0.280 0.640 0.290 ;
        RECT 0.750 0.280 0.780 0.290 ;
        RECT 1.190 0.280 1.220 0.290 ;
        RECT 1.350 0.290 1.360 0.310 ;
        RECT 1.350 0.280 1.380 0.290 ;
        RECT 0.330 0.260 1.160 0.280 ;
        RECT 0.330 0.240 0.340 0.260 ;
        RECT 1.150 0.240 1.160 0.260 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.370 0.870 2.440 ;
        RECT 3.220 2.370 3.510 2.440 ;
        RECT 0.580 2.230 3.510 2.370 ;
        RECT 0.580 2.150 0.870 2.230 ;
        RECT 3.220 2.150 3.510 2.230 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.080 0.290 0.090 0.310 ;
        RECT 0.060 0.280 0.090 0.290 ;
      LAYER li1 ;
        RECT 0.180 0.290 0.200 0.310 ;
      LAYER li1 ;
        RECT 0.200 0.290 0.210 0.310 ;
        RECT 0.180 0.280 0.210 0.290 ;
        RECT 0.320 0.290 0.330 0.310 ;
        RECT 0.460 0.290 0.470 0.310 ;
        RECT 0.490 0.290 0.500 0.310 ;
        RECT 0.750 0.290 0.760 0.310 ;
        RECT 0.780 0.290 0.790 0.310 ;
        RECT 0.800 0.290 0.810 0.310 ;
        RECT 0.320 0.280 0.350 0.290 ;
        RECT 0.460 0.280 0.500 0.290 ;
        RECT 0.610 0.280 0.640 0.290 ;
        RECT 0.750 0.280 0.810 0.290 ;
        RECT 1.180 0.290 1.190 0.310 ;
        RECT 1.210 0.290 1.220 0.310 ;
        RECT 1.180 0.280 1.220 0.290 ;
        RECT 1.350 0.290 1.360 0.310 ;
        RECT 1.380 0.290 1.390 0.310 ;
        RECT 1.350 0.280 1.390 0.290 ;
        RECT 0.610 0.260 0.620 0.280 ;
        RECT 0.630 0.260 0.640 0.280 ;
        RECT 0.060 0.240 0.110 0.250 ;
        RECT 0.180 0.240 0.210 0.250 ;
      LAYER li1 ;
        RECT 0.060 0.220 0.080 0.240 ;
      LAYER li1 ;
        RECT 0.080 0.220 0.090 0.240 ;
        RECT 0.200 0.220 0.210 0.240 ;
        RECT 0.060 0.210 0.110 0.220 ;
        RECT 0.180 0.210 0.210 0.220 ;
        RECT 0.220 0.240 0.260 0.250 ;
        RECT 0.220 0.220 0.230 0.240 ;
        RECT 0.250 0.220 0.260 0.240 ;
        RECT 0.220 0.210 0.260 0.220 ;
        RECT 0.320 0.240 0.380 0.250 ;
        RECT 0.320 0.220 0.330 0.240 ;
        RECT 0.340 0.220 0.350 0.240 ;
        RECT 0.370 0.220 0.380 0.240 ;
        RECT 0.460 0.240 0.500 0.250 ;
        RECT 0.460 0.220 0.470 0.240 ;
        RECT 0.490 0.220 0.500 0.240 ;
        RECT 0.320 0.210 0.380 0.220 ;
        RECT 0.470 0.210 0.500 0.220 ;
        RECT 0.510 0.240 0.550 0.250 ;
        RECT 0.510 0.220 0.520 0.240 ;
        RECT 0.540 0.220 0.550 0.240 ;
        RECT 0.510 0.210 0.550 0.220 ;
        RECT 0.570 0.210 0.590 0.260 ;
        RECT 0.610 0.240 0.640 0.260 ;
        RECT 0.610 0.220 0.620 0.240 ;
        RECT 0.630 0.220 0.640 0.240 ;
        RECT 0.610 0.210 0.640 0.220 ;
        RECT 0.940 0.240 0.980 0.250 ;
        RECT 0.940 0.220 0.950 0.240 ;
        RECT 0.970 0.220 0.980 0.240 ;
        RECT 0.940 0.210 0.980 0.220 ;
        RECT 1.470 0.240 1.510 0.250 ;
        RECT 1.470 0.220 1.480 0.240 ;
        RECT 1.500 0.220 1.510 0.240 ;
        RECT 1.470 0.210 1.510 0.220 ;
        RECT 0.130 0.200 0.160 0.210 ;
        RECT 0.130 0.180 0.140 0.200 ;
      LAYER li1 ;
        RECT 0.140 0.180 0.150 0.200 ;
      LAYER li1 ;
        RECT 0.150 0.180 0.160 0.200 ;
        RECT 0.130 0.170 0.160 0.180 ;
        RECT 0.270 0.200 0.310 0.210 ;
        RECT 0.420 0.200 0.450 0.210 ;
        RECT 0.270 0.180 0.280 0.200 ;
        RECT 0.300 0.180 0.310 0.200 ;
        RECT 0.440 0.180 0.450 0.200 ;
        RECT 0.270 0.170 0.310 0.180 ;
        RECT 0.420 0.170 0.450 0.180 ;
        RECT 0.560 0.200 0.590 0.210 ;
        RECT 0.700 0.200 0.740 0.210 ;
        RECT 0.560 0.180 0.570 0.200 ;
        RECT 0.700 0.180 0.710 0.200 ;
        RECT 0.730 0.180 0.740 0.200 ;
        RECT 0.560 0.170 0.590 0.180 ;
        RECT 0.700 0.170 0.740 0.180 ;
        RECT 0.850 0.200 0.880 0.210 ;
        RECT 0.850 0.180 0.860 0.200 ;
        RECT 0.870 0.180 0.880 0.200 ;
        RECT 0.850 0.170 0.880 0.180 ;
        RECT 0.990 0.200 1.030 0.210 ;
        RECT 1.140 0.200 1.170 0.210 ;
        RECT 0.990 0.180 1.000 0.200 ;
        RECT 1.020 0.180 1.030 0.200 ;
        RECT 1.160 0.180 1.170 0.200 ;
        RECT 0.990 0.170 1.030 0.180 ;
        RECT 1.140 0.170 1.170 0.180 ;
        RECT 1.420 0.200 1.460 0.210 ;
        RECT 1.420 0.180 1.430 0.200 ;
        RECT 1.450 0.180 1.460 0.200 ;
        RECT 1.420 0.170 1.460 0.180 ;
        RECT 0.140 0.110 0.150 0.170 ;
        RECT 0.280 0.140 0.300 0.170 ;
        RECT 0.280 0.110 0.300 0.130 ;
        RECT 0.130 0.100 0.160 0.110 ;
        RECT 0.130 0.090 0.140 0.100 ;
      LAYER li1 ;
        RECT 0.140 0.090 0.150 0.100 ;
      LAYER li1 ;
        RECT 0.150 0.090 0.160 0.100 ;
        RECT 0.130 0.080 0.160 0.090 ;
        RECT 0.270 0.100 0.310 0.110 ;
        RECT 0.420 0.100 0.450 0.110 ;
        RECT 0.270 0.090 0.280 0.100 ;
        RECT 0.300 0.090 0.310 0.100 ;
        RECT 0.440 0.090 0.450 0.100 ;
        RECT 0.270 0.080 0.310 0.090 ;
        RECT 0.420 0.080 0.450 0.090 ;
        RECT 0.520 0.070 0.540 0.130 ;
        RECT 0.560 0.100 0.590 0.110 ;
        RECT 0.700 0.100 0.740 0.110 ;
        RECT 0.560 0.090 0.570 0.100 ;
        RECT 0.700 0.090 0.710 0.100 ;
        RECT 0.730 0.090 0.740 0.100 ;
        RECT 0.560 0.080 0.590 0.090 ;
        RECT 0.700 0.080 0.740 0.090 ;
        RECT 0.850 0.100 0.880 0.110 ;
        RECT 0.850 0.090 0.860 0.100 ;
        RECT 0.870 0.090 0.880 0.100 ;
        RECT 0.850 0.080 0.880 0.090 ;
        RECT 0.990 0.100 1.030 0.110 ;
        RECT 1.140 0.100 1.170 0.110 ;
        RECT 0.990 0.090 1.000 0.100 ;
        RECT 1.020 0.090 1.030 0.100 ;
        RECT 1.160 0.090 1.170 0.100 ;
        RECT 0.990 0.080 1.030 0.090 ;
        RECT 1.140 0.080 1.170 0.090 ;
        RECT 1.420 0.100 1.460 0.110 ;
        RECT 1.420 0.090 1.430 0.100 ;
        RECT 1.450 0.090 1.460 0.100 ;
        RECT 1.420 0.080 1.460 0.090 ;
        RECT 0.060 0.060 0.110 0.070 ;
        RECT 0.320 0.060 0.380 0.070 ;
      LAYER li1 ;
        RECT 0.060 0.050 0.080 0.060 ;
      LAYER li1 ;
        RECT 0.080 0.050 0.090 0.060 ;
        RECT 0.320 0.050 0.330 0.060 ;
        RECT 0.340 0.050 0.350 0.060 ;
        RECT 0.370 0.050 0.380 0.060 ;
        RECT 0.060 0.040 0.110 0.050 ;
        RECT 0.320 0.040 0.380 0.050 ;
        RECT 0.460 0.060 0.500 0.070 ;
        RECT 0.460 0.050 0.470 0.060 ;
        RECT 0.490 0.050 0.500 0.060 ;
        RECT 0.460 0.040 0.500 0.050 ;
        RECT 0.510 0.060 0.550 0.070 ;
        RECT 0.510 0.050 0.520 0.060 ;
        RECT 0.540 0.050 0.550 0.060 ;
        RECT 0.510 0.040 0.550 0.050 ;
        RECT 0.610 0.060 0.640 0.070 ;
        RECT 0.610 0.050 0.620 0.060 ;
        RECT 0.630 0.050 0.640 0.060 ;
        RECT 0.610 0.040 0.640 0.050 ;
        RECT 1.040 0.060 1.070 0.070 ;
        RECT 1.470 0.060 1.510 0.070 ;
        RECT 1.040 0.050 1.050 0.060 ;
        RECT 1.470 0.050 1.480 0.060 ;
        RECT 1.500 0.050 1.510 0.060 ;
        RECT 1.040 0.040 1.070 0.050 ;
        RECT 1.470 0.040 1.510 0.050 ;
      LAYER li1 ;
        RECT 0.180 0.020 0.200 0.040 ;
      LAYER li1 ;
        RECT 0.200 0.020 0.210 0.040 ;
        RECT 0.180 0.010 0.210 0.020 ;
        RECT 0.320 0.020 0.330 0.040 ;
        RECT 0.320 0.010 0.350 0.020 ;
        RECT 0.460 0.010 0.470 0.040 ;
        RECT 0.490 0.010 0.500 0.040 ;
        RECT 0.610 0.010 0.620 0.040 ;
        RECT 0.630 0.010 0.640 0.040 ;
        RECT 0.750 0.020 0.760 0.040 ;
        RECT 0.780 0.020 0.790 0.040 ;
        RECT 0.750 0.010 0.790 0.020 ;
        RECT 0.800 0.010 0.810 0.040 ;
        RECT 0.940 0.020 0.950 0.040 ;
        RECT 0.970 0.020 0.980 0.040 ;
        RECT 1.180 0.020 1.190 0.040 ;
        RECT 1.210 0.020 1.220 0.040 ;
        RECT 0.940 0.010 1.220 0.020 ;
        RECT 1.350 0.010 1.360 0.040 ;
        RECT 1.380 0.010 1.390 0.040 ;
  END
END NAND2X1
END LIBRARY

