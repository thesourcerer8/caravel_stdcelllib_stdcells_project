VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INV
  CLASS CORE ;
  FOREIGN INV ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 2.880 3.570 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.880 0.240 ;
    END
  END vssd1
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.200 0.870 2.490 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 0.580 0.440 0.870 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 2.760 2.090 3.090 ;
        RECT 0.560 2.180 0.890 2.510 ;
        RECT 1.280 1.760 1.610 2.090 ;
        RECT 1.280 0.830 1.610 1.160 ;
        RECT 0.560 0.420 0.890 0.750 ;
        RECT 1.760 0.240 2.090 0.570 ;
  END
END INV
END LIBRARY

