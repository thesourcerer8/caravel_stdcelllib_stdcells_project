magic
tech sky130A
magscale 1 2
timestamp 1636962384
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1152 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 931 134 989 146
rect 931 132 943 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 48 561 132
rect 591 48 849 132
rect 879 100 943 132
rect 977 132 989 134
rect 977 100 1037 132
rect 879 48 1037 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 593 561 618
rect 303 559 367 593
rect 401 559 561 593
rect 303 450 561 559
rect 591 485 849 618
rect 591 451 655 485
rect 689 451 849 485
rect 591 450 849 451
rect 879 593 1037 618
rect 879 559 943 593
rect 977 559 1037 593
rect 879 450 1037 559
rect 115 439 173 450
rect 643 439 701 450
<< ndiffc >>
rect 127 100 161 134
rect 943 100 977 134
<< pdiffc >>
rect 127 451 161 485
rect 367 559 401 593
rect 655 451 689 485
rect 943 559 977 593
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1152 683
rect 31 643 1121 649
rect 31 618 893 643
rect 1027 618 1121 643
rect 351 593 417 618
rect 351 559 367 593
rect 401 559 417 593
rect 351 543 417 559
rect 927 593 993 609
rect 927 559 943 593
rect 977 559 993 593
rect 927 543 993 559
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 111 435 177 451
rect 639 485 705 501
rect 639 451 655 485
rect 689 451 705 485
rect 639 435 705 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 605 418
rect 543 368 559 402
rect 593 401 605 402
rect 831 402 897 418
rect 593 368 609 401
rect 543 352 609 368
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 881 181 893 184
rect 831 165 893 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 927 134 993 150
rect 927 100 943 134
rect 977 100 993 134
rect 927 84 993 100
rect 31 17 1121 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1152 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 367 559 401 593
rect 943 559 977 593
rect 127 451 161 485
rect 655 451 689 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 127 100 161 134
rect 943 100 977 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1152 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1152 683
rect 0 618 1152 649
rect 355 593 413 618
rect 355 559 367 593
rect 401 559 413 593
rect 355 547 413 559
rect 931 593 989 618
rect 931 559 943 593
rect 977 559 989 593
rect 931 547 989 559
rect 115 485 173 497
rect 115 451 127 485
rect 161 482 173 485
rect 643 485 701 497
rect 643 482 655 485
rect 161 454 655 482
rect 161 451 173 454
rect 115 439 173 451
rect 643 451 655 454
rect 689 451 701 485
rect 643 439 701 451
rect 130 146 158 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 274 227 302 356
rect 562 227 590 356
rect 850 227 878 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 835 215 893 227
rect 835 181 847 215
rect 881 181 893 215
rect 835 169 893 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 931 134 989 146
rect 931 100 943 134
rect 977 100 989 134
rect 931 88 989 100
rect 946 48 974 88
rect 0 17 1152 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1152 17
rect 0 -48 1152 -17
<< labels >>
rlabel metal1 0 618 1152 714 0 VPWR
port 4 se
rlabel metal1 0 618 1152 714 0 VPWR
port 4 se
rlabel metal1 0 -48 1152 48 0 VGND
port 3 se
rlabel metal1 0 -48 1152 48 0 VGND
port 3 se
rlabel metal1 115 88 173 146 0 Y
port 5 se
rlabel metal1 130 146 158 439 0 Y
port 5 se
rlabel metal1 115 439 173 454 0 Y
port 5 se
rlabel metal1 643 439 701 454 0 Y
port 5 se
rlabel metal1 115 454 701 482 0 Y
port 5 se
rlabel metal1 115 482 173 497 0 Y
port 5 se
rlabel metal1 643 482 701 497 0 Y
port 5 se
rlabel metal1 547 169 605 227 0 B
port 1 se
rlabel metal1 562 227 590 356 0 B
port 1 se
rlabel metal1 547 356 605 414 0 B
port 1 se
rlabel metal1 835 169 893 227 0 A
port 0 se
rlabel metal1 850 227 878 356 0 A
port 0 se
rlabel metal1 835 356 893 414 0 A
port 0 se
rlabel metal1 259 169 317 227 0 C
port 2 se
rlabel metal1 274 227 302 356 0 C
port 2 se
rlabel metal1 259 356 317 414 0 C
port 2 se
rlabel locali 0 -17 1152 17 4 VGND
port 3 se ground default abutment
rlabel locali 31 17 1121 48 4 VGND
port 3 se ground default abutment
rlabel locali 0 649 1152 683 4 VPWR
port 4 se power default abutment
rlabel metal1 31 618 1121 649 4 VGND
port 3 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1152 666
<< end >>
