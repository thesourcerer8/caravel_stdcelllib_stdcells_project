magic
tech sky130A
timestamp 1623602984
<< nwell >>
rect 0 179 576 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
<< ndiff >>
rect 58 66 87 69
rect 58 63 137 66
rect 58 46 64 63
rect 81 46 137 63
rect 58 24 137 46
rect 152 24 281 66
rect 296 24 425 66
rect 440 36 519 66
rect 440 24 472 36
rect 466 19 472 24
rect 489 24 519 36
rect 489 19 495 24
rect 466 13 495 19
<< pdiff >>
rect 178 309 207 312
rect 466 309 495 312
rect 58 238 137 309
rect 58 221 64 238
rect 81 225 137 238
rect 152 306 281 309
rect 152 289 184 306
rect 201 289 281 306
rect 152 225 281 289
rect 296 238 425 309
rect 296 225 328 238
rect 81 221 87 225
rect 58 215 87 221
rect 322 221 328 225
rect 345 225 425 238
rect 440 306 519 309
rect 440 289 472 306
rect 489 289 519 306
rect 440 225 519 289
rect 345 221 351 225
rect 322 215 351 221
<< ndiffc >>
rect 64 46 81 63
rect 472 19 489 36
<< pdiffc >>
rect 64 221 81 238
rect 184 289 201 306
rect 328 221 345 238
rect 472 289 489 306
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 464 306 497 314
rect 464 289 472 306
rect 489 289 497 306
rect 464 281 497 289
rect 56 238 89 246
rect 56 221 64 238
rect 81 221 89 238
rect 56 213 89 221
rect 320 238 353 246
rect 320 221 328 238
rect 345 221 353 238
rect 320 213 353 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 303 206
rect 272 181 280 198
rect 297 196 303 198
rect 416 198 449 206
rect 297 181 305 196
rect 272 173 305 181
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 56 63 89 71
rect 56 46 64 63
rect 81 46 89 63
rect 56 38 89 46
rect 464 36 497 44
rect 464 19 472 36
rect 489 19 497 36
rect 464 11 497 19
<< viali >>
rect 184 289 201 306
rect 472 289 489 306
rect 64 221 81 238
rect 328 221 345 238
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 64 46 81 63
rect 472 19 489 36
<< metal1 >>
rect 0 309 576 357
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 466 306 495 309
rect 466 289 472 306
rect 489 289 495 306
rect 466 283 495 289
rect 58 238 87 244
rect 58 221 64 238
rect 81 237 87 238
rect 322 238 351 244
rect 322 237 328 238
rect 81 223 328 237
rect 81 221 87 223
rect 58 215 87 221
rect 322 221 328 223
rect 345 221 351 238
rect 322 215 351 221
rect 65 69 79 215
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 274 198 303 204
rect 274 181 280 198
rect 297 181 303 198
rect 274 175 303 181
rect 418 198 447 204
rect 418 181 424 198
rect 441 181 447 198
rect 418 175 447 181
rect 137 109 151 175
rect 281 109 295 175
rect 425 109 439 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 86 159 103
rect 130 80 159 86
rect 274 103 303 109
rect 274 86 280 103
rect 297 86 303 103
rect 274 80 303 86
rect 418 103 447 109
rect 418 86 424 103
rect 441 86 447 103
rect 418 80 447 86
rect 58 63 87 69
rect 58 46 64 63
rect 81 46 87 63
rect 58 40 87 46
rect 466 36 495 42
rect 466 24 472 36
rect 0 19 472 24
rect 489 24 495 36
rect 489 19 576 24
rect 0 -24 576 19
<< labels >>
rlabel metal1 0 309 576 357 0 VDD
port 1 se
rlabel metal1 0 -24 576 24 0 GND
port 2 se
rlabel metal1 58 40 87 69 0 Y
port 3 se
rlabel metal1 65 69 79 215 0 Y
port 4 se
rlabel metal1 58 215 87 223 0 Y
port 5 se
rlabel metal1 322 215 351 223 0 Y
port 6 se
rlabel metal1 58 223 351 237 0 Y
port 7 se
rlabel metal1 58 237 87 244 0 Y
port 8 se
rlabel metal1 322 237 351 244 0 Y
port 9 se
rlabel metal1 418 80 447 109 0 A
port 10 se
rlabel metal1 425 109 439 175 0 A
port 11 se
rlabel metal1 418 175 447 204 0 A
port 12 se
rlabel metal1 130 80 159 109 0 C
port 13 se
rlabel metal1 137 109 151 175 0 C
port 14 se
rlabel metal1 130 175 159 204 0 C
port 15 se
rlabel metal1 274 80 303 109 0 B
port 16 se
rlabel metal1 281 109 295 175 0 B
port 17 se
rlabel metal1 274 175 303 204 0 B
port 18 se
<< properties >>
string FIXED_BBOX 0 0 576 333
<< end >>
