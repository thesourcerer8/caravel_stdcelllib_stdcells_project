VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.995 1.585 2.070 ;
        RECT 5.615 1.995 5.905 2.070 ;
        RECT 1.295 1.855 5.905 1.995 ;
        RECT 1.295 1.780 1.585 1.855 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 4.250 1.135 4.390 1.855 ;
        RECT 5.615 1.780 5.905 1.855 ;
        RECT 1.295 0.845 1.585 1.135 ;
        RECT 4.175 0.845 4.465 1.135 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
      LAYER mcon ;
        RECT 4.235 0.905 4.405 1.075 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.275 1.760 1.605 2.090 ;
      LAYER mcon ;
        RECT 1.355 1.840 1.525 2.010 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.595 1.760 5.925 2.090 ;
      LAYER mcon ;
        RECT 5.675 1.840 5.845 2.010 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 2.815 3.025 2.890 ;
        RECT 2.735 2.675 8.710 2.815 ;
        RECT 2.735 2.600 3.025 2.675 ;
        RECT 8.570 2.070 8.710 2.675 ;
        RECT 8.495 1.780 8.785 2.070 ;
        RECT 2.735 1.385 3.025 1.675 ;
        RECT 2.810 1.135 2.950 1.385 ;
        RECT 2.735 0.845 3.025 1.135 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.795 2.090 2.965 2.830 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 2.795 1.445 2.965 1.760 ;
      LAYER mcon ;
        RECT 2.795 2.660 2.965 2.830 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.240 2.065 0.570 ;
        RECT 7.535 0.240 7.825 0.570 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.755 0.240 2.085 0.590 ;
        RECT 7.515 0.240 7.845 0.590 ;
        RECT 0.155 0.085 9.925 0.240 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 1.835 0.340 2.005 0.510 ;
        RECT 7.595 0.340 7.765 0.510 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.775 2.760 2.065 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 2.167200 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.155 3.090 9.925 3.245 ;
        RECT 1.755 2.740 2.085 3.090 ;
        RECT 7.515 2.740 7.845 3.090 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 1.835 2.820 2.005 2.990 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 4.655 0.440 4.945 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 10.080 3.330 ;
      LAYER li1 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 4.235 2.090 4.405 2.425 ;
        RECT 4.635 2.260 4.965 2.505 ;
        RECT 8.955 2.260 9.285 2.505 ;
        RECT 4.655 2.175 4.965 2.260 ;
        RECT 8.975 2.175 9.285 2.260 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 4.715 0.750 4.885 2.175 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 8.555 1.155 8.725 1.760 ;
        RECT 5.595 0.825 5.925 1.155 ;
        RECT 7.035 0.825 7.365 1.155 ;
        RECT 8.475 0.825 8.805 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 8.975 0.655 9.285 0.750 ;
        RECT 8.955 0.420 9.285 0.655 ;
      LAYER mcon ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 4.235 2.255 4.405 2.425 ;
        RECT 9.035 2.255 9.205 2.425 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 7.115 1.840 7.285 2.010 ;
        RECT 8.555 1.840 8.725 2.010 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 7.115 0.905 7.285 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 9.035 0.500 9.205 0.670 ;
      LAYER met1 ;
        RECT 0.575 2.410 0.865 2.485 ;
        RECT 4.175 2.410 4.465 2.485 ;
        RECT 0.575 2.270 6.310 2.410 ;
        RECT 0.575 2.195 0.865 2.270 ;
        RECT 4.175 2.195 4.465 2.270 ;
        RECT 0.650 0.730 0.790 2.195 ;
        RECT 5.615 1.060 5.905 1.135 ;
        RECT 6.170 1.060 6.310 2.270 ;
        RECT 8.975 2.195 9.265 2.485 ;
        RECT 7.055 1.780 7.345 2.070 ;
        RECT 7.130 1.135 7.270 1.780 ;
        RECT 5.615 0.920 6.310 1.060 ;
        RECT 7.055 1.060 7.345 1.135 ;
        RECT 9.050 1.060 9.190 2.195 ;
        RECT 7.055 0.920 9.190 1.060 ;
        RECT 5.615 0.845 5.905 0.920 ;
        RECT 7.055 0.845 7.345 0.920 ;
        RECT 9.050 0.730 9.190 0.920 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 8.975 0.440 9.265 0.730 ;
  END
END XOR2X1
END LIBRARY

