VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 1.780 3.010 2.070 3.090 ;
        RECT 1.780 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.070 3.010 ;
        RECT 1.780 2.780 2.070 2.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.490 2.070 0.550 ;
        RECT 1.780 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.070 0.490 ;
        RECT 1.780 0.240 2.070 0.320 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
  END vssd1
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.820 2.410 1.110 2.490 ;
        RECT 3.220 2.410 3.510 2.490 ;
        RECT 0.820 2.270 3.510 2.410 ;
        RECT 0.820 2.200 1.110 2.270 ;
        RECT 3.220 2.200 3.510 2.270 ;
        RECT 0.890 0.730 1.030 2.200 ;
        RECT 3.290 0.730 3.430 2.200 ;
        RECT 0.820 0.440 1.110 0.730 ;
        RECT 3.220 0.440 3.510 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 1.300 1.060 1.590 1.140 ;
        RECT 2.740 1.060 3.030 1.140 ;
        RECT 1.300 0.920 3.030 1.060 ;
        RECT 1.300 0.850 1.590 0.920 ;
        RECT 2.740 0.850 3.030 0.920 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 3.010 2.090 3.090 ;
        RECT 1.760 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.090 3.010 ;
        RECT 1.760 2.760 2.090 2.840 ;
        RECT 0.800 2.430 1.130 2.510 ;
        RECT 0.800 2.260 0.880 2.430 ;
        RECT 1.050 2.260 1.130 2.430 ;
        RECT 3.200 2.430 3.530 2.510 ;
        RECT 3.200 2.260 3.280 2.430 ;
        RECT 3.450 2.260 3.530 2.430 ;
        RECT 0.800 2.180 1.110 2.260 ;
        RECT 3.220 2.180 3.530 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.920 1.360 1.080 ;
        RECT 1.300 0.910 1.360 0.920 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.300 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 0.800 0.670 1.130 0.750 ;
        RECT 0.800 0.500 0.880 0.670 ;
        RECT 1.050 0.500 1.130 0.670 ;
        RECT 3.220 0.670 3.530 0.750 ;
        RECT 3.220 0.660 3.280 0.670 ;
        RECT 0.800 0.420 1.130 0.500 ;
        RECT 1.760 0.490 2.090 0.570 ;
        RECT 1.760 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.090 0.490 ;
        RECT 3.200 0.500 3.280 0.660 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
        RECT 1.760 0.240 2.090 0.320 ;
  END
END INVX4
END LIBRARY

