magic
tech sky130A
timestamp 1621277262
<< end >>
