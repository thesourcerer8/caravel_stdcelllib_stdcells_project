magic
tech sky130A
timestamp 1623602966
<< nwell >>
rect 0 179 720 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
<< ndiff >>
rect 58 66 87 69
rect 322 66 351 69
rect 610 66 639 69
rect 58 63 137 66
rect 58 46 64 63
rect 81 46 137 63
rect 58 24 137 46
rect 152 36 281 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 281 36
rect 296 63 425 66
rect 296 46 328 63
rect 345 46 425 63
rect 296 24 425 46
rect 440 36 569 66
rect 440 24 472 36
rect 201 19 207 24
rect 178 13 207 19
rect 466 19 472 24
rect 489 24 569 36
rect 584 63 663 66
rect 584 46 616 63
rect 633 46 663 63
rect 584 24 663 46
rect 489 19 495 24
rect 466 13 495 19
<< pdiff >>
rect 178 309 207 312
rect 466 309 495 312
rect 58 238 137 309
rect 58 221 64 238
rect 81 225 137 238
rect 152 306 281 309
rect 152 289 184 306
rect 201 289 281 306
rect 152 225 281 289
rect 296 238 425 309
rect 296 225 328 238
rect 81 221 87 225
rect 58 215 87 221
rect 322 221 328 225
rect 345 225 425 238
rect 440 306 569 309
rect 440 289 472 306
rect 489 289 569 306
rect 440 225 569 289
rect 584 238 663 309
rect 584 225 616 238
rect 345 221 351 225
rect 322 215 351 221
rect 610 221 616 225
rect 633 225 663 238
rect 633 221 639 225
rect 610 215 639 221
<< ndiffc >>
rect 64 46 81 63
rect 184 19 201 36
rect 328 46 345 63
rect 472 19 489 36
rect 616 46 633 63
<< pdiffc >>
rect 64 221 81 238
rect 184 289 201 306
rect 328 221 345 238
rect 472 289 489 306
rect 616 221 633 238
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 569 309 584 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 569 206 584 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 569 66 584 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 464 306 497 314
rect 464 289 472 306
rect 489 289 497 306
rect 464 281 497 289
rect 56 238 89 246
rect 56 221 64 238
rect 81 221 89 238
rect 320 238 353 246
rect 320 223 328 238
rect 56 213 89 221
rect 322 221 328 223
rect 345 221 353 238
rect 608 238 641 246
rect 608 223 616 238
rect 322 213 353 221
rect 610 221 616 223
rect 633 221 641 238
rect 610 213 641 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 88 305 103
rect 416 103 449 111
rect 297 86 303 88
rect 272 78 303 86
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 56 63 89 71
rect 56 46 64 63
rect 81 46 89 63
rect 56 38 89 46
rect 320 63 353 71
rect 320 46 328 63
rect 345 46 353 63
rect 610 63 641 71
rect 610 61 616 63
rect 176 36 209 44
rect 320 38 353 46
rect 608 46 616 61
rect 633 46 641 63
rect 176 11 184 36
rect 201 11 209 36
rect 464 36 497 44
rect 608 38 641 46
rect 464 11 472 36
rect 489 11 497 36
<< viali >>
rect 184 289 201 306
rect 472 289 489 306
rect 64 221 81 238
rect 328 221 345 238
rect 616 221 633 238
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
rect 64 46 81 63
rect 328 46 345 63
rect 616 46 633 63
rect 184 19 201 22
rect 184 5 201 19
rect 472 19 489 22
rect 472 5 489 19
<< metal1 >>
rect 0 309 720 357
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 466 306 495 309
rect 466 289 472 306
rect 489 289 495 306
rect 466 283 495 289
rect 58 238 87 244
rect 58 221 64 238
rect 81 237 87 238
rect 322 238 351 244
rect 322 237 328 238
rect 81 223 328 237
rect 81 221 87 223
rect 58 215 87 221
rect 322 221 328 223
rect 345 221 351 238
rect 322 215 351 221
rect 610 238 639 244
rect 610 221 616 238
rect 633 221 639 238
rect 610 215 639 221
rect 65 69 79 215
rect 130 198 159 204
rect 130 181 136 198
rect 153 196 159 198
rect 274 198 303 204
rect 274 196 280 198
rect 153 182 280 196
rect 153 181 159 182
rect 130 175 159 181
rect 274 181 280 182
rect 297 196 303 198
rect 418 198 447 204
rect 418 196 424 198
rect 297 182 424 196
rect 297 181 303 182
rect 274 175 303 181
rect 418 181 424 182
rect 441 196 447 198
rect 562 198 591 204
rect 562 196 568 198
rect 441 182 568 196
rect 441 181 447 182
rect 418 175 447 181
rect 562 181 568 182
rect 585 181 591 198
rect 562 175 591 181
rect 137 109 151 175
rect 281 109 295 175
rect 425 109 439 175
rect 569 109 583 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 86 159 103
rect 130 80 159 86
rect 274 103 303 109
rect 274 86 280 103
rect 297 86 303 103
rect 274 80 303 86
rect 418 103 447 109
rect 418 86 424 103
rect 441 86 447 103
rect 418 80 447 86
rect 562 103 591 109
rect 562 86 568 103
rect 585 86 591 103
rect 562 80 591 86
rect 617 69 631 215
rect 58 63 87 69
rect 58 46 64 63
rect 81 61 87 63
rect 322 63 351 69
rect 322 61 328 63
rect 81 47 328 61
rect 81 46 87 47
rect 58 40 87 46
rect 322 46 328 47
rect 345 61 351 63
rect 610 63 639 69
rect 610 61 616 63
rect 345 47 616 61
rect 345 46 351 47
rect 322 40 351 46
rect 610 46 616 47
rect 633 46 639 63
rect 610 40 639 46
rect 178 24 207 28
rect 466 24 495 28
rect 0 22 720 24
rect 0 5 184 22
rect 201 5 472 22
rect 489 5 720 22
rect 0 -24 720 5
<< labels >>
rlabel metal1 0 309 720 357 0 VDD
port 1 se
rlabel metal1 0 -24 720 24 0 GND
port 2 se
rlabel metal1 58 40 87 47 0 Y
port 3 se
rlabel metal1 322 40 351 47 0 Y
port 4 se
rlabel metal1 610 40 639 47 0 Y
port 5 se
rlabel metal1 58 47 639 61 0 Y
port 6 se
rlabel metal1 58 61 87 69 0 Y
port 7 se
rlabel metal1 322 61 351 69 0 Y
port 8 se
rlabel metal1 610 61 639 69 0 Y
port 9 se
rlabel metal1 65 69 79 215 0 Y
port 10 se
rlabel metal1 617 69 631 215 0 Y
port 11 se
rlabel metal1 58 215 87 223 0 Y
port 12 se
rlabel metal1 322 215 351 223 0 Y
port 13 se
rlabel metal1 58 223 351 237 0 Y
port 14 se
rlabel metal1 58 237 87 244 0 Y
port 15 se
rlabel metal1 322 237 351 244 0 Y
port 16 se
rlabel metal1 610 215 639 244 0 Y
port 17 se
rlabel metal1 130 80 159 109 0 A
port 18 se
rlabel metal1 274 80 303 109 0 A
port 19 se
rlabel metal1 418 80 447 109 0 A
port 20 se
rlabel metal1 562 80 591 109 0 A
port 21 se
rlabel metal1 137 109 151 175 0 A
port 22 se
rlabel metal1 281 109 295 175 0 A
port 23 se
rlabel metal1 425 109 439 175 0 A
port 24 se
rlabel metal1 569 109 583 175 0 A
port 25 se
rlabel metal1 130 175 159 182 0 A
port 26 se
rlabel metal1 274 175 303 182 0 A
port 27 se
rlabel metal1 418 175 447 182 0 A
port 28 se
rlabel metal1 562 175 591 182 0 A
port 29 se
rlabel metal1 130 182 591 196 0 A
port 30 se
rlabel metal1 130 196 159 204 0 A
port 31 se
rlabel metal1 274 196 303 204 0 A
port 32 se
rlabel metal1 418 196 447 204 0 A
port 33 se
rlabel metal1 562 196 591 204 0 A
port 34 se
<< properties >>
string FIXED_BBOX 0 0 720 333
<< end >>
