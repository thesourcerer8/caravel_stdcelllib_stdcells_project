VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
        RECT 1.780 3.060 2.070 3.090 ;
        RECT 1.780 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.070 3.060 ;
        RECT 1.780 2.830 2.070 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.220 0.240 3.510 0.280 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.150 4.950 2.440 ;
        RECT 0.820 0.610 1.110 0.690 ;
        RECT 4.730 0.610 4.870 2.150 ;
        RECT 6.100 0.610 6.390 0.690 ;
        RECT 0.820 0.470 6.390 0.610 ;
        RECT 0.820 0.400 1.110 0.470 ;
        RECT 6.100 0.400 6.390 0.470 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END A
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.750 4.470 2.040 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 4.180 0.800 4.470 1.090 ;
    END
  END C
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.750 5.910 2.040 ;
        RECT 5.690 1.090 5.830 1.750 ;
        RECT 5.620 0.800 5.910 1.090 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 1.760 3.060 2.090 3.140 ;
        RECT 1.760 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.090 3.060 ;
        RECT 1.760 2.810 2.090 2.890 ;
        RECT 6.080 2.790 6.410 2.870 ;
        RECT 6.080 2.620 6.160 2.790 ;
        RECT 6.330 2.620 6.410 2.790 ;
        RECT 6.080 2.540 6.410 2.620 ;
        RECT 0.800 2.380 1.130 2.460 ;
        RECT 0.800 2.210 0.880 2.380 ;
        RECT 1.050 2.210 1.130 2.380 ;
        RECT 3.200 2.380 3.530 2.460 ;
        RECT 3.200 2.230 3.280 2.380 ;
        RECT 0.800 2.130 1.130 2.210 ;
        RECT 3.220 2.210 3.280 2.230 ;
        RECT 3.450 2.210 3.530 2.380 ;
        RECT 4.640 2.380 4.970 2.460 ;
        RECT 4.640 2.230 4.720 2.380 ;
        RECT 3.220 2.130 3.530 2.210 ;
        RECT 4.660 2.210 4.720 2.230 ;
        RECT 4.890 2.210 4.970 2.380 ;
        RECT 4.660 2.130 4.970 2.210 ;
        RECT 1.300 1.980 1.610 2.060 ;
        RECT 1.300 1.960 1.360 1.980 ;
        RECT 1.280 1.810 1.360 1.960 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 2.720 1.980 3.050 2.060 ;
        RECT 2.720 1.810 2.800 1.980 ;
        RECT 2.970 1.810 3.050 1.980 ;
        RECT 2.720 1.730 3.050 1.810 ;
        RECT 4.160 1.980 4.490 2.060 ;
        RECT 4.160 1.810 4.240 1.980 ;
        RECT 4.410 1.810 4.490 1.980 ;
        RECT 4.160 1.730 4.490 1.810 ;
        RECT 5.600 1.980 5.930 2.060 ;
        RECT 5.600 1.810 5.680 1.980 ;
        RECT 5.850 1.810 5.930 1.980 ;
        RECT 5.600 1.730 5.930 1.810 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.860 1.360 1.030 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.280 0.780 1.610 0.860 ;
        RECT 2.720 1.030 3.050 1.110 ;
        RECT 2.720 0.860 2.800 1.030 ;
        RECT 2.970 0.860 3.050 1.030 ;
        RECT 2.720 0.780 3.050 0.860 ;
        RECT 4.160 1.030 4.490 1.110 ;
        RECT 4.160 0.860 4.240 1.030 ;
        RECT 4.410 0.860 4.490 1.030 ;
        RECT 4.160 0.780 4.490 0.860 ;
        RECT 5.600 1.030 5.930 1.110 ;
        RECT 5.600 0.860 5.680 1.030 ;
        RECT 5.850 0.880 5.930 1.030 ;
        RECT 5.850 0.860 5.910 0.880 ;
        RECT 5.600 0.780 5.910 0.860 ;
        RECT 0.800 0.630 1.110 0.710 ;
        RECT 0.800 0.460 0.880 0.630 ;
        RECT 1.050 0.610 1.110 0.630 ;
        RECT 6.080 0.630 6.410 0.710 ;
        RECT 1.050 0.460 1.130 0.610 ;
        RECT 0.800 0.380 1.130 0.460 ;
        RECT 6.080 0.460 6.160 0.630 ;
        RECT 6.330 0.460 6.410 0.630 ;
        RECT 3.200 0.360 3.530 0.440 ;
        RECT 6.080 0.380 6.410 0.460 ;
        RECT 3.200 0.110 3.280 0.360 ;
        RECT 3.450 0.110 3.530 0.360 ;
      LAYER met1 ;
        RECT 6.100 2.790 6.390 2.850 ;
        RECT 6.100 2.770 6.160 2.790 ;
        RECT 3.290 2.630 6.160 2.770 ;
        RECT 3.290 2.440 3.430 2.630 ;
        RECT 6.100 2.620 6.160 2.630 ;
        RECT 6.330 2.620 6.390 2.790 ;
        RECT 6.100 2.560 6.390 2.620 ;
        RECT 0.820 2.380 1.110 2.440 ;
        RECT 0.820 2.210 0.880 2.380 ;
        RECT 1.050 2.370 1.110 2.380 ;
        RECT 3.220 2.380 3.510 2.440 ;
        RECT 3.220 2.370 3.280 2.380 ;
        RECT 1.050 2.230 3.280 2.370 ;
        RECT 1.050 2.210 1.110 2.230 ;
        RECT 0.820 2.150 1.110 2.210 ;
        RECT 3.220 2.210 3.280 2.230 ;
        RECT 3.450 2.210 3.510 2.380 ;
        RECT 3.220 2.150 3.510 2.210 ;
  END
END AOI22X1
END LIBRARY

