magic
tech sky130A
timestamp 1621277560
<< end >>
