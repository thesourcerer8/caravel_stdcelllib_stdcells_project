magic
tech sky130A
timestamp 1621277284
<< end >>
