MACRO INV
 CLASS CORE ;
 FOREIGN INV 0 0 ;
 SIZE 2.88 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 2.88000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 2.88000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 2.88000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 2.88000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.57500000 0.44000000 0.86500000 0.73000000 ;
        RECT 0.65000000 0.73000000 0.79000000 2.19500000 ;
        RECT 0.57500000 2.19500000 0.86500000 2.48500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 1.83500000 2.79500000 2.00500000 2.96500000 ;

    LAYER ndiffc ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 1.83500000 0.50000000 2.00500000 0.67000000 ;

    LAYER li1 ;
     RECT 0.00000000 -0.24000000 2.88000000 0.24000000 ;
     RECT 0.55500000 0.42000000 0.88500000 0.75000000 ;
     RECT 1.75500000 0.42000000 2.08500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 0.55500000 2.17500000 0.88500000 2.50500000 ;
     RECT 1.75500000 2.71500000 2.08500000 3.04500000 ;
     RECT 0.00000000 3.09000000 2.88000000 3.57000000 ;

    LAYER viali ;
     RECT 1.83500000 -0.08500000 2.00500000 0.08500000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 1.83500000 0.50000000 2.00500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 1.83500000 2.79500000 2.00500000 2.96500000 ;
     RECT 1.83500000 3.24500000 2.00500000 3.41500000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 2.88000000 0.24000000 ;
     RECT 1.85000000 0.24000000 1.99000000 0.44000000 ;
     RECT 1.77500000 0.44000000 2.06500000 0.73000000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
     RECT 0.57500000 0.44000000 0.86500000 0.73000000 ;
     RECT 0.65000000 0.73000000 0.79000000 2.19500000 ;
     RECT 0.57500000 2.19500000 0.86500000 2.48500000 ;
     RECT 1.77500000 2.73500000 2.06500000 3.09000000 ;
     RECT 0.00000000 3.09000000 2.88000000 3.57000000 ;

 END
END INV
