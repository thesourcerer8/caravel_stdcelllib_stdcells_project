MACRO HAX1
 CLASS CORE ;
 FOREIGN HAX1 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 15.84000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 15.84000000 0.24000000 ;
    END
  END GND

  PIN YS
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 14.73500000 0.39500000 15.02500000 0.68500000 ;
        RECT 14.81000000 0.68500000 14.95000000 2.15000000 ;
        RECT 14.73500000 2.15000000 15.02500000 2.44000000 ;
    END
  END YS

  PIN YC
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.77500000 0.39500000 2.06500000 0.47000000 ;
        RECT 0.89000000 0.47000000 2.06500000 0.61000000 ;
        RECT 1.77500000 0.61000000 2.06500000 0.68500000 ;
        RECT 0.89000000 0.61000000 1.03000000 2.22500000 ;
        RECT 1.77500000 2.15000000 2.06500000 2.22500000 ;
        RECT 0.89000000 2.22500000 2.06500000 2.36500000 ;
        RECT 1.77500000 2.36500000 2.06500000 2.44000000 ;
    END
  END YC

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 4.25000000 0.47000000 9.19000000 0.53000000 ;
        RECT 4.25000000 0.53000000 9.26500000 0.61000000 ;
        RECT 4.25000000 0.61000000 4.39000000 0.80000000 ;
        RECT 8.97500000 0.61000000 9.26500000 0.82000000 ;
        RECT 4.17500000 0.80000000 4.46500000 1.09000000 ;
        RECT 4.25000000 1.09000000 4.39000000 1.74500000 ;
        RECT 4.17500000 1.74500000 4.46500000 2.03500000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 5.61500000 0.80000000 5.90500000 1.01000000 ;
        RECT 11.37500000 0.80000000 11.66500000 1.01000000 ;
        RECT 5.61500000 1.01000000 11.66500000 1.09000000 ;
        RECT 5.69000000 1.09000000 11.59000000 1.15000000 ;
        RECT 5.69000000 1.15000000 5.83000000 1.74500000 ;
        RECT 11.45000000 1.15000000 11.59000000 1.74500000 ;
        RECT 5.61500000 1.74500000 5.90500000 2.03500000 ;
        RECT 11.37500000 1.74500000 11.66500000 2.03500000 ;
    END
  END A


END HAX1
