magic
tech sky130A
timestamp 1621277438
<< end >>
