magic
tech sky130A
magscale 1 2
timestamp 1636962388
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1152 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 451 134 509 146
rect 451 132 463 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 463 132
rect 497 132 509 134
rect 643 134 701 146
rect 643 132 655 134
rect 497 100 561 132
rect 303 48 561 100
rect 591 100 655 132
rect 689 132 701 134
rect 931 134 989 146
rect 931 132 943 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 977 100 1037 132
rect 879 48 1037 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 175 485
rect 209 451 273 485
rect 115 450 273 451
rect 303 450 561 618
rect 591 593 849 618
rect 591 559 655 593
rect 689 559 849 593
rect 591 450 849 559
rect 879 485 1037 618
rect 879 451 943 485
rect 977 451 1037 485
rect 879 450 1037 451
rect 163 439 221 450
rect 931 439 989 450
<< ndiffc >>
rect 127 100 161 134
rect 463 100 497 134
rect 655 100 689 134
rect 943 100 977 134
<< pdiffc >>
rect 175 451 209 485
rect 655 559 689 593
rect 943 451 977 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1152 683
rect 31 618 1121 649
rect 639 593 705 618
rect 639 559 655 593
rect 689 559 705 593
rect 639 543 705 559
rect 159 485 225 501
rect 159 451 175 485
rect 209 452 225 485
rect 927 485 993 501
rect 209 451 221 452
rect 159 435 221 451
rect 927 451 943 485
rect 977 451 993 485
rect 927 435 993 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 893 418
rect 831 368 847 402
rect 881 401 893 402
rect 881 368 897 401
rect 831 352 897 368
rect 271 231 305 352
rect 559 231 593 262
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 543 215 609 231
rect 543 184 559 215
rect 255 165 321 181
rect 547 181 559 184
rect 593 181 609 215
rect 547 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 881 181 893 184
rect 831 165 893 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 447 134 513 150
rect 447 100 463 134
rect 497 100 513 134
rect 643 134 705 150
rect 643 131 655 134
rect 447 84 513 100
rect 639 100 655 131
rect 689 100 705 134
rect 639 84 705 100
rect 927 134 993 150
rect 927 100 943 134
rect 977 100 993 134
rect 927 84 993 100
rect 31 17 1121 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1152 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 655 559 689 593
rect 175 451 209 485
rect 943 451 977 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 559 262 593 296
rect 847 181 881 215
rect 127 100 161 134
rect 463 100 497 134
rect 655 100 689 134
rect 943 100 977 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1152 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1152 683
rect 0 618 1152 649
rect 643 593 701 618
rect 643 559 655 593
rect 689 559 701 593
rect 643 547 701 559
rect 163 485 221 497
rect 163 451 175 485
rect 209 451 221 485
rect 163 439 221 451
rect 931 485 989 497
rect 931 451 943 485
rect 977 451 989 485
rect 931 439 989 451
rect 178 212 206 439
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 562 308 590 356
rect 547 296 605 308
rect 547 262 559 296
rect 593 262 605 296
rect 547 250 605 262
rect 850 227 878 356
rect 835 215 893 227
rect 835 212 847 215
rect 178 184 847 212
rect 466 146 494 184
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 946 146 974 439
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 451 134 509 146
rect 451 100 463 134
rect 497 100 509 134
rect 451 88 509 100
rect 643 134 701 146
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 931 134 989 146
rect 931 100 943 134
rect 977 100 989 134
rect 931 88 989 100
rect 130 48 158 88
rect 658 48 686 88
rect 0 17 1152 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1152 17
rect 0 -48 1152 -17
<< labels >>
rlabel metal1 0 618 1152 714 0 VPWR
port 3 se
rlabel metal1 0 618 1152 714 0 VPWR
port 3 se
rlabel metal1 0 -48 1152 48 0 VGND
port 2 se
rlabel metal1 0 -48 1152 48 0 VGND
port 2 se
rlabel metal1 931 88 989 146 0 Y
port 4 se
rlabel metal1 946 146 974 439 0 Y
port 4 se
rlabel metal1 931 439 989 497 0 Y
port 4 se
rlabel metal1 547 250 605 308 0 B
port 1 se
rlabel metal1 562 308 590 356 0 B
port 1 se
rlabel metal1 547 356 605 414 0 B
port 1 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel locali 0 -17 1152 17 4 VGND
port 2 se ground default abutment
rlabel locali 31 17 1121 48 4 VGND
port 2 se ground default abutment
rlabel locali 0 649 1152 683 4 VPWR
port 3 se power default abutment
rlabel locali 31 618 1121 649 4 VGND
port 2 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1152 666
<< end >>
