* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_ls__decap_8 abstract view
.subckt sky130_fd_sc_ls__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_ls__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__decap_4 abstract view
.subckt sky130_fd_sc_ls__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__fill_1 abstract view
.subckt sky130_fd_sc_ls__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__fill_2 abstract view
.subckt sky130_fd_sc_ls__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__diode_2 abstract view
.subckt sky130_fd_sc_ls__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__conb_1 abstract view
.subckt sky130_fd_sc_ls__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__clkbuf_4 abstract view
.subckt sky130_fd_sc_ls__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 VPWR VGND Y B A
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 VPWR VGND Y B A
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 VPWR VGND Y C B A
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 VPWR VGND Y A B
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 VPWR VGND Y A
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 VPWR VGND Y A
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 VPWR VGND Y B A
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 VPWR VGND Y A
.ends

* Black-box entry subcircuit for OR2X1 abstract view
.subckt OR2X1 VPWR VGND Y B A
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 VPWR VGND Y A B
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 VPWR VGND Y A
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 VPWR VGND Y C B D A
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__clkbuf_2 abstract view
.subckt sky130_fd_sc_ls__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 VPWR VGND Y A
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__buf_2 abstract view
.subckt sky130_fd_sc_ls__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 VPWR VGND Y B A C
.ends

* Black-box entry subcircuit for INV abstract view
.subckt INV VPWR VGND Y A
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 VPWR VGND Y A
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__buf_1 abstract view
.subckt sky130_fd_sc_ls__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__buf_4 abstract view
.subckt sky130_fd_sc_ls__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 VPWR VGND Y B A D C
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 VPWR VGND Y A
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 VPWR VGND Y B S A
.ends

* Black-box entry subcircuit for AND2X1 abstract view
.subckt AND2X1 VPWR VGND Y B A
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 VPWR VGND Y B A
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 VPWR VGND Y C A B
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_188 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output56_A NAND2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AND2X2_A AND2X2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_38_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_OAI22X1_A input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_200_ vssd1 vssd1 vccd1 vccd1 _200_/HI wbs_dat_o[17] sky130_fd_sc_ls__conb_1
XFILLER_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_131_ vssd1 vssd1 vccd1 vccd1 _131_/HI la_data_out[77] sky130_fd_sc_ls__conb_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_062_ vssd1 vssd1 vccd1 vccd1 _062_/HI la_data_out[0] sky130_fd_sc_ls__conb_1
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_9_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_114_ vssd1 vssd1 vccd1 vccd1 _114_/HI la_data_out[60] sky130_fd_sc_ls__conb_1
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_045_ vssd1 vssd1 vccd1 vccd1 _045_/HI io_out[13] sky130_fd_sc_ls__conb_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_507 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input18_A io_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_028_ vssd1 vssd1 vccd1 vccd1 _028_/HI io_oeb[22] sky130_fd_sc_ls__conb_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_326 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_20_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_871 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_893 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput53 AND2X1/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_ls__clkbuf_4
Xoutput64 XOR2X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_ls__clkbuf_4
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_189 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output49_A INV/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XNAND2X1 vccd1 vssd1 NAND2X1/Y input19/X input18/X NAND2X1
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AND2X2_B AND2X2/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OAI22X1_B input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_130_ vssd1 vssd1 vccd1 vccd1 _130_/HI la_data_out[76] sky130_fd_sc_ls__conb_1
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_061_ vssd1 vssd1 vccd1 vccd1 _061_/HI irq[2] sky130_fd_sc_ls__conb_1
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_113_ vssd1 vssd1 vccd1 vccd1 _113_/HI la_data_out[59] sky130_fd_sc_ls__conb_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_044_ vssd1 vssd1 vccd1 vccd1 _044_/HI io_out[12] sky130_fd_sc_ls__conb_1
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_027_ vssd1 vssd1 vccd1 vccd1 _027_/HI io_oeb[20] sky130_fd_sc_ls__conb_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_316 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_13_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_850 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INVX1_A INVX1/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
Xoutput54 INVX8/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_ls__clkbuf_4
Xoutput65 NAND3X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_ls__clkbuf_4
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input30_A la_data_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_168 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI21X1_Y AOI21X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output61_A OR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_OAI22X1_C input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_060_ vssd1 vssd1 vccd1 vccd1 _060_/HI irq[1] sky130_fd_sc_ls__conb_1
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_189_ vssd1 vssd1 vccd1 vccd1 _189_/HI wbs_dat_o[6] sky130_fd_sc_ls__conb_1
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_112_ vssd1 vssd1 vccd1 vccd1 _112_/HI la_data_out[58] sky130_fd_sc_ls__conb_1
X_043_ vssd1 vssd1 vccd1 vccd1 _043_/HI io_out[11] sky130_fd_sc_ls__conb_1
XFILLER_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_026_ vssd1 vssd1 vccd1 vccd1 _026_/HI io_oeb[18] sky130_fd_sc_ls__conb_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_328 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput55 MUX2X1/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_ls__clkbuf_4
Xoutput66 NOR2X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_ls__clkbuf_4
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input23_A io_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_009_ vssd1 vssd1 vccd1 vccd1 io_oeb[27] _009_/LO sky130_fd_sc_ls__conb_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_BUFX4_Y BUFX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INVX4_Y INVX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_72_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI22X1_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output54_A INVX8/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_OAI22X1_D input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_188_ vssd1 vssd1 vccd1 vccd1 _188_/HI wbs_dat_o[5] sky130_fd_sc_ls__conb_1
XFILLER_36_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_111_ vssd1 vssd1 vccd1 vccd1 _111_/HI la_data_out[57] sky130_fd_sc_ls__conb_1
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_042_ vssd1 vssd1 vccd1 vccd1 _042_/HI io_out[10] sky130_fd_sc_ls__conb_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_30_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_025_ vssd1 vssd1 vccd1 vccd1 _025_/HI io_oeb[16] sky130_fd_sc_ls__conb_1
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_318 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_852 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_OR2X2_A OR2X2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput45 AOI22X1/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_ls__clkbuf_4
Xoutput56 NAND2X1/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_ls__clkbuf_4
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input16_A io_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_008_ vssd1 vssd1 vccd1 vccd1 io_oeb[25] _008_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input8_A io_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_671 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XXNOR2X1 vccd1 vssd1 XNOR2X1/Y input36/X input35/X XNOR2X1
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI22X1_B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_output47_A BUFX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_187_ vssd1 vssd1 vccd1 vccd1 _187_/HI wbs_dat_o[4] sky130_fd_sc_ls__conb_1
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_110_ vssd1 vssd1 vccd1 vccd1 _110_/HI la_data_out[56] sky130_fd_sc_ls__conb_1
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_041_ vssd1 vssd1 vccd1 vccd1 _041_/HI io_out[8] sky130_fd_sc_ls__conb_1
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_024_ vssd1 vssd1 vccd1 vccd1 _024_/HI io_oeb[14] sky130_fd_sc_ls__conb_1
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_853 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OR2X2_B OR2X2/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput46 BUFX2/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_ls__clkbuf_4
Xoutput57 AND2X2/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_ls__clkbuf_4
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_007_ vssd1 vssd1 vccd1 vccd1 io_oeb[23] _007_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI22X1_C input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XAOI21X1 vccd1 vssd1 AOI21X1/Y input24/X input23/X input22/X AOI21X1
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_37_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_186_ vssd1 vssd1 vccd1 vccd1 _186_/HI wbs_dat_o[3] sky130_fd_sc_ls__conb_1
XFILLER_6_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_040_ vssd1 vssd1 vccd1 vccd1 _040_/HI io_out[7] sky130_fd_sc_ls__conb_1
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input39_A la_data_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_169_ vssd1 vssd1 vccd1 vccd1 _169_/HI la_data_out[115] sky130_fd_sc_ls__conb_1
XFILLER_41_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_023_ vssd1 vssd1 vccd1 vccd1 io_oeb[10] _023_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XXOR2X1 vccd1 vssd1 XOR2X1/Y XOR2X1/A XOR2X1/B XOR2X1
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1081 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput58 AOI21X1/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_ls__clkbuf_4
Xoutput47 BUFX4/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_ls__clkbuf_4
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_006_ vssd1 vssd1 vccd1 vccd1 io_oeb[21] _006_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_640 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input21_A io_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_8_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XANTENNA_AOI22X1_D input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_BUFX2_Y BUFX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_INVX2_Y INVX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_185_ vssd1 vssd1 vccd1 vccd1 _185_/HI wbs_dat_o[2] sky130_fd_sc_ls__conb_1
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INV_A INV/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_output52_A INVX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_NOR2X1_Y NOR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_CLKBUF1_A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_51_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_168_ vssd1 vssd1 vccd1 vccd1 _168_/HI la_data_out[114] sky130_fd_sc_ls__conb_1
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_099_ vssd1 vssd1 vccd1 vccd1 _099_/HI la_data_out[45] sky130_fd_sc_ls__conb_1
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_022_ vssd1 vssd1 vccd1 vccd1 io_oeb[8] _022_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1082 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput48 CLKBUF1/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_ls__clkbuf_4
Xoutput59 OAI21X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_ls__clkbuf_4
XFILLER_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_005_ vssd1 vssd1 vccd1 vccd1 io_oeb[19] _005_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input14_A io_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_NAND2X1_Y NAND2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input6_A io_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XINVX1 vccd1 vssd1 INVX1/Y INVX1/A INVX1
XTAP_290 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_184_ vssd1 vssd1 vccd1 vccd1 _184_/HI wbs_dat_o[1] sky130_fd_sc_ls__conb_1
XFILLER_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_output45_A AOI22X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_167_ vssd1 vssd1 vccd1 vccd1 _167_/HI la_data_out[113] sky130_fd_sc_ls__conb_1
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_098_ vssd1 vssd1 vccd1 vccd1 _098_/HI la_data_out[44] sky130_fd_sc_ls__conb_1
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_021_ vssd1 vssd1 vccd1 vccd1 io_oeb[7] _021_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input44_A la_data_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XANTENNA_AND2X1_Y AND2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_80_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput49 INV/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_ls__clkbuf_4
XFILLER_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_72_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_004_ vssd1 vssd1 vccd1 vccd1 io_oeb[17] _004_/LO sky130_fd_sc_ls__conb_1
XFILLER_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_697 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_NAND3X1_A input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_450 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_461 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XINVX2 vccd1 vssd1 INVX2/Y INVX2/A INVX2
XFILLER_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_183_ vssd1 vssd1 vccd1 vccd1 _183_/HI wbs_dat_o[0] sky130_fd_sc_ls__conb_1
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_166_ vssd1 vssd1 vccd1 vccd1 _166_/HI la_data_out[112] sky130_fd_sc_ls__conb_1
X_097_ vssd1 vssd1 vccd1 vccd1 _097_/HI la_data_out[43] sky130_fd_sc_ls__conb_1
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_020_ vssd1 vssd1 vccd1 vccd1 io_oeb[6] _020_/LO sky130_fd_sc_ls__conb_1
XFILLER_20_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INVX8_A INVX8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input37_A la_data_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1073 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_149_ vssd1 vssd1 vccd1 vccd1 _149_/HI la_data_out[95] sky130_fd_sc_ls__conb_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XNOR2X1 vccd1 vssd1 NOR2X1/Y NOR2X1/B NOR2X1/A NOR2X1
XFILLER_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_72_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_003_ vssd1 vssd1 vccd1 vccd1 io_oeb[15] _003_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_NAND3X1_B input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_440 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_64_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_182_ vssd1 vssd1 vccd1 vccd1 _182_/HI wbs_ack_o sky130_fd_sc_ls__conb_1
XFILLER_10_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_165_ vssd1 vssd1 vccd1 vccd1 _165_/HI la_data_out[111] sky130_fd_sc_ls__conb_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_096_ vssd1 vssd1 vccd1 vccd1 _096_/HI la_data_out[42] sky130_fd_sc_ls__conb_1
XFILLER_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output50_A INVX1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_MUX2X1_A MUX2X1/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_217_ vssd1 vssd1 vccd1 vccd1 _217_/HI io_oeb[9] sky130_fd_sc_ls__conb_1
X_148_ vssd1 vssd1 vccd1 vccd1 _148_/HI la_data_out[94] sky130_fd_sc_ls__conb_1
X_079_ vssd1 vssd1 vccd1 vccd1 _079_/HI la_data_out[23] sky130_fd_sc_ls__conb_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_32_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_869 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_002_ vssd1 vssd1 vccd1 vccd1 io_oeb[13] _002_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_688 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_NAND3X1_C input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_441 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input12_A io_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input4_A io_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XINVX4 vccd1 vssd1 INVX4/Y INVX4/A INVX4
XTAP_293 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_181_ vssd1 vssd1 vccd1 vccd1 _181_/HI la_data_out[127] sky130_fd_sc_ls__conb_1
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_10_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_164_ vssd1 vssd1 vccd1 vccd1 _164_/HI la_data_out[110] sky130_fd_sc_ls__conb_1
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_095_ vssd1 vssd1 vccd1 vccd1 _095_/HI la_data_out[41] sky130_fd_sc_ls__conb_1
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_XOR2X1_A XOR2X1/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_MUX2X1_B MUX2X1/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_216_ vssd1 vssd1 vccd1 vccd1 _216_/HI io_oeb[5] sky130_fd_sc_ls__conb_1
XFILLER_51_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_147_ vssd1 vssd1 vccd1 vccd1 _147_/HI la_data_out[93] sky130_fd_sc_ls__conb_1
X_078_ vssd1 vssd1 vccd1 vccd1 _078_/HI la_data_out[22] sky130_fd_sc_ls__conb_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_001_ vssd1 vssd1 vccd1 vccd1 io_oeb[12] _001_/LO sky130_fd_sc_ls__conb_1
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input42_A la_data_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_601 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_420 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XOR2X1 vccd1 vssd1 OR2X1/Y OR2X1/B OR2X1/A OR2X1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OAI21X1_A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_48_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_283 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_294 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_OR2X1_Y OR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_180_ vssd1 vssd1 vccd1 vccd1 _180_/HI la_data_out[126] sky130_fd_sc_ls__conb_1
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_163_ vssd1 vssd1 vccd1 vccd1 _163_/HI la_data_out[109] sky130_fd_sc_ls__conb_1
X_094_ vssd1 vssd1 vccd1 vccd1 _094_/HI la_data_out[40] sky130_fd_sc_ls__conb_1
XFILLER_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_19_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_XOR2X1_B XOR2X1/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_215_ vssd1 vssd1 vccd1 vccd1 _215_/HI io_oeb[2] sky130_fd_sc_ls__conb_1
XFILLER_11_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_146_ vssd1 vssd1 vccd1 vccd1 _146_/HI la_data_out[92] sky130_fd_sc_ls__conb_1
XFILLER_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_077_ vssd1 vssd1 vccd1 vccd1 _077_/HI la_data_out[20] sky130_fd_sc_ls__conb_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_000_ vssd1 vssd1 vccd1 vccd1 io_oeb[11] _000_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input35_A la_data_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_129_ vssd1 vssd1 vccd1 vccd1 _129_/HI la_data_out[75] sky130_fd_sc_ls__conb_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XOR2X2 vccd1 vssd1 OR2X2/Y OR2X2/A OR2X2/B OR2X2
XFILLER_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output66_A NOR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OAI21X1_B input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_162_ vssd1 vssd1 vccd1 vccd1 _162_/HI la_data_out[108] sky130_fd_sc_ls__conb_1
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_093_ vssd1 vssd1 vccd1 vccd1 _093_/HI la_data_out[39] sky130_fd_sc_ls__conb_1
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_ls__clkbuf_4
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1077 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_214_ vssd1 vssd1 vccd1 vccd1 _214_/HI wbs_dat_o[31] sky130_fd_sc_ls__conb_1
XFILLER_42_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_145_ vssd1 vssd1 vccd1 vccd1 _145_/HI la_data_out[91] sky130_fd_sc_ls__conb_1
X_076_ vssd1 vssd1 vccd1 vccd1 _076_/HI la_data_out[19] sky130_fd_sc_ls__conb_1
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_839 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input28_A la_data_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_128_ vssd1 vssd1 vccd1 vccd1 _128_/HI la_data_out[74] sky130_fd_sc_ls__conb_1
X_059_ vssd1 vssd1 vccd1 vccd1 _059_/HI irq[0] sky130_fd_sc_ls__conb_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_603 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_636 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_400 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_477 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output59_A OAI21X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_OAI21X1_C input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_241 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input10_A io_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input2_A io_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_161_ vssd1 vssd1 vccd1 vccd1 _161_/HI la_data_out[107] sky130_fd_sc_ls__conb_1
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_092_ vssd1 vssd1 vccd1 vccd1 _092_/HI la_data_out[38] sky130_fd_sc_ls__conb_1
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_ls__clkbuf_4
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1078 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_213_ vssd1 vssd1 vccd1 vccd1 _213_/HI wbs_dat_o[30] sky130_fd_sc_ls__conb_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_144_ vssd1 vssd1 vccd1 vccd1 _144_/HI la_data_out[90] sky130_fd_sc_ls__conb_1
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_075_ vssd1 vssd1 vccd1 vccd1 _075_/HI la_data_out[17] sky130_fd_sc_ls__conb_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_127_ vssd1 vssd1 vccd1 vccd1 _127_/HI la_data_out[73] sky130_fd_sc_ls__conb_1
XFILLER_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_058_ vssd1 vssd1 vccd1 vccd1 _058_/HI io_out[36] sky130_fd_sc_ls__conb_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input40_A la_data_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_401 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_445 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_AOI21X1_A input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_78_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_990 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_242 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XINVX8 vccd1 vssd1 INVX8/Y INVX8/A INVX8
XTAP_297 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_160_ vssd1 vssd1 vccd1 vccd1 _160_/HI la_data_out[106] sky130_fd_sc_ls__conb_1
XFILLER_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_091_ vssd1 vssd1 vccd1 vccd1 _091_/HI la_data_out[37] sky130_fd_sc_ls__conb_1
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_ls__clkbuf_4
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_212_ vssd1 vssd1 vccd1 vccd1 _212_/HI wbs_dat_o[29] sky130_fd_sc_ls__conb_1
XFILLER_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_143_ vssd1 vssd1 vccd1 vccd1 _143_/HI la_data_out[89] sky130_fd_sc_ls__conb_1
XFILLER_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_074_ vssd1 vssd1 vccd1 vccd1 _074_/HI la_data_out[16] sky130_fd_sc_ls__conb_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_126_ vssd1 vssd1 vccd1 vccd1 _126_/HI la_data_out[72] sky130_fd_sc_ls__conb_1
XFILLER_11_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_057_ vssd1 vssd1 vccd1 vccd1 _057_/HI io_out[35] sky130_fd_sc_ls__conb_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_BUFX4_A BUFX4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INVX4_A INVX4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XANTENNA_input33_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XOAI22X1 vccd1 vssd1 OAI22X1/Y input28/X input27/X input29/X input26/X OAI22X1
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_109_ vssd1 vssd1 vccd1 vccd1 _109_/HI la_data_out[55] sky130_fd_sc_ls__conb_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI21X1_B input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_232 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output64_A XOR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_76_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_090_ vssd1 vssd1 vccd1 vccd1 _090_/HI la_data_out[36] sky130_fd_sc_ls__conb_1
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_ls__clkbuf_4
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1069 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_211_ vssd1 vssd1 vccd1 vccd1 _211_/HI wbs_dat_o[28] sky130_fd_sc_ls__conb_1
XFILLER_11_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_142_ vssd1 vssd1 vccd1 vccd1 _142_/HI la_data_out[88] sky130_fd_sc_ls__conb_1
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_073_ vssd1 vssd1 vccd1 vccd1 _073_/HI la_data_out[14] sky130_fd_sc_ls__conb_1
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_809 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_125_ vssd1 vssd1 vccd1 vccd1 _125_/HI la_data_out[71] sky130_fd_sc_ls__conb_1
X_056_ vssd1 vssd1 vccd1 vccd1 _056_/HI io_out[33] sky130_fd_sc_ls__conb_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_606 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput40 la_data_in[4] vssd1 vssd1 vccd1 vccd1 NOR2X1/A sky130_fd_sc_ls__clkbuf_2
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input26_A la_data_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_108_ vssd1 vssd1 vccd1 vccd1 _108_/HI la_data_out[54] sky130_fd_sc_ls__conb_1
X_039_ vssd1 vssd1 vccd1 vccd1 _039_/HI io_out[6] sky130_fd_sc_ls__conb_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI21X1_C input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_992 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_233 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output57_A AND2X2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_ls__clkbuf_4
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XBUFX2 vccd1 vssd1 BUFX2/Y BUFX2/A BUFX2
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1026 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_210_ vssd1 vssd1 vccd1 vccd1 _210_/HI wbs_dat_o[27] sky130_fd_sc_ls__conb_1
X_141_ vssd1 vssd1 vccd1 vccd1 _141_/HI la_data_out[87] sky130_fd_sc_ls__conb_1
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_072_ vssd1 vssd1 vccd1 vccd1 _072_/HI la_data_out[13] sky130_fd_sc_ls__conb_1
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_124_ vssd1 vssd1 vccd1 vccd1 _124_/HI la_data_out[70] sky130_fd_sc_ls__conb_1
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_055_ vssd1 vssd1 vccd1 vccd1 _055_/HI io_out[32] sky130_fd_sc_ls__conb_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput30 la_data_in[16] vssd1 vssd1 vccd1 vccd1 OR2X1/A sky130_fd_sc_ls__buf_2
Xinput41 la_data_in[5] vssd1 vssd1 vccd1 vccd1 NOR2X1/B sky130_fd_sc_ls__clkbuf_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_input19_A io_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_107_ vssd1 vssd1 vccd1 vccd1 _107_/HI la_data_out[53] sky130_fd_sc_ls__conb_1
XFILLER_7_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_038_ vssd1 vssd1 vccd1 vccd1 _038_/HI io_out[4] sky130_fd_sc_ls__conb_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_21_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_459 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_54_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_223 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_256 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_790 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XNAND3X1 vccd1 vssd1 NAND3X1/Y input33/X input25/X input39/X NAND3X1
XFILLER_14_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput6 io_in[15] vssd1 vssd1 vccd1 vccd1 BUFX2/A sky130_fd_sc_ls__clkbuf_4
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_140_ vssd1 vssd1 vccd1 vccd1 _140_/HI la_data_out[86] sky130_fd_sc_ls__conb_1
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_071_ vssd1 vssd1 vccd1 vccd1 _071_/HI la_data_out[12] sky130_fd_sc_ls__conb_1
XFILLER_2_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XINV vccd1 vssd1 INV/Y INV/A INV
XFILLER_20_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_123_ vssd1 vssd1 vccd1 vccd1 _123_/HI la_data_out[69] sky130_fd_sc_ls__conb_1
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_054_ vssd1 vssd1 vccd1 vccd1 _054_/HI io_out[31] sky130_fd_sc_ls__conb_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput20 io_in[3] vssd1 vssd1 vccd1 vccd1 AND2X2/A sky130_fd_sc_ls__clkbuf_4
Xinput31 la_data_in[17] vssd1 vssd1 vccd1 vccd1 OR2X1/B sky130_fd_sc_ls__buf_2
Xinput42 la_data_in[7] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_ls__clkbuf_2
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_106_ vssd1 vssd1 vccd1 vccd1 _106_/HI la_data_out[52] sky130_fd_sc_ls__conb_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_037_ vssd1 vssd1 vccd1 vccd1 _037_/HI io_out[3] sky130_fd_sc_ls__conb_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_961 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XANTENNA_BUFX2_A BUFX2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INVX2_A INVX2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input31_A la_data_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_224 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_202 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_780 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_NOR2X1_A NOR2X1/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_output62_A OR2X2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput7 io_in[17] vssd1 vssd1 vccd1 vccd1 BUFX4/A sky130_fd_sc_ls__clkbuf_4
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XBUFX4 vccd1 vssd1 BUFX4/Y BUFX4/A BUFX4
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1028 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1039 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_070_ vssd1 vssd1 vccd1 vccd1 _070_/HI la_data_out[11] sky130_fd_sc_ls__conb_1
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_199_ vssd1 vssd1 vccd1 vccd1 _199_/HI wbs_dat_o[16] sky130_fd_sc_ls__conb_1
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_122_ vssd1 vssd1 vccd1 vccd1 _122_/HI la_data_out[68] sky130_fd_sc_ls__conb_1
X_053_ vssd1 vssd1 vccd1 vccd1 _053_/HI io_out[29] sky130_fd_sc_ls__conb_1
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput10 io_in[21] vssd1 vssd1 vccd1 vccd1 INV/A sky130_fd_sc_ls__clkbuf_4
Xinput21 io_in[4] vssd1 vssd1 vccd1 vccd1 AND2X2/B sky130_fd_sc_ls__clkbuf_4
Xinput43 la_data_in[8] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_ls__clkbuf_2
Xinput32 la_data_in[19] vssd1 vssd1 vccd1 vccd1 OR2X2/A sky130_fd_sc_ls__buf_2
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_105_ vssd1 vssd1 vccd1 vccd1 _105_/HI la_data_out[51] sky130_fd_sc_ls__conb_1
X_036_ vssd1 vssd1 vccd1 vccd1 _036_/HI io_out[1] sky130_fd_sc_ls__conb_1
XANTENNA_NAND2X1_A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_995 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input24_A io_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_8_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_019_ vssd1 vssd1 vccd1 vccd1 io_oeb[4] _019_/LO sky130_fd_sc_ls__conb_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_770 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_781 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_NOR2X1_B NOR2X1/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput8 io_in[19] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_ls__clkbuf_4
XANTENNA_output55_A MUX2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_198_ vssd1 vssd1 vccd1 vccd1 _198_/HI wbs_dat_o[15] sky130_fd_sc_ls__conb_1
XFILLER_10_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_AND2X1_A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_37_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_121_ vssd1 vssd1 vccd1 vccd1 _121_/HI la_data_out[67] sky130_fd_sc_ls__conb_1
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_052_ vssd1 vssd1 vccd1 vccd1 _052_/HI io_out[27] sky130_fd_sc_ls__conb_1
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput11 io_in[23] vssd1 vssd1 vccd1 vccd1 INVX1/A sky130_fd_sc_ls__clkbuf_4
Xinput22 io_in[6] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_ls__buf_2
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput44 la_data_in[9] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_ls__clkbuf_2
Xinput33 la_data_in[1] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_ls__buf_1
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_16_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_104_ vssd1 vssd1 vccd1 vccd1 _104_/HI la_data_out[50] sky130_fd_sc_ls__conb_1
X_035_ vssd1 vssd1 vccd1 vccd1 _035_/HI io_out[0] sky130_fd_sc_ls__conb_1
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_NAND2X1_B input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_407 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_941 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input17_A io_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_018_ vssd1 vssd1 vccd1 vccd1 io_oeb[3] _018_/LO sky130_fd_sc_ls__conb_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_259 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input9_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_26_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output48_A CLKBUF1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
Xinput9 io_in[1] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_ls__clkbuf_4
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1019 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_197_ vssd1 vssd1 vccd1 vccd1 _197_/HI wbs_dat_o[14] sky130_fd_sc_ls__conb_1
XANTENNA_AND2X1_B input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_120_ vssd1 vssd1 vccd1 vccd1 _120_/HI la_data_out[66] sky130_fd_sc_ls__conb_1
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_051_ vssd1 vssd1 vccd1 vccd1 _051_/HI io_out[25] sky130_fd_sc_ls__conb_1
XFILLER_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput12 io_in[25] vssd1 vssd1 vccd1 vccd1 INVX2/A sky130_fd_sc_ls__buf_4
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput23 io_in[7] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_ls__clkbuf_4
Xinput34 la_data_in[20] vssd1 vssd1 vccd1 vccd1 OR2X2/B sky130_fd_sc_ls__buf_2
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_32_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_103_ vssd1 vssd1 vccd1 vccd1 _103_/HI la_data_out[49] sky130_fd_sc_ls__conb_1
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_034_ vssd1 vssd1 vccd1 vccd1 _034_/HI io_oeb[37] sky130_fd_sc_ls__conb_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_942 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_017_ vssd1 vssd1 vccd1 vccd1 io_oeb[1] _017_/LO sky130_fd_sc_ls__conb_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_238 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_750 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XAOI22X1 vccd1 vssd1 AOI22X1/Y input3/X input2/X input5/X input4/X AOI22X1
XFILLER_40_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_XNOR2X1_Y XNOR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_196_ vssd1 vssd1 vccd1 vccd1 _196_/HI wbs_dat_o[13] sky130_fd_sc_ls__conb_1
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_output60_A OAI22X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_050_ vssd1 vssd1 vccd1 vccd1 _050_/HI io_out[23] sky130_fd_sc_ls__conb_1
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_3_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput13 io_in[27] vssd1 vssd1 vccd1 vccd1 INVX4/A sky130_fd_sc_ls__buf_4
Xinput24 io_in[8] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_ls__clkbuf_4
Xinput35 la_data_in[22] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_ls__buf_2
X_179_ vssd1 vssd1 vccd1 vccd1 _179_/HI la_data_out[125] sky130_fd_sc_ls__conb_1
XFILLER_42_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_102_ vssd1 vssd1 vccd1 vccd1 _102_/HI la_data_out[48] sky130_fd_sc_ls__conb_1
X_033_ vssd1 vssd1 vccd1 vccd1 _033_/HI io_oeb[34] sky130_fd_sc_ls__conb_1
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_932 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_016_ vssd1 vssd1 vccd1 vccd1 io_oeb[0] _016_/LO sky130_fd_sc_ls__conb_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_762 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input22_A io_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_570 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_65_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_195_ vssd1 vssd1 vccd1 vccd1 _195_/HI wbs_dat_o[12] sky130_fd_sc_ls__conb_1
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output53_A AND2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput14 io_in[29] vssd1 vssd1 vccd1 vccd1 INVX8/A sky130_fd_sc_ls__buf_4
Xinput25 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_ls__buf_1
Xinput36 la_data_in[23] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_ls__buf_2
X_178_ vssd1 vssd1 vccd1 vccd1 _178_/HI la_data_out[124] sky130_fd_sc_ls__conb_1
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_101_ vssd1 vssd1 vccd1 vccd1 _101_/HI la_data_out[47] sky130_fd_sc_ls__conb_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_032_ vssd1 vssd1 vccd1 vccd1 _032_/HI io_oeb[30] sky130_fd_sc_ls__conb_1
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_900 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_015_ vssd1 vssd1 vccd1 vccd1 io_oeb[36] _015_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_OR2X1_A OR2X1/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input15_A io_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_63_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input7_A io_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_194_ vssd1 vssd1 vccd1 vccd1 _194_/HI wbs_dat_o[11] sky130_fd_sc_ls__conb_1
XFILLER_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_output46_A BUFX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_32_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput15 io_in[31] vssd1 vssd1 vccd1 vccd1 MUX2X1/A sky130_fd_sc_ls__buf_4
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput26 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_ls__clkbuf_2
Xinput37 la_data_in[25] vssd1 vssd1 vccd1 vccd1 XOR2X1/A sky130_fd_sc_ls__buf_2
X_177_ vssd1 vssd1 vccd1 vccd1 _177_/HI la_data_out[123] sky130_fd_sc_ls__conb_1
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_100_ vssd1 vssd1 vccd1 vccd1 _100_/HI la_data_out[46] sky130_fd_sc_ls__conb_1
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_031_ vssd1 vssd1 vccd1 vccd1 _031_/HI io_oeb[28] sky130_fd_sc_ls__conb_1
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AND2X2_Y AND2X2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_945 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OAI22X1_Y OAI22X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_014_ vssd1 vssd1 vccd1 vccd1 io_oeb[35] _014_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_219 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OR2X1_B OR2X1/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_380 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_193_ vssd1 vssd1 vccd1 vccd1 _193_/HI wbs_dat_o[10] sky130_fd_sc_ls__conb_1
XFILLER_41_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput16 io_in[32] vssd1 vssd1 vccd1 vccd1 MUX2X1/B sky130_fd_sc_ls__buf_4
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput27 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_ls__clkbuf_2
X_176_ vssd1 vssd1 vccd1 vccd1 _176_/HI la_data_out[122] sky130_fd_sc_ls__conb_1
Xinput38 la_data_in[26] vssd1 vssd1 vccd1 vccd1 XOR2X1/B sky130_fd_sc_ls__buf_2
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_030_ vssd1 vssd1 vccd1 vccd1 _030_/HI io_oeb[26] sky130_fd_sc_ls__conb_1
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input38_A la_data_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_159_ vssd1 vssd1 vccd1 vccd1 _159_/HI la_data_out[105] sky130_fd_sc_ls__conb_1
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_935 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_013_ vssd1 vssd1 vccd1 vccd1 io_oeb[33] _013_/LO sky130_fd_sc_ls__conb_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_34_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input20_A io_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_192_ vssd1 vssd1 vccd1 vccd1 _192_/HI wbs_dat_o[9] sky130_fd_sc_ls__conb_1
XFILLER_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_INVX1_Y INVX1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput17 io_in[33] vssd1 vssd1 vccd1 vccd1 MUX2X1/S sky130_fd_sc_ls__buf_4
Xinput28 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_ls__clkbuf_2
XFILLER_10_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput39 la_data_in[2] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_ls__buf_1
X_175_ vssd1 vssd1 vccd1 vccd1 _175_/HI la_data_out[121] sky130_fd_sc_ls__conb_1
XFILLER_6_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output51_A INVX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XCLKBUF1 vccd1 vssd1 CLKBUF1/Y input8/X CLKBUF1
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_158_ vssd1 vssd1 vccd1 vccd1 _158_/HI la_data_out[104] sky130_fd_sc_ls__conb_1
X_089_ vssd1 vssd1 vccd1 vccd1 _089_/HI la_data_out[35] sky130_fd_sc_ls__conb_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_33_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_969 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_012_ vssd1 vssd1 vccd1 vccd1 io_oeb[32] _012_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_700 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_563 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input13_A io_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input5_A io_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_191_ vssd1 vssd1 vccd1 vccd1 _191_/HI wbs_dat_o[8] sky130_fd_sc_ls__conb_1
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput18 io_in[35] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_ls__buf_4
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput29 la_data_in[14] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_ls__clkbuf_2
X_174_ vssd1 vssd1 vccd1 vccd1 _174_/HI la_data_out[120] sky130_fd_sc_ls__conb_1
XFILLER_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XMUX2X1 vccd1 vssd1 MUX2X1/Y MUX2X1/B MUX2X1/S MUX2X1/A MUX2X1
XFILLER_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_AOI22X1_Y AOI22X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_24_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_42_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_157_ vssd1 vssd1 vccd1 vccd1 _157_/HI la_data_out[103] sky130_fd_sc_ls__conb_1
X_088_ vssd1 vssd1 vccd1 vccd1 _088_/HI la_data_out[34] sky130_fd_sc_ls__conb_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_011_ vssd1 vssd1 vccd1 vccd1 io_oeb[31] _011_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_input43_A la_data_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_209_ vssd1 vssd1 vccd1 vccd1 _209_/HI wbs_dat_o[26] sky130_fd_sc_ls__conb_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_778 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_520 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_MUX2X1_S MUX2X1/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OR2X2_Y OR2X2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_190_ vssd1 vssd1 vccd1 vccd1 _190_/HI wbs_dat_o[7] sky130_fd_sc_ls__conb_1
XFILLER_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_191 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput19 io_in[36] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_ls__buf_4
X_173_ vssd1 vssd1 vccd1 vccd1 _173_/HI la_data_out[119] sky130_fd_sc_ls__conb_1
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_156_ vssd1 vssd1 vccd1 vccd1 _156_/HI la_data_out[102] sky130_fd_sc_ls__conb_1
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_087_ vssd1 vssd1 vccd1 vccd1 _087_/HI la_data_out[33] sky130_fd_sc_ls__conb_1
XFILLER_6_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_010_ vssd1 vssd1 vccd1 vccd1 io_oeb[29] _010_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_input36_A la_data_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_208_ vssd1 vssd1 vccd1 vccd1 _208_/HI wbs_dat_o[25] sky130_fd_sc_ls__conb_1
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_139_ vssd1 vssd1 vccd1 vccd1 _139_/HI la_data_out[85] sky130_fd_sc_ls__conb_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_779 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_510 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_351 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_170 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_172_ vssd1 vssd1 vccd1 vccd1 _172_/HI la_data_out[118] sky130_fd_sc_ls__conb_1
XFILLER_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_77_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XAND2X1 vccd1 vssd1 AND2X1/Y input9/X input1/X AND2X1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_155_ vssd1 vssd1 vccd1 vccd1 _155_/HI la_data_out[101] sky130_fd_sc_ls__conb_1
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_086_ vssd1 vssd1 vccd1 vccd1 _086_/HI la_data_out[32] sky130_fd_sc_ls__conb_1
XFILLER_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input29_A la_data_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_207_ vssd1 vssd1 vccd1 vccd1 _207_/HI wbs_dat_o[24] sky130_fd_sc_ls__conb_1
X_138_ vssd1 vssd1 vccd1 vccd1 _138_/HI la_data_out[84] sky130_fd_sc_ls__conb_1
X_069_ vssd1 vssd1 vccd1 vccd1 _069_/HI la_data_out[9] sky130_fd_sc_ls__conb_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_736 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_769 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_500 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_577 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_38_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_330 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input11_A io_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_31_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input3_A io_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_171 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_171_ vssd1 vssd1 vccd1 vccd1 _171_/HI la_data_out[117] sky130_fd_sc_ls__conb_1
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_77_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XAND2X2 vccd1 vssd1 AND2X2/Y AND2X2/B AND2X2/A AND2X2
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_154_ vssd1 vssd1 vccd1 vccd1 _154_/HI la_data_out[100] sky130_fd_sc_ls__conb_1
X_085_ vssd1 vssd1 vccd1 vccd1 _085_/HI la_data_out[31] sky130_fd_sc_ls__conb_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_206_ vssd1 vssd1 vccd1 vccd1 _206_/HI wbs_dat_o[23] sky130_fd_sc_ls__conb_1
X_137_ vssd1 vssd1 vccd1 vccd1 _137_/HI la_data_out[83] sky130_fd_sc_ls__conb_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_068_ vssd1 vssd1 vccd1 vccd1 _068_/HI la_data_out[8] sky130_fd_sc_ls__conb_1
XANTENNA_INV_Y INV/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_CLKBUF1_Y CLKBUF1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input41_A la_data_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_320 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_172 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_170_ vssd1 vssd1 vccd1 vccd1 _170_/HI la_data_out[116] sky130_fd_sc_ls__conb_1
XFILLER_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_153_ vssd1 vssd1 vccd1 vccd1 _153_/HI la_data_out[99] sky130_fd_sc_ls__conb_1
X_084_ vssd1 vssd1 vccd1 vccd1 _084_/HI la_data_out[30] sky130_fd_sc_ls__conb_1
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_908 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_919 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_52_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_205_ vssd1 vssd1 vccd1 vccd1 _205_/HI wbs_dat_o[22] sky130_fd_sc_ls__conb_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_136_ vssd1 vssd1 vccd1 vccd1 _136_/HI la_data_out[82] sky130_fd_sc_ls__conb_1
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_067_ vssd1 vssd1 vccd1 vccd1 _067_/HI la_data_out[7] sky130_fd_sc_ls__conb_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_60_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input34_A la_data_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_119_ vssd1 vssd1 vccd1 vccd1 _119_/HI la_data_out[65] sky130_fd_sc_ls__conb_1
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_502 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output65_A NAND3X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_173 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_18_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_NAND3X1_Y NAND3X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_47_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_22_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_152_ vssd1 vssd1 vccd1 vccd1 _152_/HI la_data_out[98] sky130_fd_sc_ls__conb_1
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_083_ vssd1 vssd1 vccd1 vccd1 _083_/HI la_data_out[29] sky130_fd_sc_ls__conb_1
XFILLER_10_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_52_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_204_ vssd1 vssd1 vccd1 vccd1 _204_/HI wbs_dat_o[21] sky130_fd_sc_ls__conb_1
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_135_ vssd1 vssd1 vccd1 vccd1 _135_/HI la_data_out[81] sky130_fd_sc_ls__conb_1
X_066_ vssd1 vssd1 vccd1 vccd1 _066_/HI la_data_out[5] sky130_fd_sc_ls__conb_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_717 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_34_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input27_A la_data_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_118_ vssd1 vssd1 vccd1 vccd1 _118_/HI la_data_out[64] sky130_fd_sc_ls__conb_1
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_049_ vssd1 vssd1 vccd1 vccd1 _049_/HI io_out[21] sky130_fd_sc_ls__conb_1
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_INVX8_Y INVX8/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput60 OAI22X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_ls__clkbuf_4
XANTENNA_output58_A AOI21X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
X_151_ vssd1 vssd1 vccd1 vccd1 _151_/HI la_data_out[97] sky130_fd_sc_ls__conb_1
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_082_ vssd1 vssd1 vccd1 vccd1 _082_/HI la_data_out[28] sky130_fd_sc_ls__conb_1
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_74_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_203_ vssd1 vssd1 vccd1 vccd1 _203_/HI wbs_dat_o[20] sky130_fd_sc_ls__conb_1
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_134_ vssd1 vssd1 vccd1 vccd1 _134_/HI la_data_out[80] sky130_fd_sc_ls__conb_1
X_065_ vssd1 vssd1 vccd1 vccd1 _065_/HI la_data_out[4] sky130_fd_sc_ls__conb_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_28_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_117_ vssd1 vssd1 vccd1 vccd1 _117_/HI la_data_out[63] sky130_fd_sc_ls__conb_1
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_048_ vssd1 vssd1 vccd1 vccd1 _048_/HI io_out[19] sky130_fd_sc_ls__conb_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_22_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_MUX2X1_Y MUX2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_XNOR2X1_A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput50 INVX1/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_ls__clkbuf_4
Xoutput61 OR2X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_ls__clkbuf_4
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_164 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_67_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_150_ vssd1 vssd1 vccd1 vccd1 _150_/HI la_data_out[96] sky130_fd_sc_ls__conb_1
XFILLER_50_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_081_ vssd1 vssd1 vccd1 vccd1 _081_/HI la_data_out[26] sky130_fd_sc_ls__conb_1
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_202_ vssd1 vssd1 vccd1 vccd1 _202_/HI wbs_dat_o[19] sky130_fd_sc_ls__conb_1
XFILLER_51_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_133_ vssd1 vssd1 vccd1 vccd1 _133_/HI la_data_out[79] sky130_fd_sc_ls__conb_1
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_064_ vssd1 vssd1 vccd1 vccd1 _064_/HI la_data_out[2] sky130_fd_sc_ls__conb_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_116_ vssd1 vssd1 vccd1 vccd1 _116_/HI la_data_out[62] sky130_fd_sc_ls__conb_1
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_047_ vssd1 vssd1 vccd1 vccd1 _047_/HI io_out[17] sky130_fd_sc_ls__conb_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input32_A la_data_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_XOR2X1_Y XOR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XOAI21X1 vccd1 vssd1 OAI21X1/Y input44/X input42/X input43/X OAI21X1
XFILLER_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_XNOR2X1_B input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XTAP_313 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput51 INVX2/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_ls__clkbuf_4
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput62 OR2X2/Y vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_ls__clkbuf_4
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_165 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_187 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_output63_A XNOR2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_080_ vssd1 vssd1 vccd1 vccd1 _080_/HI la_data_out[25] sky130_fd_sc_ls__conb_1
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_OAI21X1_Y OAI21X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_201_ vssd1 vssd1 vccd1 vccd1 _201_/HI wbs_dat_o[18] sky130_fd_sc_ls__conb_1
X_132_ vssd1 vssd1 vccd1 vccd1 _132_/HI la_data_out[78] sky130_fd_sc_ls__conb_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_063_ vssd1 vssd1 vccd1 vccd1 _063_/HI la_data_out[1] sky130_fd_sc_ls__conb_1
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_115_ vssd1 vssd1 vccd1 vccd1 _115_/HI la_data_out[61] sky130_fd_sc_ls__conb_1
X_046_ vssd1 vssd1 vccd1 vccd1 _046_/HI io_out[15] sky130_fd_sc_ls__conb_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_input25_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_48_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_029_ vssd1 vssd1 vccd1 vccd1 _029_/HI io_oeb[24] sky130_fd_sc_ls__conb_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_22_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_870 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
Xoutput52 INVX4/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_ls__clkbuf_4
Xoutput63 XNOR2X1/Y vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_ls__clkbuf_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_2
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XTAP_166 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
.ends

