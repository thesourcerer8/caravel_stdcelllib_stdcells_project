magic
tech sky130A
magscale 1 2
timestamp 1623610208
<< locali >>
rect 29407 52742 29441 52856
rect 16255 51410 16289 51524
rect 11167 50784 11551 50818
rect 11167 50744 11201 50784
rect 34399 50152 34433 50340
rect 22207 41420 22241 41460
rect 22207 41386 22399 41420
rect 21089 34874 21343 34908
rect 21089 34800 21343 34834
rect 8897 33024 9151 33058
rect 7999 19442 8033 19778
rect 21823 12264 21857 12452
rect 23167 10192 23201 10454
rect 12415 9452 12449 9862
rect 13375 7528 13409 7716
rect 17023 6788 17057 7124
rect 8863 6270 8897 6458
rect 27391 4864 27425 4978
rect 20191 3606 20225 3794
rect 19903 3014 19937 3128
rect 19903 2980 20129 3014
rect 20095 2866 20129 2980
rect 21727 2866 21761 2980
rect 22399 2980 22687 3014
rect 22399 2940 22433 2980
rect 41119 2940 41153 3054
rect 44095 2940 44129 3054
<< viali >>
rect 13951 57000 13985 57034
rect 16159 57000 16193 57034
rect 17983 57000 18017 57034
rect 19327 57000 19361 57034
rect 32575 57000 32609 57034
rect 57055 57000 57089 57034
rect 1567 56926 1601 56960
rect 2335 56926 2369 56960
rect 3199 56926 3233 56960
rect 4927 56926 4961 56960
rect 7039 56926 7073 56960
rect 8095 56926 8129 56960
rect 9727 56926 9761 56960
rect 11263 56926 11297 56960
rect 12799 56926 12833 56960
rect 15103 56926 15137 56960
rect 21055 56926 21089 56960
rect 23167 56926 23201 56960
rect 23935 56926 23969 56960
rect 25951 56926 25985 56960
rect 27007 56926 27041 56960
rect 28639 56926 28673 56960
rect 30079 56926 30113 56960
rect 31711 56926 31745 56960
rect 34303 56926 34337 56960
rect 34879 56926 34913 56960
rect 36607 56926 36641 56960
rect 38047 56926 38081 56960
rect 41983 56926 42017 56960
rect 43231 56926 43265 56960
rect 44671 56926 44705 56960
rect 47551 56926 47585 56960
rect 49087 56926 49121 56960
rect 51103 56926 51137 56960
rect 53887 56926 53921 56960
rect 55423 56926 55457 56960
rect 5599 56852 5633 56886
rect 5887 56852 5921 56886
rect 14047 56852 14081 56886
rect 20863 56852 20897 56886
rect 21439 56852 21473 56886
rect 21727 56852 21761 56886
rect 32671 56852 32705 56886
rect 34111 56852 34145 56886
rect 40063 56852 40097 56886
rect 40831 56852 40865 56886
rect 43039 56852 43073 56886
rect 46303 56852 46337 56886
rect 48895 56852 48929 56886
rect 50911 56852 50945 56886
rect 53119 56852 53153 56886
rect 1855 56778 1889 56812
rect 11455 56778 11489 56812
rect 2623 56704 2657 56738
rect 5215 56704 5249 56738
rect 5791 56704 5825 56738
rect 7327 56704 7361 56738
rect 10015 56704 10049 56738
rect 13087 56704 13121 56738
rect 13663 56704 13697 56738
rect 16063 56704 16097 56738
rect 17887 56704 17921 56738
rect 19231 56704 19265 56738
rect 21631 56704 21665 56738
rect 24223 56704 24257 56738
rect 27295 56704 27329 56738
rect 28927 56704 28961 56738
rect 36895 56704 36929 56738
rect 39775 56704 39809 56738
rect 40735 56704 40769 56738
rect 46015 56704 46049 56738
rect 52831 56704 52865 56738
rect 55711 56704 55745 56738
rect 56959 56704 56993 56738
rect 1663 56482 1697 56516
rect 2911 56482 2945 56516
rect 4447 56482 4481 56516
rect 5503 56482 5537 56516
rect 6271 56482 6305 56516
rect 7135 56482 7169 56516
rect 8479 56482 8513 56516
rect 10303 56482 10337 56516
rect 11071 56482 11105 56516
rect 11839 56482 11873 56516
rect 12607 56482 12641 56516
rect 13471 56482 13505 56516
rect 15007 56482 15041 56516
rect 15775 56482 15809 56516
rect 17119 56482 17153 56516
rect 18655 56482 18689 56516
rect 20287 56482 20321 56516
rect 21343 56482 21377 56516
rect 22207 56482 22241 56516
rect 22879 56482 22913 56516
rect 24319 56482 24353 56516
rect 26047 56482 26081 56516
rect 26815 56482 26849 56516
rect 27679 56482 27713 56516
rect 28543 56482 28577 56516
rect 29695 56482 29729 56516
rect 30847 56482 30881 56516
rect 31615 56482 31649 56516
rect 32383 56482 32417 56516
rect 33151 56482 33185 56516
rect 33919 56482 33953 56516
rect 34783 56482 34817 56516
rect 36127 56482 36161 56516
rect 36991 56482 37025 56516
rect 37663 56482 37697 56516
rect 38815 56482 38849 56516
rect 40159 56482 40193 56516
rect 41983 56482 42017 56516
rect 43519 56482 43553 56516
rect 44287 56482 44321 56516
rect 45055 56482 45089 56516
rect 46687 56482 46721 56516
rect 48223 56482 48257 56516
rect 48991 56482 49025 56516
rect 49759 56482 49793 56516
rect 50623 56482 50657 56516
rect 52927 56482 52961 56516
rect 53791 56482 53825 56516
rect 54463 56482 54497 56516
rect 55327 56482 55361 56516
rect 55999 56482 56033 56516
rect 33247 56334 33281 56368
rect 42751 56334 42785 56368
rect 54943 56334 54977 56368
rect 55231 56334 55265 56368
rect 56095 56334 56129 56368
rect 26911 56260 26945 56294
rect 31711 56260 31745 56294
rect 49855 56260 49889 56294
rect 53023 56260 53057 56294
rect 54271 56260 54305 56294
rect 54559 56260 54593 56294
rect 57823 56260 57857 56294
rect 1759 56186 1793 56220
rect 3007 56186 3041 56220
rect 4255 56186 4289 56220
rect 4543 56186 4577 56220
rect 5599 56186 5633 56220
rect 6367 56186 6401 56220
rect 7231 56186 7265 56220
rect 8575 56186 8609 56220
rect 10111 56186 10145 56220
rect 10399 56186 10433 56220
rect 11167 56186 11201 56220
rect 11647 56186 11681 56220
rect 11935 56186 11969 56220
rect 12319 56186 12353 56220
rect 12703 56186 12737 56220
rect 13567 56186 13601 56220
rect 15103 56186 15137 56220
rect 15871 56186 15905 56220
rect 16831 56186 16865 56220
rect 17215 56186 17249 56220
rect 18751 56186 18785 56220
rect 20383 56186 20417 56220
rect 21439 56186 21473 56220
rect 21919 56186 21953 56220
rect 22111 56186 22145 56220
rect 22975 56186 23009 56220
rect 24415 56186 24449 56220
rect 26143 56186 26177 56220
rect 27775 56186 27809 56220
rect 28255 56186 28289 56220
rect 28447 56186 28481 56220
rect 29407 56186 29441 56220
rect 29599 56186 29633 56220
rect 30943 56186 30977 56220
rect 32479 56186 32513 56220
rect 33727 56186 33761 56220
rect 34015 56186 34049 56220
rect 34399 56186 34433 56220
rect 34687 56186 34721 56220
rect 34975 56186 35009 56220
rect 36223 56186 36257 56220
rect 36607 56186 36641 56220
rect 36895 56186 36929 56220
rect 37471 56186 37505 56220
rect 37759 56186 37793 56220
rect 38527 56186 38561 56220
rect 38719 56186 38753 56220
rect 40255 56186 40289 56220
rect 41599 56186 41633 56220
rect 41887 56186 41921 56220
rect 42655 56186 42689 56220
rect 43231 56186 43265 56220
rect 43423 56186 43457 56220
rect 43903 56186 43937 56220
rect 44191 56186 44225 56220
rect 44767 56186 44801 56220
rect 45151 56186 45185 56220
rect 46783 56186 46817 56220
rect 47839 56186 47873 56220
rect 48127 56186 48161 56220
rect 48415 56186 48449 56220
rect 48607 56186 48641 56220
rect 48895 56186 48929 56220
rect 50239 56186 50273 56220
rect 50527 56186 50561 56220
rect 51679 56186 51713 56220
rect 51967 56186 52001 56220
rect 52063 56186 52097 56220
rect 53407 56186 53441 56220
rect 53695 56186 53729 56220
rect 1663 55668 1697 55702
rect 4447 55668 4481 55702
rect 7615 55668 7649 55702
rect 9247 55668 9281 55702
rect 14047 55668 14081 55702
rect 20287 55668 20321 55702
rect 23551 55668 23585 55702
rect 24991 55668 25025 55702
rect 42463 55668 42497 55702
rect 45631 55668 45665 55702
rect 47167 55668 47201 55702
rect 51871 55668 51905 55702
rect 56575 55668 56609 55702
rect 57727 55668 57761 55702
rect 1759 55520 1793 55554
rect 4543 55520 4577 55554
rect 7423 55520 7457 55554
rect 7711 55520 7745 55554
rect 9343 55520 9377 55554
rect 12127 55520 12161 55554
rect 12415 55520 12449 55554
rect 13951 55520 13985 55554
rect 20383 55520 20417 55554
rect 23455 55520 23489 55554
rect 24799 55520 24833 55554
rect 25087 55520 25121 55554
rect 42559 55520 42593 55554
rect 45343 55520 45377 55554
rect 45535 55520 45569 55554
rect 47071 55520 47105 55554
rect 47359 55520 47393 55554
rect 51967 55520 52001 55554
rect 55807 55520 55841 55554
rect 56671 55520 56705 55554
rect 57631 55520 57665 55554
rect 57919 55520 57953 55554
rect 2047 55372 2081 55406
rect 13759 55372 13793 55406
rect 23167 55372 23201 55406
rect 46879 55372 46913 55406
rect 55615 55372 55649 55406
rect 57343 55372 57377 55406
rect 39199 55150 39233 55184
rect 57823 55150 57857 55184
rect 39295 54854 39329 54888
rect 57919 54854 57953 54888
rect 55615 54780 55649 54814
rect 55807 54780 55841 54814
rect 35839 54706 35873 54740
rect 36031 54706 36065 54740
rect 39775 54706 39809 54740
rect 39871 54706 39905 54740
rect 53887 54706 53921 54740
rect 54079 54706 54113 54740
rect 42655 54484 42689 54518
rect 57823 54336 57857 54370
rect 36511 54188 36545 54222
rect 57919 54188 57953 54222
rect 33919 54040 33953 54074
rect 36319 54040 36353 54074
rect 57919 53818 57953 53852
rect 57631 53522 57665 53556
rect 57823 53522 57857 53556
rect 22303 53374 22337 53408
rect 22591 53374 22625 53408
rect 44959 53374 44993 53408
rect 45247 53374 45281 53408
rect 29407 52856 29441 52890
rect 29695 52856 29729 52890
rect 56191 52856 56225 52890
rect 56287 52856 56321 52890
rect 29407 52708 29441 52742
rect 29503 52708 29537 52742
rect 19999 52116 20033 52150
rect 20191 52116 20225 52150
rect 17695 52042 17729 52076
rect 17983 52042 18017 52076
rect 32383 52042 32417 52076
rect 32671 52042 32705 52076
rect 13471 51598 13505 51632
rect 4543 51524 4577 51558
rect 15871 51524 15905 51558
rect 16159 51524 16193 51558
rect 16255 51524 16289 51558
rect 23263 51524 23297 51558
rect 23455 51524 23489 51558
rect 16255 51376 16289 51410
rect 20767 51154 20801 51188
rect 11551 50784 11585 50818
rect 10687 50710 10721 50744
rect 11167 50710 11201 50744
rect 27199 50710 27233 50744
rect 27487 50710 27521 50744
rect 47551 50414 47585 50448
rect 29983 50340 30017 50374
rect 34399 50340 34433 50374
rect 26335 50192 26369 50226
rect 26623 50192 26657 50226
rect 54463 50192 54497 50226
rect 23359 50118 23393 50152
rect 29311 50118 29345 50152
rect 34399 50118 34433 50152
rect 6943 50044 6977 50078
rect 47359 50044 47393 50078
rect 54367 50044 54401 50078
rect 26719 49526 26753 49560
rect 12223 49378 12257 49412
rect 12415 49378 12449 49412
rect 23071 49378 23105 49412
rect 23167 49378 23201 49412
rect 31903 49378 31937 49412
rect 32095 49378 32129 49412
rect 23167 49156 23201 49190
rect 55807 49156 55841 49190
rect 54367 48934 54401 48968
rect 54655 48934 54689 48968
rect 6943 48860 6977 48894
rect 6847 48712 6881 48746
rect 12703 48712 12737 48746
rect 31999 47528 32033 47562
rect 32191 47528 32225 47562
rect 51679 46714 51713 46748
rect 51871 46714 51905 46748
rect 50911 46270 50945 46304
rect 12895 46196 12929 46230
rect 13951 46196 13985 46230
rect 23455 46196 23489 46230
rect 26047 46196 26081 46230
rect 26335 46196 26369 46230
rect 12607 46122 12641 46156
rect 13759 46122 13793 46156
rect 23167 46122 23201 46156
rect 35647 46048 35681 46082
rect 50047 46048 50081 46082
rect 49087 45678 49121 45712
rect 27967 45382 28001 45416
rect 28255 45382 28289 45416
rect 38911 45382 38945 45416
rect 39103 45382 39137 45416
rect 26335 44864 26369 44898
rect 26623 44864 26657 44898
rect 27103 44050 27137 44084
rect 27391 44050 27425 44084
rect 32479 44050 32513 44084
rect 32767 44050 32801 44084
rect 33151 44050 33185 44084
rect 33343 44050 33377 44084
rect 34783 44050 34817 44084
rect 34879 44050 34913 44084
rect 45631 44050 45665 44084
rect 55039 44050 55073 44084
rect 55327 44050 55361 44084
rect 28255 43532 28289 43566
rect 28351 43532 28385 43566
rect 45919 43532 45953 43566
rect 46207 43532 46241 43566
rect 50527 43014 50561 43048
rect 14815 42718 14849 42752
rect 15103 42718 15137 42752
rect 34687 42718 34721 42752
rect 34879 42718 34913 42752
rect 52543 42718 52577 42752
rect 52735 42718 52769 42752
rect 30175 42200 30209 42234
rect 54943 42200 54977 42234
rect 55135 42200 55169 42234
rect 28063 42126 28097 42160
rect 30079 42052 30113 42086
rect 22207 41460 22241 41494
rect 22399 41386 22433 41420
rect 42271 41386 42305 41420
rect 42463 41386 42497 41420
rect 57151 41386 57185 41420
rect 57247 41386 57281 41420
rect 45727 40942 45761 40976
rect 23359 40868 23393 40902
rect 30175 40868 30209 40902
rect 23071 40794 23105 40828
rect 49567 40350 49601 40384
rect 16735 40276 16769 40310
rect 52063 40276 52097 40310
rect 12127 39536 12161 39570
rect 12415 39536 12449 39570
rect 5887 38722 5921 38756
rect 21247 38722 21281 38756
rect 21343 38722 21377 38756
rect 26911 38722 26945 38756
rect 27199 38722 27233 38756
rect 46399 38722 46433 38756
rect 15967 38352 16001 38386
rect 52063 38278 52097 38312
rect 30271 38204 30305 38238
rect 30559 38204 30593 38238
rect 57727 38204 57761 38238
rect 57823 38204 57857 38238
rect 41503 37464 41537 37498
rect 43039 37464 43073 37498
rect 16351 37390 16385 37424
rect 16447 37390 16481 37424
rect 41791 37390 41825 37424
rect 43231 37390 43265 37424
rect 53887 37390 53921 37424
rect 54079 37390 54113 37424
rect 2719 36206 2753 36240
rect 1663 36058 1697 36092
rect 1951 36058 1985 36092
rect 22399 36058 22433 36092
rect 22591 36058 22625 36092
rect 38527 36058 38561 36092
rect 54751 36058 54785 36092
rect 54847 36058 54881 36092
rect 2335 35540 2369 35574
rect 2623 35540 2657 35574
rect 20479 35540 20513 35574
rect 21343 35540 21377 35574
rect 21631 35540 21665 35574
rect 45055 35540 45089 35574
rect 49183 35540 49217 35574
rect 51391 35540 51425 35574
rect 9439 35466 9473 35500
rect 44863 35392 44897 35426
rect 48991 35392 49025 35426
rect 51199 35392 51233 35426
rect 4543 35022 4577 35056
rect 21055 34874 21089 34908
rect 21343 34874 21377 34908
rect 21055 34800 21089 34834
rect 21343 34800 21377 34834
rect 17791 34726 17825 34760
rect 20863 34726 20897 34760
rect 50047 34726 50081 34760
rect 50239 34726 50273 34760
rect 21343 34208 21377 34242
rect 36703 34208 36737 34242
rect 52543 33468 52577 33502
rect 52735 33468 52769 33502
rect 45631 33394 45665 33428
rect 57343 33172 57377 33206
rect 8863 33024 8897 33058
rect 9151 33024 9185 33058
rect 13087 32062 13121 32096
rect 26527 31692 26561 31726
rect 57343 31692 57377 31726
rect 23071 30878 23105 30912
rect 20863 30360 20897 30394
rect 46783 30286 46817 30320
rect 27967 29398 28001 29432
rect 28255 29398 28289 29432
rect 9343 28880 9377 28914
rect 28927 28880 28961 28914
rect 9055 28806 9089 28840
rect 46399 28510 46433 28544
rect 46591 28362 46625 28396
rect 38047 28214 38081 28248
rect 38143 28214 38177 28248
rect 6271 28066 6305 28100
rect 57343 28066 57377 28100
rect 58015 28066 58049 28100
rect 37759 27030 37793 27064
rect 38047 27030 38081 27064
rect 12511 26734 12545 26768
rect 40159 26216 40193 26250
rect 47743 26216 47777 26250
rect 54655 26216 54689 26250
rect 13567 25698 13601 25732
rect 13855 25698 13889 25732
rect 4447 25476 4481 25510
rect 4735 25476 4769 25510
rect 5407 25402 5441 25436
rect 39775 25402 39809 25436
rect 15679 24958 15713 24992
rect 26623 24884 26657 24918
rect 26911 24884 26945 24918
rect 36703 24884 36737 24918
rect 8575 23552 8609 23586
rect 13663 23552 13697 23586
rect 41887 23552 41921 23586
rect 45535 23552 45569 23586
rect 20479 23034 20513 23068
rect 20767 23034 20801 23068
rect 8671 22738 8705 22772
rect 24031 22738 24065 22772
rect 36319 22738 36353 22772
rect 57343 22738 57377 22772
rect 15103 22220 15137 22254
rect 20575 22220 20609 22254
rect 34975 22220 35009 22254
rect 5119 21406 5153 21440
rect 15103 21406 15137 21440
rect 37087 20888 37121 20922
rect 47647 20888 47681 20922
rect 47743 20888 47777 20922
rect 7999 19778 8033 19812
rect 1759 19556 1793 19590
rect 8479 19556 8513 19590
rect 13951 19556 13985 19590
rect 28255 19556 28289 19590
rect 38911 19556 38945 19590
rect 7999 19408 8033 19442
rect 5503 18816 5537 18850
rect 34015 18224 34049 18258
rect 27103 17558 27137 17592
rect 27295 17558 27329 17592
rect 54079 17484 54113 17518
rect 23167 17410 23201 17444
rect 46783 17410 46817 17444
rect 2815 16966 2849 17000
rect 3103 16966 3137 17000
rect 10495 16892 10529 16926
rect 35551 16892 35585 16926
rect 46111 16892 46145 16926
rect 54655 16892 54689 16926
rect 53503 16226 53537 16260
rect 53311 16078 53345 16112
rect 9823 15856 9857 15890
rect 32287 14746 32321 14780
rect 48991 14524 49025 14558
rect 49183 14524 49217 14558
rect 46591 14450 46625 14484
rect 44671 14080 44705 14114
rect 44863 14080 44897 14114
rect 12415 13488 12449 13522
rect 5311 13414 5345 13448
rect 57727 13192 57761 13226
rect 57823 13192 57857 13226
rect 9727 12970 9761 13004
rect 29887 12970 29921 13004
rect 49375 12970 49409 13004
rect 57343 12526 57377 12560
rect 21823 12452 21857 12486
rect 57631 12378 57665 12412
rect 20767 12230 20801 12264
rect 21055 12230 21089 12264
rect 21823 12230 21857 12264
rect 29791 12230 29825 12264
rect 57727 12230 57761 12264
rect 9631 12082 9665 12116
rect 9919 12082 9953 12116
rect 39871 11860 39905 11894
rect 40063 11860 40097 11894
rect 56191 11860 56225 11894
rect 22687 11786 22721 11820
rect 29311 11786 29345 11820
rect 56479 11712 56513 11746
rect 56575 11712 56609 11746
rect 39487 11638 39521 11672
rect 56959 11638 56993 11672
rect 57247 11638 57281 11672
rect 14623 11564 14657 11598
rect 57327 11564 57361 11598
rect 31135 11194 31169 11228
rect 31423 11194 31457 11228
rect 57343 11046 57377 11080
rect 56095 10972 56129 11006
rect 55999 10898 56033 10932
rect 57247 10898 57281 10932
rect 6943 10750 6977 10784
rect 15679 10750 15713 10784
rect 42655 10750 42689 10784
rect 54367 10750 54401 10784
rect 56287 10528 56321 10562
rect 23167 10454 23201 10488
rect 12607 10232 12641 10266
rect 54847 10380 54881 10414
rect 55039 10380 55073 10414
rect 55327 10380 55361 10414
rect 55903 10380 55937 10414
rect 56575 10380 56609 10414
rect 57439 10380 57473 10414
rect 38815 10232 38849 10266
rect 23167 10158 23201 10192
rect 55135 10084 55169 10118
rect 55807 10084 55841 10118
rect 56671 10084 56705 10118
rect 57343 10084 57377 10118
rect 12415 9862 12449 9896
rect 4447 9492 4481 9526
rect 26239 9714 26273 9748
rect 26431 9714 26465 9748
rect 54847 9714 54881 9748
rect 55135 9714 55169 9748
rect 55711 9714 55745 9748
rect 55903 9714 55937 9748
rect 56191 9714 56225 9748
rect 57631 9640 57665 9674
rect 54367 9566 54401 9600
rect 54463 9566 54497 9600
rect 55231 9566 55265 9600
rect 55999 9566 56033 9600
rect 53407 9492 53441 9526
rect 53599 9492 53633 9526
rect 12415 9418 12449 9452
rect 45631 9418 45665 9452
rect 46783 9418 46817 9452
rect 54271 9196 54305 9230
rect 38815 9048 38849 9082
rect 53119 9048 53153 9082
rect 53311 9048 53345 9082
rect 53407 9048 53441 9082
rect 54655 9048 54689 9082
rect 55039 8974 55073 9008
rect 55327 8974 55361 9008
rect 56575 8974 56609 9008
rect 57247 8974 57281 9008
rect 1759 8900 1793 8934
rect 3487 8900 3521 8934
rect 52735 8900 52769 8934
rect 54559 8900 54593 8934
rect 10975 8752 11009 8786
rect 11263 8752 11297 8786
rect 55423 8752 55457 8786
rect 2143 8530 2177 8564
rect 39103 8530 39137 8564
rect 42271 8530 42305 8564
rect 44095 8530 44129 8564
rect 48223 8530 48257 8564
rect 52255 8530 52289 8564
rect 52927 8530 52961 8564
rect 2527 8382 2561 8416
rect 4255 8382 4289 8416
rect 4543 8382 4577 8416
rect 10783 8382 10817 8416
rect 11263 8382 11297 8416
rect 11551 8382 11585 8416
rect 12319 8382 12353 8416
rect 16255 8382 16289 8416
rect 16735 8382 16769 8416
rect 17023 8382 17057 8416
rect 39295 8382 39329 8416
rect 42559 8382 42593 8416
rect 44383 8382 44417 8416
rect 47551 8382 47585 8416
rect 47839 8382 47873 8416
rect 48511 8382 48545 8416
rect 49375 8382 49409 8416
rect 50143 8382 50177 8416
rect 52447 8382 52481 8416
rect 53215 8382 53249 8416
rect 54079 8382 54113 8416
rect 2911 8308 2945 8342
rect 3295 8308 3329 8342
rect 55231 8308 55265 8342
rect 55999 8308 56033 8342
rect 57151 8308 57185 8342
rect 1663 8234 1697 8268
rect 1759 8234 1793 8268
rect 2431 8234 2465 8268
rect 3199 8234 3233 8268
rect 4447 8234 4481 8268
rect 10687 8234 10721 8268
rect 11455 8234 11489 8268
rect 12223 8234 12257 8268
rect 12991 8234 13025 8268
rect 13087 8234 13121 8268
rect 16159 8234 16193 8268
rect 16927 8234 16961 8268
rect 39391 8234 39425 8268
rect 42655 8234 42689 8268
rect 44479 8234 44513 8268
rect 47743 8234 47777 8268
rect 48607 8234 48641 8268
rect 49279 8234 49313 8268
rect 50047 8234 50081 8268
rect 52543 8234 52577 8268
rect 53311 8234 53345 8268
rect 53983 8234 54017 8268
rect 2047 8160 2081 8194
rect 40159 8160 40193 8194
rect 7519 8086 7553 8120
rect 13855 8086 13889 8120
rect 43423 8086 43457 8120
rect 12127 7864 12161 7898
rect 12799 7864 12833 7898
rect 13567 7864 13601 7898
rect 15103 7864 15137 7898
rect 17695 7864 17729 7898
rect 17983 7864 18017 7898
rect 27967 7864 28001 7898
rect 30847 7864 30881 7898
rect 32383 7864 32417 7898
rect 35839 7864 35873 7898
rect 39967 7864 40001 7898
rect 43711 7864 43745 7898
rect 44479 7864 44513 7898
rect 45247 7864 45281 7898
rect 46879 7864 46913 7898
rect 48991 7864 49025 7898
rect 49759 7864 49793 7898
rect 4543 7790 4577 7824
rect 3967 7716 4001 7750
rect 4735 7716 4769 7750
rect 4831 7716 4865 7750
rect 10111 7716 10145 7750
rect 10591 7716 10625 7750
rect 10879 7716 10913 7750
rect 12319 7716 12353 7750
rect 12415 7716 12449 7750
rect 13375 7716 13409 7750
rect 13951 7716 13985 7750
rect 15391 7716 15425 7750
rect 15967 7716 16001 7750
rect 16255 7716 16289 7750
rect 20671 7716 20705 7750
rect 20959 7716 20993 7750
rect 23935 7716 23969 7750
rect 24415 7716 24449 7750
rect 24703 7716 24737 7750
rect 25471 7716 25505 7750
rect 26239 7716 26273 7750
rect 27007 7716 27041 7750
rect 28351 7716 28385 7750
rect 29119 7716 29153 7750
rect 29407 7716 29441 7750
rect 29887 7716 29921 7750
rect 30175 7716 30209 7750
rect 31135 7716 31169 7750
rect 34303 7716 34337 7750
rect 34591 7716 34625 7750
rect 35359 7716 35393 7750
rect 36031 7716 36065 7750
rect 36607 7716 36641 7750
rect 36799 7716 36833 7750
rect 38815 7716 38849 7750
rect 39295 7716 39329 7750
rect 39487 7716 39521 7750
rect 40255 7716 40289 7750
rect 41119 7716 41153 7750
rect 41887 7716 41921 7750
rect 42367 7716 42401 7750
rect 42655 7716 42689 7750
rect 44095 7716 44129 7750
rect 44767 7716 44801 7750
rect 45535 7716 45569 7750
rect 46399 7716 46433 7750
rect 47071 7716 47105 7750
rect 47935 7716 47969 7750
rect 49279 7716 49313 7750
rect 50047 7716 50081 7750
rect 51103 7716 51137 7750
rect 52639 7716 52673 7750
rect 53407 7716 53441 7750
rect 1567 7642 1601 7676
rect 2239 7642 2273 7676
rect 2527 7642 2561 7676
rect 5599 7642 5633 7676
rect 3007 7568 3041 7602
rect 3295 7568 3329 7602
rect 4063 7568 4097 7602
rect 9343 7568 9377 7602
rect 13087 7568 13121 7602
rect 53119 7642 53153 7676
rect 53311 7642 53345 7676
rect 55135 7642 55169 7676
rect 55807 7642 55841 7676
rect 56575 7642 56609 7676
rect 57343 7642 57377 7676
rect 18655 7568 18689 7602
rect 21727 7568 21761 7602
rect 33823 7568 33857 7602
rect 51871 7568 51905 7602
rect 13375 7494 13409 7528
rect 2431 7420 2465 7454
rect 3199 7420 3233 7454
rect 5503 7420 5537 7454
rect 9247 7420 9281 7454
rect 10015 7420 10049 7454
rect 10783 7420 10817 7454
rect 13183 7420 13217 7454
rect 13855 7420 13889 7454
rect 15487 7420 15521 7454
rect 16159 7420 16193 7454
rect 20863 7420 20897 7454
rect 23839 7420 23873 7454
rect 24607 7420 24641 7454
rect 25375 7420 25409 7454
rect 26143 7420 26177 7454
rect 26911 7420 26945 7454
rect 28255 7420 28289 7454
rect 29311 7420 29345 7454
rect 30079 7420 30113 7454
rect 31231 7420 31265 7454
rect 33727 7420 33761 7454
rect 34495 7420 34529 7454
rect 35263 7420 35297 7454
rect 36127 7420 36161 7454
rect 36895 7420 36929 7454
rect 38719 7420 38753 7454
rect 39583 7420 39617 7454
rect 40351 7420 40385 7454
rect 41023 7420 41057 7454
rect 41791 7420 41825 7454
rect 42559 7420 42593 7454
rect 43999 7420 44033 7454
rect 44863 7420 44897 7454
rect 45631 7420 45665 7454
rect 46303 7420 46337 7454
rect 47167 7420 47201 7454
rect 47839 7420 47873 7454
rect 49375 7420 49409 7454
rect 50143 7420 50177 7454
rect 51007 7420 51041 7454
rect 51775 7420 51809 7454
rect 52543 7420 52577 7454
rect 17215 7198 17249 7232
rect 31615 7198 31649 7232
rect 33919 7198 33953 7232
rect 42175 7198 42209 7232
rect 6463 7124 6497 7158
rect 7999 7124 8033 7158
rect 17023 7124 17057 7158
rect 22303 7124 22337 7158
rect 28351 7124 28385 7158
rect 38911 7124 38945 7158
rect 6847 7050 6881 7084
rect 7327 7050 7361 7084
rect 7615 7050 7649 7084
rect 8383 7050 8417 7084
rect 9823 7050 9857 7084
rect 15103 7050 15137 7084
rect 15871 7050 15905 7084
rect 1663 6976 1697 7010
rect 2527 6976 2561 7010
rect 4255 6976 4289 7010
rect 4543 6976 4577 7010
rect 11263 6976 11297 7010
rect 12703 6976 12737 7010
rect 4447 6902 4481 6936
rect 5215 6902 5249 6936
rect 5311 6902 5345 6936
rect 5983 6902 6017 6936
rect 6079 6902 6113 6936
rect 6751 6902 6785 6936
rect 7519 6902 7553 6936
rect 8287 6902 8321 6936
rect 9727 6902 9761 6936
rect 10495 6902 10529 6936
rect 10591 6902 10625 6936
rect 13567 6902 13601 6936
rect 13663 6902 13697 6936
rect 15007 6902 15041 6936
rect 15775 6902 15809 6936
rect 5791 6828 5825 6862
rect 10303 6828 10337 6862
rect 17791 7050 17825 7084
rect 18079 7050 18113 7084
rect 18847 7050 18881 7084
rect 20095 7050 20129 7084
rect 20383 7050 20417 7084
rect 21151 7050 21185 7084
rect 21919 7050 21953 7084
rect 22591 7050 22625 7084
rect 23455 7050 23489 7084
rect 24223 7050 24257 7084
rect 25663 7050 25697 7084
rect 26431 7050 26465 7084
rect 27199 7050 27233 7084
rect 27967 7050 28001 7084
rect 28639 7050 28673 7084
rect 29503 7050 29537 7084
rect 31711 7050 31745 7084
rect 32479 7050 32513 7084
rect 33247 7050 33281 7084
rect 34015 7050 34049 7084
rect 36703 7050 36737 7084
rect 36895 7050 36929 7084
rect 37183 7050 37217 7084
rect 37471 7050 37505 7084
rect 37663 7050 37697 7084
rect 38527 7050 38561 7084
rect 39295 7050 39329 7084
rect 40063 7050 40097 7084
rect 41503 7050 41537 7084
rect 42271 7050 42305 7084
rect 42751 7050 42785 7084
rect 42943 7050 42977 7084
rect 43727 7050 43761 7084
rect 44287 7050 44321 7084
rect 44575 7050 44609 7084
rect 46783 7050 46817 7084
rect 47167 7050 47201 7084
rect 47455 7050 47489 7084
rect 48319 7050 48353 7084
rect 49087 7050 49121 7084
rect 50335 7050 50369 7084
rect 52063 7050 52097 7084
rect 52447 7050 52481 7084
rect 52735 7050 52769 7084
rect 23375 6976 23409 7010
rect 30943 6976 30977 7010
rect 36223 6976 36257 7010
rect 54079 6976 54113 7010
rect 54751 6976 54785 7010
rect 55519 6976 55553 7010
rect 57823 6976 57857 7010
rect 17311 6902 17345 6936
rect 17983 6902 18017 6936
rect 18751 6902 18785 6936
rect 20287 6902 20321 6936
rect 21055 6902 21089 6936
rect 21823 6902 21857 6936
rect 22687 6902 22721 6936
rect 24127 6902 24161 6936
rect 25567 6902 25601 6936
rect 26335 6902 26369 6936
rect 27103 6902 27137 6936
rect 27871 6902 27905 6936
rect 28735 6902 28769 6936
rect 29407 6902 29441 6936
rect 30847 6902 30881 6936
rect 32383 6902 32417 6936
rect 33151 6902 33185 6936
rect 34687 6902 34721 6936
rect 34783 6902 34817 6936
rect 36127 6902 36161 6936
rect 36991 6902 37025 6936
rect 37759 6902 37793 6936
rect 38431 6902 38465 6936
rect 39199 6902 39233 6936
rect 39967 6902 40001 6936
rect 41407 6902 41441 6936
rect 43039 6902 43073 6936
rect 43807 6902 43841 6936
rect 44479 6902 44513 6936
rect 45247 6902 45281 6936
rect 45343 6902 45377 6936
rect 46687 6902 46721 6936
rect 47551 6902 47585 6936
rect 48223 6902 48257 6936
rect 48991 6902 49025 6936
rect 50239 6902 50273 6936
rect 51967 6902 52001 6936
rect 52831 6902 52865 6936
rect 17023 6754 17057 6788
rect 18943 6532 18977 6566
rect 33151 6532 33185 6566
rect 36895 6532 36929 6566
rect 50623 6532 50657 6566
rect 8383 6458 8417 6492
rect 8863 6458 8897 6492
rect 9151 6458 9185 6492
rect 7135 6384 7169 6418
rect 1567 6310 1601 6344
rect 2335 6310 2369 6344
rect 3199 6310 3233 6344
rect 3967 6310 4001 6344
rect 4735 6310 4769 6344
rect 5695 6310 5729 6344
rect 9343 6384 9377 6418
rect 9439 6384 9473 6418
rect 13951 6384 13985 6418
rect 14719 6384 14753 6418
rect 15199 6384 15233 6418
rect 15487 6384 15521 6418
rect 18463 6384 18497 6418
rect 19231 6384 19265 6418
rect 19711 6384 19745 6418
rect 19999 6384 20033 6418
rect 20479 6384 20513 6418
rect 20767 6384 20801 6418
rect 21247 6384 21281 6418
rect 21535 6384 21569 6418
rect 22687 6384 22721 6418
rect 22975 6384 23009 6418
rect 23743 6384 23777 6418
rect 24223 6384 24257 6418
rect 24511 6384 24545 6418
rect 27967 6384 28001 6418
rect 28159 6384 28193 6418
rect 28735 6384 28769 6418
rect 29023 6384 29057 6418
rect 30655 6384 30689 6418
rect 32191 6384 32225 6418
rect 50815 6384 50849 6418
rect 51679 6384 51713 6418
rect 52351 6384 52385 6418
rect 10111 6310 10145 6344
rect 10879 6310 10913 6344
rect 12223 6310 12257 6344
rect 12991 6310 13025 6344
rect 16351 6310 16385 6344
rect 25663 6310 25697 6344
rect 26815 6310 26849 6344
rect 29695 6310 29729 6344
rect 31231 6310 31265 6344
rect 34223 6310 34257 6344
rect 36319 6310 36353 6344
rect 37263 6310 37297 6344
rect 38911 6310 38945 6344
rect 40351 6310 40385 6344
rect 41503 6310 41537 6344
rect 42271 6310 42305 6344
rect 43903 6310 43937 6344
rect 44767 6310 44801 6344
rect 45535 6310 45569 6344
rect 46975 6310 47009 6344
rect 47743 6310 47777 6344
rect 49183 6310 49217 6344
rect 49951 6310 49985 6344
rect 53311 6310 53345 6344
rect 54463 6310 54497 6344
rect 55231 6310 55265 6344
rect 55999 6310 56033 6344
rect 57055 6310 57089 6344
rect 57823 6310 57857 6344
rect 7903 6236 7937 6270
rect 8671 6236 8705 6270
rect 8863 6236 8897 6270
rect 17695 6236 17729 6270
rect 33535 6236 33569 6270
rect 34303 6236 34337 6270
rect 35071 6236 35105 6270
rect 37183 6236 37217 6270
rect 52447 6236 52481 6270
rect 5599 6088 5633 6122
rect 7039 6088 7073 6122
rect 7807 6088 7841 6122
rect 8575 6088 8609 6122
rect 13855 6088 13889 6122
rect 14623 6088 14657 6122
rect 15391 6088 15425 6122
rect 17599 6088 17633 6122
rect 18367 6088 18401 6122
rect 19135 6088 19169 6122
rect 19903 6088 19937 6122
rect 20671 6088 20705 6122
rect 21439 6088 21473 6122
rect 22879 6088 22913 6122
rect 23647 6088 23681 6122
rect 24415 6088 24449 6122
rect 28255 6088 28289 6122
rect 28927 6088 28961 6122
rect 30559 6088 30593 6122
rect 32095 6088 32129 6122
rect 33439 6088 33473 6122
rect 34975 6088 35009 6122
rect 50911 6088 50945 6122
rect 51583 6088 51617 6122
rect 55039 5866 55073 5900
rect 55231 5866 55265 5900
rect 6079 5718 6113 5752
rect 1567 5644 1601 5678
rect 2911 5644 2945 5678
rect 4447 5644 4481 5678
rect 5119 5644 5153 5678
rect 7231 5644 7265 5678
rect 7999 5644 8033 5678
rect 9631 5644 9665 5678
rect 10399 5644 10433 5678
rect 11167 5644 11201 5678
rect 12607 5644 12641 5678
rect 13375 5644 13409 5678
rect 15007 5644 15041 5678
rect 15871 5644 15905 5678
rect 16543 5644 16577 5678
rect 17983 5644 18017 5678
rect 18751 5644 18785 5678
rect 20191 5644 20225 5678
rect 20959 5644 20993 5678
rect 21727 5644 21761 5678
rect 22495 5644 22529 5678
rect 23263 5644 23297 5678
rect 24031 5644 24065 5678
rect 25471 5644 25505 5678
rect 26239 5644 26273 5678
rect 27007 5644 27041 5678
rect 27775 5644 27809 5678
rect 28543 5644 28577 5678
rect 29311 5644 29345 5678
rect 30751 5644 30785 5678
rect 31519 5644 31553 5678
rect 32287 5644 32321 5678
rect 33151 5644 33185 5678
rect 33823 5644 33857 5678
rect 34687 5644 34721 5678
rect 36127 5644 36161 5678
rect 36799 5644 36833 5678
rect 37567 5644 37601 5678
rect 38335 5644 38369 5678
rect 39103 5644 39137 5678
rect 39871 5644 39905 5678
rect 41311 5644 41345 5678
rect 43903 5644 43937 5678
rect 44671 5644 44705 5678
rect 46591 5644 46625 5678
rect 47359 5644 47393 5678
rect 48127 5644 48161 5678
rect 48991 5644 49025 5678
rect 49663 5644 49697 5678
rect 50527 5644 50561 5678
rect 52159 5644 52193 5678
rect 52927 5644 52961 5678
rect 53695 5644 53729 5678
rect 54463 5644 54497 5678
rect 55999 5644 56033 5678
rect 57439 5644 57473 5678
rect 5983 5570 6017 5604
rect 11839 5422 11873 5456
rect 12127 5422 12161 5456
rect 17215 5422 17249 5456
rect 17503 5422 17537 5456
rect 1567 4978 1601 5012
rect 2335 4978 2369 5012
rect 3103 4978 3137 5012
rect 4159 4978 4193 5012
rect 5407 4978 5441 5012
rect 6943 4978 6977 5012
rect 7711 4978 7745 5012
rect 8479 4978 8513 5012
rect 9247 4978 9281 5012
rect 10111 4978 10145 5012
rect 10783 4978 10817 5012
rect 12223 4978 12257 5012
rect 12991 4978 13025 5012
rect 13951 4978 13985 5012
rect 14719 4978 14753 5012
rect 15487 4978 15521 5012
rect 16351 4978 16385 5012
rect 17503 4978 17537 5012
rect 18271 4978 18305 5012
rect 19039 4978 19073 5012
rect 19807 4978 19841 5012
rect 20575 4978 20609 5012
rect 21343 4978 21377 5012
rect 22783 4978 22817 5012
rect 23551 4978 23585 5012
rect 24319 4978 24353 5012
rect 25087 4978 25121 5012
rect 25855 4978 25889 5012
rect 26623 4978 26657 5012
rect 27391 4978 27425 5012
rect 28063 4978 28097 5012
rect 28927 4978 28961 5012
rect 29599 4978 29633 5012
rect 30367 4978 30401 5012
rect 31135 4978 31169 5012
rect 31903 4978 31937 5012
rect 33343 4978 33377 5012
rect 34111 4978 34145 5012
rect 34879 4978 34913 5012
rect 35647 4978 35681 5012
rect 36415 4978 36449 5012
rect 37183 4978 37217 5012
rect 38623 4978 38657 5012
rect 39391 4978 39425 5012
rect 40159 4978 40193 5012
rect 40927 4978 40961 5012
rect 41695 4978 41729 5012
rect 42463 4978 42497 5012
rect 43903 4978 43937 5012
rect 44671 4978 44705 5012
rect 45439 4978 45473 5012
rect 46207 4978 46241 5012
rect 46975 4978 47009 5012
rect 47839 4978 47873 5012
rect 49375 4978 49409 5012
rect 50431 4978 50465 5012
rect 51103 4978 51137 5012
rect 51871 4978 51905 5012
rect 52639 4978 52673 5012
rect 54463 4978 54497 5012
rect 55615 4978 55649 5012
rect 56383 4978 56417 5012
rect 57055 4978 57089 5012
rect 58015 4904 58049 4938
rect 27391 4830 27425 4864
rect 15775 4534 15809 4568
rect 19135 4534 19169 4568
rect 38143 4534 38177 4568
rect 38335 4534 38369 4568
rect 16543 4460 16577 4494
rect 17311 4460 17345 4494
rect 1567 4312 1601 4346
rect 2335 4312 2369 4346
rect 3103 4312 3137 4346
rect 4351 4312 4385 4346
rect 5119 4312 5153 4346
rect 5887 4312 5921 4346
rect 6655 4312 6689 4346
rect 7423 4312 7457 4346
rect 8191 4312 8225 4346
rect 9631 4312 9665 4346
rect 10399 4312 10433 4346
rect 11167 4312 11201 4346
rect 11935 4312 11969 4346
rect 12703 4312 12737 4346
rect 13567 4312 13601 4346
rect 15487 4312 15521 4346
rect 16255 4312 16289 4346
rect 17023 4312 17057 4346
rect 17791 4312 17825 4346
rect 18847 4312 18881 4346
rect 20191 4312 20225 4346
rect 21055 4312 21089 4346
rect 21823 4312 21857 4346
rect 23263 4312 23297 4346
rect 24031 4312 24065 4346
rect 25471 4312 25505 4346
rect 26239 4312 26273 4346
rect 27007 4312 27041 4346
rect 28351 4312 28385 4346
rect 29119 4312 29153 4346
rect 30943 4312 30977 4346
rect 31711 4312 31745 4346
rect 32767 4312 32801 4346
rect 33919 4312 33953 4346
rect 34687 4312 34721 4346
rect 36031 4312 36065 4346
rect 36799 4312 36833 4346
rect 37567 4312 37601 4346
rect 39007 4312 39041 4346
rect 39775 4312 39809 4346
rect 41983 4312 42017 4346
rect 42751 4312 42785 4346
rect 43519 4312 43553 4346
rect 44959 4312 44993 4346
rect 46783 4312 46817 4346
rect 47551 4312 47585 4346
rect 48319 4312 48353 4346
rect 49087 4312 49121 4346
rect 49855 4312 49889 4346
rect 50623 4312 50657 4346
rect 51871 4312 51905 4346
rect 52639 4312 52673 4346
rect 53407 4312 53441 4346
rect 54175 4312 54209 4346
rect 55615 4312 55649 4346
rect 57151 4312 57185 4346
rect 22783 4238 22817 4272
rect 55135 4238 55169 4272
rect 41503 4164 41537 4198
rect 20191 3794 20225 3828
rect 13567 3720 13601 3754
rect 15295 3720 15329 3754
rect 17695 3720 17729 3754
rect 18559 3720 18593 3754
rect 1567 3646 1601 3680
rect 2335 3646 2369 3680
rect 3103 3646 3137 3680
rect 3871 3646 3905 3680
rect 4639 3646 4673 3680
rect 5599 3646 5633 3680
rect 6943 3646 6977 3680
rect 7711 3646 7745 3680
rect 8479 3646 8513 3680
rect 9247 3646 9281 3680
rect 10015 3646 10049 3680
rect 10783 3646 10817 3680
rect 12703 3646 12737 3680
rect 13759 3646 13793 3680
rect 14623 3646 14657 3680
rect 15871 3646 15905 3680
rect 17887 3646 17921 3680
rect 18751 3646 18785 3680
rect 19231 3646 19265 3680
rect 20671 3646 20705 3680
rect 21151 3646 21185 3680
rect 22783 3646 22817 3680
rect 23551 3646 23585 3680
rect 24319 3646 24353 3680
rect 25087 3646 25121 3680
rect 25855 3646 25889 3680
rect 26623 3646 26657 3680
rect 28063 3646 28097 3680
rect 28831 3646 28865 3680
rect 29599 3646 29633 3680
rect 30367 3646 30401 3680
rect 31135 3646 31169 3680
rect 31903 3646 31937 3680
rect 33343 3646 33377 3680
rect 34111 3646 34145 3680
rect 34879 3646 34913 3680
rect 35647 3646 35681 3680
rect 36415 3646 36449 3680
rect 37183 3646 37217 3680
rect 38623 3646 38657 3680
rect 39391 3646 39425 3680
rect 40159 3646 40193 3680
rect 40927 3646 40961 3680
rect 41695 3646 41729 3680
rect 42463 3646 42497 3680
rect 43903 3646 43937 3680
rect 44671 3646 44705 3680
rect 45439 3646 45473 3680
rect 46207 3646 46241 3680
rect 46975 3646 47009 3680
rect 47743 3646 47777 3680
rect 49183 3646 49217 3680
rect 50527 3646 50561 3680
rect 51199 3646 51233 3680
rect 51967 3646 52001 3680
rect 52735 3646 52769 3680
rect 54463 3646 54497 3680
rect 55231 3646 55265 3680
rect 55999 3646 56033 3680
rect 56767 3646 56801 3680
rect 57535 3646 57569 3680
rect 14431 3572 14465 3606
rect 20191 3572 20225 3606
rect 20479 3572 20513 3606
rect 15199 3424 15233 3458
rect 21631 3202 21665 3236
rect 19903 3128 19937 3162
rect 51391 3128 51425 3162
rect 15295 3054 15329 3088
rect 18847 3054 18881 3088
rect 41119 3054 41153 3088
rect 1567 2980 1601 3014
rect 2335 2980 2369 3014
rect 3103 2980 3137 3014
rect 4927 2980 4961 3014
rect 5695 2980 5729 3014
rect 7039 2980 7073 3014
rect 7807 2980 7841 3014
rect 9727 2980 9761 3014
rect 10495 2980 10529 3014
rect 13375 2980 13409 3014
rect 13951 2980 13985 3014
rect 15487 2980 15521 3014
rect 16639 2980 16673 3014
rect 18175 2980 18209 3014
rect 19039 2980 19073 3014
rect 20863 2980 20897 3014
rect 21343 2980 21377 3014
rect 21727 2980 21761 3014
rect 13183 2906 13217 2940
rect 17983 2906 18017 2940
rect 20671 2906 20705 2940
rect 20095 2832 20129 2866
rect 22687 2980 22721 3014
rect 23167 2980 23201 3014
rect 23935 2980 23969 3014
rect 25855 2980 25889 3014
rect 26623 2980 26657 3014
rect 28543 2980 28577 3014
rect 29311 2980 29345 3014
rect 31231 2980 31265 3014
rect 31999 2980 32033 3014
rect 33919 2980 33953 3014
rect 34687 2980 34721 3014
rect 36607 2980 36641 3014
rect 37375 2980 37409 3014
rect 39295 2980 39329 3014
rect 40063 2980 40097 3014
rect 22399 2906 22433 2940
rect 44095 3054 44129 3088
rect 46399 3054 46433 3088
rect 51583 3054 51617 3088
rect 41983 2980 42017 3014
rect 42751 2980 42785 3014
rect 41119 2906 41153 2940
rect 44671 2980 44705 3014
rect 45439 2980 45473 3014
rect 47359 2980 47393 3014
rect 48127 2980 48161 3014
rect 50047 2980 50081 3014
rect 50815 2980 50849 3014
rect 52735 2980 52769 3014
rect 53503 2980 53537 3014
rect 55423 2980 55457 3014
rect 56191 2980 56225 3014
rect 44095 2906 44129 2940
rect 21727 2832 21761 2866
rect 57151 2832 57185 2866
rect 24895 2758 24929 2792
rect 54463 2758 54497 2792
<< metal1 >>
rect 1152 57302 58848 57324
rect 1152 57250 4294 57302
rect 4346 57250 4358 57302
rect 4410 57250 4422 57302
rect 4474 57250 4486 57302
rect 4538 57250 35014 57302
rect 35066 57250 35078 57302
rect 35130 57250 35142 57302
rect 35194 57250 35206 57302
rect 35258 57250 58848 57302
rect 1152 57228 58848 57250
rect 16432 57105 16438 57117
rect 13954 57077 16438 57105
rect 13954 57040 13982 57077
rect 16432 57065 16438 57077
rect 16490 57065 16496 57117
rect 13939 57034 13997 57040
rect 13939 57000 13951 57034
rect 13985 57000 13997 57034
rect 13939 56994 13997 57000
rect 15952 56991 15958 57043
rect 16010 57031 16016 57043
rect 16147 57034 16205 57040
rect 16147 57031 16159 57034
rect 16010 57003 16159 57031
rect 16010 56991 16016 57003
rect 16147 57000 16159 57003
rect 16193 57000 16205 57034
rect 16147 56994 16205 57000
rect 17488 56991 17494 57043
rect 17546 57031 17552 57043
rect 17971 57034 18029 57040
rect 17971 57031 17983 57034
rect 17546 57003 17983 57031
rect 17546 56991 17552 57003
rect 17971 57000 17983 57003
rect 18017 57000 18029 57034
rect 17971 56994 18029 57000
rect 19120 56991 19126 57043
rect 19178 57031 19184 57043
rect 19315 57034 19373 57040
rect 19315 57031 19327 57034
rect 19178 57003 19327 57031
rect 19178 56991 19184 57003
rect 19315 57000 19327 57003
rect 19361 57000 19373 57034
rect 19315 56994 19373 57000
rect 29104 56991 29110 57043
rect 29162 57031 29168 57043
rect 32563 57034 32621 57040
rect 32563 57031 32575 57034
rect 29162 57003 32575 57031
rect 29162 56991 29168 57003
rect 32563 57000 32575 57003
rect 32609 57000 32621 57034
rect 57040 57031 57046 57043
rect 57001 57003 57046 57031
rect 32563 56994 32621 57000
rect 57040 56991 57046 57003
rect 57098 56991 57104 57043
rect 208 56917 214 56969
rect 266 56957 272 56969
rect 1555 56960 1613 56966
rect 1555 56957 1567 56960
rect 266 56929 1567 56957
rect 266 56917 272 56929
rect 1555 56926 1567 56929
rect 1601 56926 1613 56960
rect 1555 56920 1613 56926
rect 1744 56917 1750 56969
rect 1802 56957 1808 56969
rect 2323 56960 2381 56966
rect 2323 56957 2335 56960
rect 1802 56929 2335 56957
rect 1802 56917 1808 56929
rect 2323 56926 2335 56929
rect 2369 56926 2381 56960
rect 2323 56920 2381 56926
rect 3187 56960 3245 56966
rect 3187 56926 3199 56960
rect 3233 56957 3245 56960
rect 3280 56957 3286 56969
rect 3233 56929 3286 56957
rect 3233 56926 3245 56929
rect 3187 56920 3245 56926
rect 3280 56917 3286 56929
rect 3338 56917 3344 56969
rect 4912 56957 4918 56969
rect 4873 56929 4918 56957
rect 4912 56917 4918 56929
rect 4970 56917 4976 56969
rect 6448 56917 6454 56969
rect 6506 56957 6512 56969
rect 7027 56960 7085 56966
rect 7027 56957 7039 56960
rect 6506 56929 7039 56957
rect 6506 56917 6512 56929
rect 7027 56926 7039 56929
rect 7073 56926 7085 56960
rect 8080 56957 8086 56969
rect 8041 56929 8086 56957
rect 7027 56920 7085 56926
rect 8080 56917 8086 56929
rect 8138 56917 8144 56969
rect 9616 56917 9622 56969
rect 9674 56957 9680 56969
rect 9715 56960 9773 56966
rect 9715 56957 9727 56960
rect 9674 56929 9727 56957
rect 9674 56917 9680 56929
rect 9715 56926 9727 56929
rect 9761 56926 9773 56960
rect 11248 56957 11254 56969
rect 11209 56929 11254 56957
rect 9715 56920 9773 56926
rect 11248 56917 11254 56929
rect 11306 56917 11312 56969
rect 12784 56957 12790 56969
rect 12745 56929 12790 56957
rect 12784 56917 12790 56929
rect 12842 56917 12848 56969
rect 14416 56917 14422 56969
rect 14474 56957 14480 56969
rect 15091 56960 15149 56966
rect 15091 56957 15103 56960
rect 14474 56929 15103 56957
rect 14474 56917 14480 56929
rect 15091 56926 15103 56929
rect 15137 56926 15149 56960
rect 15091 56920 15149 56926
rect 20656 56917 20662 56969
rect 20714 56957 20720 56969
rect 21043 56960 21101 56966
rect 21043 56957 21055 56960
rect 20714 56929 21055 56957
rect 20714 56917 20720 56929
rect 21043 56926 21055 56929
rect 21089 56926 21101 56960
rect 21043 56920 21101 56926
rect 22288 56917 22294 56969
rect 22346 56957 22352 56969
rect 23155 56960 23213 56966
rect 23155 56957 23167 56960
rect 22346 56929 23167 56957
rect 22346 56917 22352 56929
rect 23155 56926 23167 56929
rect 23201 56926 23213 56960
rect 23155 56920 23213 56926
rect 23824 56917 23830 56969
rect 23882 56957 23888 56969
rect 23923 56960 23981 56966
rect 23923 56957 23935 56960
rect 23882 56929 23935 56957
rect 23882 56917 23888 56929
rect 23923 56926 23935 56929
rect 23969 56926 23981 56960
rect 23923 56920 23981 56926
rect 25456 56917 25462 56969
rect 25514 56957 25520 56969
rect 25939 56960 25997 56966
rect 25939 56957 25951 56960
rect 25514 56929 25951 56957
rect 25514 56917 25520 56929
rect 25939 56926 25951 56929
rect 25985 56926 25997 56960
rect 26992 56957 26998 56969
rect 26953 56929 26998 56957
rect 25939 56920 25997 56926
rect 26992 56917 26998 56929
rect 27050 56917 27056 56969
rect 28624 56957 28630 56969
rect 28585 56929 28630 56957
rect 28624 56917 28630 56929
rect 28682 56917 28688 56969
rect 30067 56960 30125 56966
rect 30067 56926 30079 56960
rect 30113 56957 30125 56960
rect 30160 56957 30166 56969
rect 30113 56929 30166 56957
rect 30113 56926 30125 56929
rect 30067 56920 30125 56926
rect 30160 56917 30166 56929
rect 30218 56917 30224 56969
rect 31696 56957 31702 56969
rect 31657 56929 31702 56957
rect 31696 56917 31702 56929
rect 31754 56917 31760 56969
rect 33328 56917 33334 56969
rect 33386 56957 33392 56969
rect 34291 56960 34349 56966
rect 34291 56957 34303 56960
rect 33386 56929 34303 56957
rect 33386 56917 33392 56929
rect 34291 56926 34303 56929
rect 34337 56926 34349 56960
rect 34864 56957 34870 56969
rect 34825 56929 34870 56957
rect 34291 56920 34349 56926
rect 34864 56917 34870 56929
rect 34922 56917 34928 56969
rect 36496 56917 36502 56969
rect 36554 56957 36560 56969
rect 36595 56960 36653 56966
rect 36595 56957 36607 56960
rect 36554 56929 36607 56957
rect 36554 56917 36560 56929
rect 36595 56926 36607 56929
rect 36641 56926 36653 56960
rect 38032 56957 38038 56969
rect 37993 56929 38038 56957
rect 36595 56920 36653 56926
rect 38032 56917 38038 56929
rect 38090 56917 38096 56969
rect 41200 56917 41206 56969
rect 41258 56957 41264 56969
rect 41971 56960 42029 56966
rect 41971 56957 41983 56960
rect 41258 56929 41983 56957
rect 41258 56917 41264 56929
rect 41971 56926 41983 56929
rect 42017 56926 42029 56960
rect 41971 56920 42029 56926
rect 42832 56917 42838 56969
rect 42890 56957 42896 56969
rect 43219 56960 43277 56966
rect 43219 56957 43231 56960
rect 42890 56929 43231 56957
rect 42890 56917 42896 56929
rect 43219 56926 43231 56929
rect 43265 56926 43277 56960
rect 43219 56920 43277 56926
rect 44368 56917 44374 56969
rect 44426 56957 44432 56969
rect 44659 56960 44717 56966
rect 44659 56957 44671 56960
rect 44426 56929 44671 56957
rect 44426 56917 44432 56929
rect 44659 56926 44671 56929
rect 44705 56926 44717 56960
rect 44659 56920 44717 56926
rect 47536 56917 47542 56969
rect 47594 56957 47600 56969
rect 49072 56957 49078 56969
rect 47594 56929 47639 56957
rect 49033 56929 49078 56957
rect 47594 56917 47600 56929
rect 49072 56917 49078 56929
rect 49130 56917 49136 56969
rect 50704 56917 50710 56969
rect 50762 56957 50768 56969
rect 51091 56960 51149 56966
rect 51091 56957 51103 56960
rect 50762 56929 51103 56957
rect 50762 56917 50768 56929
rect 51091 56926 51103 56929
rect 51137 56926 51149 56960
rect 53872 56957 53878 56969
rect 53833 56929 53878 56957
rect 51091 56920 51149 56926
rect 53872 56917 53878 56929
rect 53930 56917 53936 56969
rect 55408 56957 55414 56969
rect 55369 56929 55414 56957
rect 55408 56917 55414 56929
rect 55466 56917 55472 56969
rect 5587 56886 5645 56892
rect 5587 56852 5599 56886
rect 5633 56883 5645 56886
rect 5875 56886 5933 56892
rect 5875 56883 5887 56886
rect 5633 56855 5887 56883
rect 5633 56852 5645 56855
rect 5587 56846 5645 56852
rect 5875 56852 5887 56855
rect 5921 56883 5933 56886
rect 7888 56883 7894 56895
rect 5921 56855 7894 56883
rect 5921 56852 5933 56855
rect 5875 56846 5933 56852
rect 7888 56843 7894 56855
rect 7946 56843 7952 56895
rect 14035 56886 14093 56892
rect 14035 56883 14047 56886
rect 13666 56855 14047 56883
rect 1843 56812 1901 56818
rect 1843 56778 1855 56812
rect 1889 56809 1901 56812
rect 6064 56809 6070 56821
rect 1889 56781 6070 56809
rect 1889 56778 1901 56781
rect 1843 56772 1901 56778
rect 6064 56769 6070 56781
rect 6122 56769 6128 56821
rect 9040 56769 9046 56821
rect 9098 56809 9104 56821
rect 11443 56812 11501 56818
rect 11443 56809 11455 56812
rect 9098 56781 11455 56809
rect 9098 56769 9104 56781
rect 11443 56778 11455 56781
rect 11489 56778 11501 56812
rect 11443 56772 11501 56778
rect 13666 56747 13694 56855
rect 14035 56852 14047 56855
rect 14081 56852 14093 56886
rect 20848 56883 20854 56895
rect 20809 56855 20854 56883
rect 14035 56846 14093 56852
rect 20848 56843 20854 56855
rect 20906 56843 20912 56895
rect 21427 56886 21485 56892
rect 21427 56852 21439 56886
rect 21473 56883 21485 56886
rect 21616 56883 21622 56895
rect 21473 56855 21622 56883
rect 21473 56852 21485 56855
rect 21427 56846 21485 56852
rect 21616 56843 21622 56855
rect 21674 56883 21680 56895
rect 21715 56886 21773 56892
rect 21715 56883 21727 56886
rect 21674 56855 21727 56883
rect 21674 56843 21680 56855
rect 21715 56852 21727 56855
rect 21761 56852 21773 56886
rect 21715 56846 21773 56852
rect 32560 56843 32566 56895
rect 32618 56883 32624 56895
rect 32659 56886 32717 56892
rect 32659 56883 32671 56886
rect 32618 56855 32671 56883
rect 32618 56843 32624 56855
rect 32659 56852 32671 56855
rect 32705 56852 32717 56886
rect 34096 56883 34102 56895
rect 34057 56855 34102 56883
rect 32659 56846 32717 56852
rect 34096 56843 34102 56855
rect 34154 56843 34160 56895
rect 39664 56843 39670 56895
rect 39722 56883 39728 56895
rect 40051 56886 40109 56892
rect 40051 56883 40063 56886
rect 39722 56855 40063 56883
rect 39722 56843 39728 56855
rect 40051 56852 40063 56855
rect 40097 56852 40109 56886
rect 40816 56883 40822 56895
rect 40777 56855 40822 56883
rect 40051 56846 40109 56852
rect 40816 56843 40822 56855
rect 40874 56843 40880 56895
rect 43024 56883 43030 56895
rect 42985 56855 43030 56883
rect 43024 56843 43030 56855
rect 43082 56843 43088 56895
rect 45904 56843 45910 56895
rect 45962 56883 45968 56895
rect 46291 56886 46349 56892
rect 46291 56883 46303 56886
rect 45962 56855 46303 56883
rect 45962 56843 45968 56855
rect 46291 56852 46303 56855
rect 46337 56852 46349 56886
rect 48880 56883 48886 56895
rect 48841 56855 48886 56883
rect 46291 56846 46349 56852
rect 48880 56843 48886 56855
rect 48938 56843 48944 56895
rect 50896 56883 50902 56895
rect 50857 56855 50902 56883
rect 50896 56843 50902 56855
rect 50954 56843 50960 56895
rect 52240 56843 52246 56895
rect 52298 56883 52304 56895
rect 53107 56886 53165 56892
rect 53107 56883 53119 56886
rect 52298 56855 53119 56883
rect 52298 56843 52304 56855
rect 53107 56852 53119 56855
rect 53153 56852 53165 56886
rect 53107 56846 53165 56852
rect 32464 56769 32470 56821
rect 32522 56809 32528 56821
rect 39856 56809 39862 56821
rect 32522 56781 39862 56809
rect 32522 56769 32528 56781
rect 39856 56769 39862 56781
rect 39914 56769 39920 56821
rect 42832 56769 42838 56821
rect 42890 56809 42896 56821
rect 54832 56809 54838 56821
rect 42890 56781 54838 56809
rect 42890 56769 42896 56781
rect 54832 56769 54838 56781
rect 54890 56769 54896 56821
rect 2611 56738 2669 56744
rect 2611 56704 2623 56738
rect 2657 56735 2669 56738
rect 4816 56735 4822 56747
rect 2657 56707 4822 56735
rect 2657 56704 2669 56707
rect 2611 56698 2669 56704
rect 4816 56695 4822 56707
rect 4874 56695 4880 56747
rect 5200 56735 5206 56747
rect 5161 56707 5206 56735
rect 5200 56695 5206 56707
rect 5258 56695 5264 56747
rect 5776 56735 5782 56747
rect 5737 56707 5782 56735
rect 5776 56695 5782 56707
rect 5834 56695 5840 56747
rect 7312 56735 7318 56747
rect 7273 56707 7318 56735
rect 7312 56695 7318 56707
rect 7370 56695 7376 56747
rect 10000 56735 10006 56747
rect 9961 56707 10006 56735
rect 10000 56695 10006 56707
rect 10058 56695 10064 56747
rect 13072 56735 13078 56747
rect 13033 56707 13078 56735
rect 13072 56695 13078 56707
rect 13130 56695 13136 56747
rect 13648 56735 13654 56747
rect 13609 56707 13654 56735
rect 13648 56695 13654 56707
rect 13706 56695 13712 56747
rect 16048 56735 16054 56747
rect 16009 56707 16054 56735
rect 16048 56695 16054 56707
rect 16106 56695 16112 56747
rect 17872 56735 17878 56747
rect 17833 56707 17878 56735
rect 17872 56695 17878 56707
rect 17930 56695 17936 56747
rect 19216 56735 19222 56747
rect 19177 56707 19222 56735
rect 19216 56695 19222 56707
rect 19274 56695 19280 56747
rect 21619 56738 21677 56744
rect 21619 56704 21631 56738
rect 21665 56735 21677 56738
rect 21808 56735 21814 56747
rect 21665 56707 21814 56735
rect 21665 56704 21677 56707
rect 21619 56698 21677 56704
rect 21808 56695 21814 56707
rect 21866 56695 21872 56747
rect 22000 56695 22006 56747
rect 22058 56735 22064 56747
rect 24211 56738 24269 56744
rect 24211 56735 24223 56738
rect 22058 56707 24223 56735
rect 22058 56695 22064 56707
rect 24211 56704 24223 56707
rect 24257 56704 24269 56738
rect 27280 56735 27286 56747
rect 27241 56707 27286 56735
rect 24211 56698 24269 56704
rect 27280 56695 27286 56707
rect 27338 56695 27344 56747
rect 28915 56738 28973 56744
rect 28915 56704 28927 56738
rect 28961 56735 28973 56738
rect 36112 56735 36118 56747
rect 28961 56707 36118 56735
rect 28961 56704 28973 56707
rect 28915 56698 28973 56704
rect 36112 56695 36118 56707
rect 36170 56695 36176 56747
rect 36880 56735 36886 56747
rect 36841 56707 36886 56735
rect 36880 56695 36886 56707
rect 36938 56695 36944 56747
rect 39664 56695 39670 56747
rect 39722 56735 39728 56747
rect 39763 56738 39821 56744
rect 39763 56735 39775 56738
rect 39722 56707 39775 56735
rect 39722 56695 39728 56707
rect 39763 56704 39775 56707
rect 39809 56704 39821 56738
rect 39763 56698 39821 56704
rect 40336 56695 40342 56747
rect 40394 56735 40400 56747
rect 40723 56738 40781 56744
rect 40723 56735 40735 56738
rect 40394 56707 40735 56735
rect 40394 56695 40400 56707
rect 40723 56704 40735 56707
rect 40769 56704 40781 56738
rect 40723 56698 40781 56704
rect 46003 56738 46061 56744
rect 46003 56704 46015 56738
rect 46049 56735 46061 56738
rect 46096 56735 46102 56747
rect 46049 56707 46102 56735
rect 46049 56704 46061 56707
rect 46003 56698 46061 56704
rect 46096 56695 46102 56707
rect 46154 56695 46160 56747
rect 52816 56735 52822 56747
rect 52777 56707 52822 56735
rect 52816 56695 52822 56707
rect 52874 56695 52880 56747
rect 55696 56735 55702 56747
rect 55657 56707 55702 56735
rect 55696 56695 55702 56707
rect 55754 56695 55760 56747
rect 56944 56735 56950 56747
rect 56905 56707 56950 56735
rect 56944 56695 56950 56707
rect 57002 56695 57008 56747
rect 1152 56636 58848 56658
rect 1152 56584 19654 56636
rect 19706 56584 19718 56636
rect 19770 56584 19782 56636
rect 19834 56584 19846 56636
rect 19898 56584 50374 56636
rect 50426 56584 50438 56636
rect 50490 56584 50502 56636
rect 50554 56584 50566 56636
rect 50618 56584 58848 56636
rect 1152 56562 58848 56584
rect 688 56473 694 56525
rect 746 56513 752 56525
rect 1651 56516 1709 56522
rect 1651 56513 1663 56516
rect 746 56485 1663 56513
rect 746 56473 752 56485
rect 1651 56482 1663 56485
rect 1697 56482 1709 56516
rect 1651 56476 1709 56482
rect 2800 56473 2806 56525
rect 2858 56513 2864 56525
rect 2899 56516 2957 56522
rect 2899 56513 2911 56516
rect 2858 56485 2911 56513
rect 2858 56473 2864 56485
rect 2899 56482 2911 56485
rect 2945 56482 2957 56516
rect 2899 56476 2957 56482
rect 3856 56473 3862 56525
rect 3914 56513 3920 56525
rect 4435 56516 4493 56522
rect 4435 56513 4447 56516
rect 3914 56485 4447 56513
rect 3914 56473 3920 56485
rect 4435 56482 4447 56485
rect 4481 56482 4493 56516
rect 4435 56476 4493 56482
rect 5392 56473 5398 56525
rect 5450 56513 5456 56525
rect 5491 56516 5549 56522
rect 5491 56513 5503 56516
rect 5450 56485 5503 56513
rect 5450 56473 5456 56485
rect 5491 56482 5503 56485
rect 5537 56482 5549 56516
rect 5491 56476 5549 56482
rect 5968 56473 5974 56525
rect 6026 56513 6032 56525
rect 6259 56516 6317 56522
rect 6259 56513 6271 56516
rect 6026 56485 6271 56513
rect 6026 56473 6032 56485
rect 6259 56482 6271 56485
rect 6305 56482 6317 56516
rect 6259 56476 6317 56482
rect 7024 56473 7030 56525
rect 7082 56513 7088 56525
rect 7123 56516 7181 56522
rect 7123 56513 7135 56516
rect 7082 56485 7135 56513
rect 7082 56473 7088 56485
rect 7123 56482 7135 56485
rect 7169 56482 7181 56516
rect 7123 56476 7181 56482
rect 8467 56516 8525 56522
rect 8467 56482 8479 56516
rect 8513 56513 8525 56516
rect 8560 56513 8566 56525
rect 8513 56485 8566 56513
rect 8513 56482 8525 56485
rect 8467 56476 8525 56482
rect 8560 56473 8566 56485
rect 8618 56473 8624 56525
rect 10192 56473 10198 56525
rect 10250 56513 10256 56525
rect 10291 56516 10349 56522
rect 10291 56513 10303 56516
rect 10250 56485 10303 56513
rect 10250 56473 10256 56485
rect 10291 56482 10303 56485
rect 10337 56482 10349 56516
rect 10291 56476 10349 56482
rect 10672 56473 10678 56525
rect 10730 56513 10736 56525
rect 11059 56516 11117 56522
rect 11059 56513 11071 56516
rect 10730 56485 11071 56513
rect 10730 56473 10736 56485
rect 11059 56482 11071 56485
rect 11105 56482 11117 56516
rect 11059 56476 11117 56482
rect 11728 56473 11734 56525
rect 11786 56513 11792 56525
rect 11827 56516 11885 56522
rect 11827 56513 11839 56516
rect 11786 56485 11839 56513
rect 11786 56473 11792 56485
rect 11827 56482 11839 56485
rect 11873 56482 11885 56516
rect 11827 56476 11885 56482
rect 12304 56473 12310 56525
rect 12362 56513 12368 56525
rect 12595 56516 12653 56522
rect 12595 56513 12607 56516
rect 12362 56485 12607 56513
rect 12362 56473 12368 56485
rect 12595 56482 12607 56485
rect 12641 56482 12653 56516
rect 12595 56476 12653 56482
rect 13360 56473 13366 56525
rect 13418 56513 13424 56525
rect 13459 56516 13517 56522
rect 13459 56513 13471 56516
rect 13418 56485 13471 56513
rect 13418 56473 13424 56485
rect 13459 56482 13471 56485
rect 13505 56482 13517 56516
rect 13459 56476 13517 56482
rect 14896 56473 14902 56525
rect 14954 56513 14960 56525
rect 14995 56516 15053 56522
rect 14995 56513 15007 56516
rect 14954 56485 15007 56513
rect 14954 56473 14960 56485
rect 14995 56482 15007 56485
rect 15041 56482 15053 56516
rect 14995 56476 15053 56482
rect 15376 56473 15382 56525
rect 15434 56513 15440 56525
rect 15763 56516 15821 56522
rect 15763 56513 15775 56516
rect 15434 56485 15775 56513
rect 15434 56473 15440 56485
rect 15763 56482 15775 56485
rect 15809 56482 15821 56516
rect 15763 56476 15821 56482
rect 17008 56473 17014 56525
rect 17066 56513 17072 56525
rect 17107 56516 17165 56522
rect 17107 56513 17119 56516
rect 17066 56485 17119 56513
rect 17066 56473 17072 56485
rect 17107 56482 17119 56485
rect 17153 56482 17165 56516
rect 17107 56476 17165 56482
rect 18544 56473 18550 56525
rect 18602 56513 18608 56525
rect 18643 56516 18701 56522
rect 18643 56513 18655 56516
rect 18602 56485 18655 56513
rect 18602 56473 18608 56485
rect 18643 56482 18655 56485
rect 18689 56482 18701 56516
rect 18643 56476 18701 56482
rect 19984 56473 19990 56525
rect 20042 56513 20048 56525
rect 20275 56516 20333 56522
rect 20275 56513 20287 56516
rect 20042 56485 20287 56513
rect 20042 56473 20048 56485
rect 20275 56482 20287 56485
rect 20321 56482 20333 56516
rect 20275 56476 20333 56482
rect 21232 56473 21238 56525
rect 21290 56513 21296 56525
rect 21331 56516 21389 56522
rect 21331 56513 21343 56516
rect 21290 56485 21343 56513
rect 21290 56473 21296 56485
rect 21331 56482 21343 56485
rect 21377 56482 21389 56516
rect 21331 56476 21389 56482
rect 21712 56473 21718 56525
rect 21770 56513 21776 56525
rect 22195 56516 22253 56522
rect 22195 56513 22207 56516
rect 21770 56485 22207 56513
rect 21770 56473 21776 56485
rect 22195 56482 22207 56485
rect 22241 56482 22253 56516
rect 22195 56476 22253 56482
rect 22768 56473 22774 56525
rect 22826 56513 22832 56525
rect 22867 56516 22925 56522
rect 22867 56513 22879 56516
rect 22826 56485 22879 56513
rect 22826 56473 22832 56485
rect 22867 56482 22879 56485
rect 22913 56482 22925 56516
rect 22867 56476 22925 56482
rect 24307 56516 24365 56522
rect 24307 56482 24319 56516
rect 24353 56513 24365 56516
rect 24400 56513 24406 56525
rect 24353 56485 24406 56513
rect 24353 56482 24365 56485
rect 24307 56476 24365 56482
rect 24400 56473 24406 56485
rect 24458 56473 24464 56525
rect 25936 56473 25942 56525
rect 25994 56513 26000 56525
rect 26035 56516 26093 56522
rect 26035 56513 26047 56516
rect 25994 56485 26047 56513
rect 25994 56473 26000 56485
rect 26035 56482 26047 56485
rect 26081 56482 26093 56516
rect 26035 56476 26093 56482
rect 26512 56473 26518 56525
rect 26570 56513 26576 56525
rect 26803 56516 26861 56522
rect 26803 56513 26815 56516
rect 26570 56485 26815 56513
rect 26570 56473 26576 56485
rect 26803 56482 26815 56485
rect 26849 56482 26861 56516
rect 26803 56476 26861 56482
rect 27568 56473 27574 56525
rect 27626 56513 27632 56525
rect 27667 56516 27725 56522
rect 27667 56513 27679 56516
rect 27626 56485 27679 56513
rect 27626 56473 27632 56485
rect 27667 56482 27679 56485
rect 27713 56482 27725 56516
rect 27667 56476 27725 56482
rect 28048 56473 28054 56525
rect 28106 56513 28112 56525
rect 28531 56516 28589 56522
rect 28531 56513 28543 56516
rect 28106 56485 28543 56513
rect 28106 56473 28112 56485
rect 28531 56482 28543 56485
rect 28577 56482 28589 56516
rect 29680 56513 29686 56525
rect 29641 56485 29686 56513
rect 28531 56476 28589 56482
rect 29680 56473 29686 56485
rect 29738 56473 29744 56525
rect 30640 56473 30646 56525
rect 30698 56513 30704 56525
rect 30835 56516 30893 56522
rect 30835 56513 30847 56516
rect 30698 56485 30847 56513
rect 30698 56473 30704 56485
rect 30835 56482 30847 56485
rect 30881 56482 30893 56516
rect 30835 56476 30893 56482
rect 31216 56473 31222 56525
rect 31274 56513 31280 56525
rect 31603 56516 31661 56522
rect 31603 56513 31615 56516
rect 31274 56485 31615 56513
rect 31274 56473 31280 56485
rect 31603 56482 31615 56485
rect 31649 56482 31661 56516
rect 31603 56476 31661 56482
rect 32272 56473 32278 56525
rect 32330 56513 32336 56525
rect 32371 56516 32429 56522
rect 32371 56513 32383 56516
rect 32330 56485 32383 56513
rect 32330 56473 32336 56485
rect 32371 56482 32383 56485
rect 32417 56482 32429 56516
rect 32371 56476 32429 56482
rect 32752 56473 32758 56525
rect 32810 56513 32816 56525
rect 33139 56516 33197 56522
rect 33139 56513 33151 56516
rect 32810 56485 33151 56513
rect 32810 56473 32816 56485
rect 33139 56482 33151 56485
rect 33185 56482 33197 56516
rect 33139 56476 33197 56482
rect 33808 56473 33814 56525
rect 33866 56513 33872 56525
rect 33907 56516 33965 56522
rect 33907 56513 33919 56516
rect 33866 56485 33919 56513
rect 33866 56473 33872 56485
rect 33907 56482 33919 56485
rect 33953 56482 33965 56516
rect 33907 56476 33965 56482
rect 34576 56473 34582 56525
rect 34634 56513 34640 56525
rect 34771 56516 34829 56522
rect 34771 56513 34783 56516
rect 34634 56485 34783 56513
rect 34634 56473 34640 56485
rect 34771 56482 34783 56485
rect 34817 56482 34829 56516
rect 34771 56476 34829 56482
rect 35440 56473 35446 56525
rect 35498 56513 35504 56525
rect 36115 56516 36173 56522
rect 36115 56513 36127 56516
rect 35498 56485 36127 56513
rect 35498 56473 35504 56485
rect 36115 56482 36127 56485
rect 36161 56482 36173 56516
rect 36115 56476 36173 56482
rect 36979 56516 37037 56522
rect 36979 56482 36991 56516
rect 37025 56482 37037 56516
rect 36979 56476 37037 56482
rect 27280 56399 27286 56451
rect 27338 56439 27344 56451
rect 32464 56439 32470 56451
rect 27338 56411 32470 56439
rect 27338 56399 27344 56411
rect 32464 56399 32470 56411
rect 32522 56399 32528 56451
rect 36016 56399 36022 56451
rect 36074 56439 36080 56451
rect 36994 56439 37022 56476
rect 37552 56473 37558 56525
rect 37610 56513 37616 56525
rect 37651 56516 37709 56522
rect 37651 56513 37663 56516
rect 37610 56485 37663 56513
rect 37610 56473 37616 56485
rect 37651 56482 37663 56485
rect 37697 56482 37709 56516
rect 37651 56476 37709 56482
rect 38608 56473 38614 56525
rect 38666 56513 38672 56525
rect 38803 56516 38861 56522
rect 38803 56513 38815 56516
rect 38666 56485 38815 56513
rect 38666 56473 38672 56485
rect 38803 56482 38815 56485
rect 38849 56482 38861 56516
rect 40144 56513 40150 56525
rect 40105 56485 40150 56513
rect 38803 56476 38861 56482
rect 40144 56473 40150 56485
rect 40202 56473 40208 56525
rect 41776 56473 41782 56525
rect 41834 56513 41840 56525
rect 41971 56516 42029 56522
rect 41971 56513 41983 56516
rect 41834 56485 41983 56513
rect 41834 56473 41840 56485
rect 41971 56482 41983 56485
rect 42017 56482 42029 56516
rect 41971 56476 42029 56482
rect 43312 56473 43318 56525
rect 43370 56513 43376 56525
rect 43507 56516 43565 56522
rect 43507 56513 43519 56516
rect 43370 56485 43519 56513
rect 43370 56473 43376 56485
rect 43507 56482 43519 56485
rect 43553 56482 43565 56516
rect 43507 56476 43565 56482
rect 43888 56473 43894 56525
rect 43946 56513 43952 56525
rect 44275 56516 44333 56522
rect 44275 56513 44287 56516
rect 43946 56485 44287 56513
rect 43946 56473 43952 56485
rect 44275 56482 44287 56485
rect 44321 56482 44333 56516
rect 44275 56476 44333 56482
rect 44944 56473 44950 56525
rect 45002 56513 45008 56525
rect 45043 56516 45101 56522
rect 45043 56513 45055 56516
rect 45002 56485 45055 56513
rect 45002 56473 45008 56485
rect 45043 56482 45055 56485
rect 45089 56482 45101 56516
rect 45043 56476 45101 56482
rect 46480 56473 46486 56525
rect 46538 56513 46544 56525
rect 46675 56516 46733 56522
rect 46675 56513 46687 56516
rect 46538 56485 46687 56513
rect 46538 56473 46544 56485
rect 46675 56482 46687 56485
rect 46721 56482 46733 56516
rect 46675 56476 46733 56482
rect 48016 56473 48022 56525
rect 48074 56513 48080 56525
rect 48211 56516 48269 56522
rect 48211 56513 48223 56516
rect 48074 56485 48223 56513
rect 48074 56473 48080 56485
rect 48211 56482 48223 56485
rect 48257 56482 48269 56516
rect 48211 56476 48269 56482
rect 48592 56473 48598 56525
rect 48650 56513 48656 56525
rect 48979 56516 49037 56522
rect 48979 56513 48991 56516
rect 48650 56485 48991 56513
rect 48650 56473 48656 56485
rect 48979 56482 48991 56485
rect 49025 56482 49037 56516
rect 48979 56476 49037 56482
rect 49648 56473 49654 56525
rect 49706 56513 49712 56525
rect 49747 56516 49805 56522
rect 49747 56513 49759 56516
rect 49706 56485 49759 56513
rect 49706 56473 49712 56485
rect 49747 56482 49759 56485
rect 49793 56482 49805 56516
rect 49747 56476 49805 56482
rect 50128 56473 50134 56525
rect 50186 56513 50192 56525
rect 50611 56516 50669 56522
rect 50611 56513 50623 56516
rect 50186 56485 50623 56513
rect 50186 56473 50192 56485
rect 50611 56482 50623 56485
rect 50657 56482 50669 56516
rect 52912 56513 52918 56525
rect 52873 56485 52918 56513
rect 50611 56476 50669 56482
rect 52912 56473 52918 56485
rect 52970 56473 52976 56525
rect 53296 56473 53302 56525
rect 53354 56513 53360 56525
rect 53779 56516 53837 56522
rect 53779 56513 53791 56516
rect 53354 56485 53791 56513
rect 53354 56473 53360 56485
rect 53779 56482 53791 56485
rect 53825 56482 53837 56516
rect 53779 56476 53837 56482
rect 54352 56473 54358 56525
rect 54410 56513 54416 56525
rect 54451 56516 54509 56522
rect 54451 56513 54463 56516
rect 54410 56485 54463 56513
rect 54410 56473 54416 56485
rect 54451 56482 54463 56485
rect 54497 56482 54509 56516
rect 54451 56476 54509 56482
rect 54928 56473 54934 56525
rect 54986 56513 54992 56525
rect 55315 56516 55373 56522
rect 55315 56513 55327 56516
rect 54986 56485 55327 56513
rect 54986 56473 54992 56485
rect 55315 56482 55327 56485
rect 55361 56482 55373 56516
rect 55984 56513 55990 56525
rect 55945 56485 55990 56513
rect 55315 56476 55373 56482
rect 55984 56473 55990 56485
rect 56042 56473 56048 56525
rect 38896 56439 38902 56451
rect 36074 56411 37022 56439
rect 37426 56411 38902 56439
rect 36074 56399 36080 56411
rect 33235 56368 33293 56374
rect 33235 56334 33247 56368
rect 33281 56365 33293 56368
rect 37426 56365 37454 56411
rect 38896 56399 38902 56411
rect 38954 56399 38960 56451
rect 46192 56399 46198 56451
rect 46250 56439 46256 56451
rect 46250 56411 56126 56439
rect 46250 56399 46256 56411
rect 33281 56337 37454 56365
rect 42739 56368 42797 56374
rect 33281 56334 33293 56337
rect 33235 56328 33293 56334
rect 42739 56334 42751 56368
rect 42785 56365 42797 56368
rect 48304 56365 48310 56377
rect 42785 56337 48310 56365
rect 42785 56334 42797 56337
rect 42739 56328 42797 56334
rect 48304 56325 48310 56337
rect 48362 56325 48368 56377
rect 54832 56325 54838 56377
rect 54890 56365 54896 56377
rect 56098 56374 56126 56411
rect 54931 56368 54989 56374
rect 54931 56365 54943 56368
rect 54890 56337 54943 56365
rect 54890 56325 54896 56337
rect 54931 56334 54943 56337
rect 54977 56365 54989 56368
rect 55219 56368 55277 56374
rect 55219 56365 55231 56368
rect 54977 56337 55231 56365
rect 54977 56334 54989 56337
rect 54931 56328 54989 56334
rect 55219 56334 55231 56337
rect 55265 56334 55277 56368
rect 55219 56328 55277 56334
rect 56083 56368 56141 56374
rect 56083 56334 56095 56368
rect 56129 56334 56141 56368
rect 56083 56328 56141 56334
rect 22864 56251 22870 56303
rect 22922 56291 22928 56303
rect 26899 56294 26957 56300
rect 26899 56291 26911 56294
rect 22922 56263 26911 56291
rect 22922 56251 22928 56263
rect 26899 56260 26911 56263
rect 26945 56260 26957 56294
rect 26899 56254 26957 56260
rect 31699 56294 31757 56300
rect 31699 56260 31711 56294
rect 31745 56291 31757 56294
rect 41776 56291 41782 56303
rect 31745 56263 41782 56291
rect 31745 56260 31757 56263
rect 31699 56254 31757 56260
rect 41776 56251 41782 56263
rect 41834 56251 41840 56303
rect 46288 56251 46294 56303
rect 46346 56291 46352 56303
rect 49843 56294 49901 56300
rect 49843 56291 49855 56294
rect 46346 56263 49855 56291
rect 46346 56251 46352 56263
rect 49843 56260 49855 56263
rect 49889 56260 49901 56294
rect 49843 56254 49901 56260
rect 50032 56251 50038 56303
rect 50090 56291 50096 56303
rect 53011 56294 53069 56300
rect 53011 56291 53023 56294
rect 50090 56263 53023 56291
rect 50090 56251 50096 56263
rect 53011 56260 53023 56263
rect 53057 56260 53069 56294
rect 53011 56254 53069 56260
rect 54259 56294 54317 56300
rect 54259 56260 54271 56294
rect 54305 56291 54317 56294
rect 54547 56294 54605 56300
rect 54547 56291 54559 56294
rect 54305 56263 54559 56291
rect 54305 56260 54317 56263
rect 54259 56254 54317 56260
rect 54547 56260 54559 56263
rect 54593 56291 54605 56294
rect 57811 56294 57869 56300
rect 54593 56263 57614 56291
rect 54593 56260 54605 56263
rect 54547 56254 54605 56260
rect 1744 56217 1750 56229
rect 1705 56189 1750 56217
rect 1744 56177 1750 56189
rect 1802 56177 1808 56229
rect 2992 56177 2998 56229
rect 3050 56217 3056 56229
rect 4243 56220 4301 56226
rect 3050 56189 3095 56217
rect 3050 56177 3056 56189
rect 4243 56186 4255 56220
rect 4289 56217 4301 56220
rect 4531 56220 4589 56226
rect 4531 56217 4543 56220
rect 4289 56189 4543 56217
rect 4289 56186 4301 56189
rect 4243 56180 4301 56186
rect 4531 56186 4543 56189
rect 4577 56217 4589 56220
rect 4720 56217 4726 56229
rect 4577 56189 4726 56217
rect 4577 56186 4589 56189
rect 4531 56180 4589 56186
rect 4720 56177 4726 56189
rect 4778 56177 4784 56229
rect 5584 56217 5590 56229
rect 5545 56189 5590 56217
rect 5584 56177 5590 56189
rect 5642 56177 5648 56229
rect 6352 56217 6358 56229
rect 6313 56189 6358 56217
rect 6352 56177 6358 56189
rect 6410 56177 6416 56229
rect 7216 56177 7222 56229
rect 7274 56217 7280 56229
rect 7274 56189 7319 56217
rect 7274 56177 7280 56189
rect 8560 56177 8566 56229
rect 8618 56217 8624 56229
rect 10096 56217 10102 56229
rect 8618 56189 8663 56217
rect 10057 56189 10102 56217
rect 8618 56177 8624 56189
rect 10096 56177 10102 56189
rect 10154 56217 10160 56229
rect 10387 56220 10445 56226
rect 10387 56217 10399 56220
rect 10154 56189 10399 56217
rect 10154 56177 10160 56189
rect 10387 56186 10399 56189
rect 10433 56186 10445 56220
rect 11152 56217 11158 56229
rect 11113 56189 11158 56217
rect 10387 56180 10445 56186
rect 11152 56177 11158 56189
rect 11210 56177 11216 56229
rect 11635 56220 11693 56226
rect 11635 56186 11647 56220
rect 11681 56217 11693 56220
rect 11920 56217 11926 56229
rect 11681 56189 11926 56217
rect 11681 56186 11693 56189
rect 11635 56180 11693 56186
rect 11920 56177 11926 56189
rect 11978 56177 11984 56229
rect 12304 56217 12310 56229
rect 12265 56189 12310 56217
rect 12304 56177 12310 56189
rect 12362 56217 12368 56229
rect 12691 56220 12749 56226
rect 12691 56217 12703 56220
rect 12362 56189 12703 56217
rect 12362 56177 12368 56189
rect 12691 56186 12703 56189
rect 12737 56186 12749 56220
rect 12691 56180 12749 56186
rect 13552 56177 13558 56229
rect 13610 56217 13616 56229
rect 15091 56220 15149 56226
rect 13610 56189 13655 56217
rect 13610 56177 13616 56189
rect 15091 56186 15103 56220
rect 15137 56217 15149 56220
rect 15184 56217 15190 56229
rect 15137 56189 15190 56217
rect 15137 56186 15149 56189
rect 15091 56180 15149 56186
rect 15184 56177 15190 56189
rect 15242 56177 15248 56229
rect 15280 56177 15286 56229
rect 15338 56217 15344 56229
rect 15859 56220 15917 56226
rect 15859 56217 15871 56220
rect 15338 56189 15871 56217
rect 15338 56177 15344 56189
rect 15859 56186 15871 56189
rect 15905 56186 15917 56220
rect 16816 56217 16822 56229
rect 16777 56189 16822 56217
rect 15859 56180 15917 56186
rect 16816 56177 16822 56189
rect 16874 56217 16880 56229
rect 17203 56220 17261 56226
rect 17203 56217 17215 56220
rect 16874 56189 17215 56217
rect 16874 56177 16880 56189
rect 17203 56186 17215 56189
rect 17249 56186 17261 56220
rect 17203 56180 17261 56186
rect 18064 56177 18070 56229
rect 18122 56217 18128 56229
rect 18739 56220 18797 56226
rect 18739 56217 18751 56220
rect 18122 56189 18751 56217
rect 18122 56177 18128 56189
rect 18739 56186 18751 56189
rect 18785 56186 18797 56220
rect 20368 56217 20374 56229
rect 20329 56189 20374 56217
rect 18739 56180 18797 56186
rect 20368 56177 20374 56189
rect 20426 56177 20432 56229
rect 21424 56217 21430 56229
rect 21385 56189 21430 56217
rect 21424 56177 21430 56189
rect 21482 56177 21488 56229
rect 21907 56220 21965 56226
rect 21907 56186 21919 56220
rect 21953 56217 21965 56220
rect 22096 56217 22102 56229
rect 21953 56189 22102 56217
rect 21953 56186 21965 56189
rect 21907 56180 21965 56186
rect 22096 56177 22102 56189
rect 22154 56177 22160 56229
rect 22672 56177 22678 56229
rect 22730 56217 22736 56229
rect 22963 56220 23021 56226
rect 22963 56217 22975 56220
rect 22730 56189 22975 56217
rect 22730 56177 22736 56189
rect 22963 56186 22975 56189
rect 23009 56186 23021 56220
rect 24400 56217 24406 56229
rect 24361 56189 24406 56217
rect 22963 56180 23021 56186
rect 24400 56177 24406 56189
rect 24458 56177 24464 56229
rect 26128 56217 26134 56229
rect 26089 56189 26134 56217
rect 26128 56177 26134 56189
rect 26186 56177 26192 56229
rect 27760 56217 27766 56229
rect 27721 56189 27766 56217
rect 27760 56177 27766 56189
rect 27818 56177 27824 56229
rect 28243 56220 28301 56226
rect 28243 56186 28255 56220
rect 28289 56217 28301 56220
rect 28432 56217 28438 56229
rect 28289 56189 28438 56217
rect 28289 56186 28301 56189
rect 28243 56180 28301 56186
rect 28432 56177 28438 56189
rect 28490 56177 28496 56229
rect 29395 56220 29453 56226
rect 29395 56186 29407 56220
rect 29441 56217 29453 56220
rect 29584 56217 29590 56229
rect 29441 56189 29590 56217
rect 29441 56186 29453 56189
rect 29395 56180 29453 56186
rect 29584 56177 29590 56189
rect 29642 56177 29648 56229
rect 30928 56217 30934 56229
rect 30889 56189 30934 56217
rect 30928 56177 30934 56189
rect 30986 56177 30992 56229
rect 32464 56217 32470 56229
rect 32425 56189 32470 56217
rect 32464 56177 32470 56189
rect 32522 56177 32528 56229
rect 33715 56220 33773 56226
rect 33715 56186 33727 56220
rect 33761 56217 33773 56220
rect 34003 56220 34061 56226
rect 34003 56217 34015 56220
rect 33761 56189 34015 56217
rect 33761 56186 33773 56189
rect 33715 56180 33773 56186
rect 34003 56186 34015 56189
rect 34049 56217 34061 56220
rect 34192 56217 34198 56229
rect 34049 56189 34198 56217
rect 34049 56186 34061 56189
rect 34003 56180 34061 56186
rect 34192 56177 34198 56189
rect 34250 56177 34256 56229
rect 34384 56217 34390 56229
rect 34345 56189 34390 56217
rect 34384 56177 34390 56189
rect 34442 56217 34448 56229
rect 34675 56220 34733 56226
rect 34675 56217 34687 56220
rect 34442 56189 34687 56217
rect 34442 56177 34448 56189
rect 34675 56186 34687 56189
rect 34721 56217 34733 56220
rect 34963 56220 35021 56226
rect 34963 56217 34975 56220
rect 34721 56189 34975 56217
rect 34721 56186 34733 56189
rect 34675 56180 34733 56186
rect 34963 56186 34975 56189
rect 35009 56186 35021 56220
rect 34963 56180 35021 56186
rect 36208 56177 36214 56229
rect 36266 56217 36272 56229
rect 36592 56217 36598 56229
rect 36266 56189 36311 56217
rect 36553 56189 36598 56217
rect 36266 56177 36272 56189
rect 36592 56177 36598 56189
rect 36650 56217 36656 56229
rect 36883 56220 36941 56226
rect 36883 56217 36895 56220
rect 36650 56189 36895 56217
rect 36650 56177 36656 56189
rect 36883 56186 36895 56189
rect 36929 56186 36941 56220
rect 36883 56180 36941 56186
rect 37459 56220 37517 56226
rect 37459 56186 37471 56220
rect 37505 56217 37517 56220
rect 37744 56217 37750 56229
rect 37505 56189 37750 56217
rect 37505 56186 37517 56189
rect 37459 56180 37517 56186
rect 37744 56177 37750 56189
rect 37802 56177 37808 56229
rect 38515 56220 38573 56226
rect 38515 56186 38527 56220
rect 38561 56217 38573 56220
rect 38704 56217 38710 56229
rect 38561 56189 38710 56217
rect 38561 56186 38573 56189
rect 38515 56180 38573 56186
rect 38704 56177 38710 56189
rect 38762 56177 38768 56229
rect 38800 56177 38806 56229
rect 38858 56217 38864 56229
rect 40243 56220 40301 56226
rect 40243 56217 40255 56220
rect 38858 56189 40255 56217
rect 38858 56177 38864 56189
rect 40243 56186 40255 56189
rect 40289 56186 40301 56220
rect 41584 56217 41590 56229
rect 41545 56189 41590 56217
rect 40243 56180 40301 56186
rect 41584 56177 41590 56189
rect 41642 56217 41648 56229
rect 41875 56220 41933 56226
rect 41875 56217 41887 56220
rect 41642 56189 41887 56217
rect 41642 56177 41648 56189
rect 41875 56186 41887 56189
rect 41921 56186 41933 56220
rect 41875 56180 41933 56186
rect 42643 56220 42701 56226
rect 42643 56186 42655 56220
rect 42689 56186 42701 56220
rect 42643 56180 42701 56186
rect 43219 56220 43277 56226
rect 43219 56186 43231 56220
rect 43265 56217 43277 56220
rect 43408 56217 43414 56229
rect 43265 56189 43414 56217
rect 43265 56186 43277 56189
rect 43219 56180 43277 56186
rect 2224 56103 2230 56155
rect 2282 56143 2288 56155
rect 5776 56143 5782 56155
rect 2282 56115 5782 56143
rect 2282 56103 2288 56115
rect 5776 56103 5782 56115
rect 5834 56103 5840 56155
rect 18160 56103 18166 56155
rect 18218 56143 18224 56155
rect 21808 56143 21814 56155
rect 18218 56115 21814 56143
rect 18218 56103 18224 56115
rect 21808 56103 21814 56115
rect 21866 56103 21872 56155
rect 37072 56103 37078 56155
rect 37130 56143 37136 56155
rect 40336 56143 40342 56155
rect 37130 56115 40342 56143
rect 37130 56103 37136 56115
rect 40336 56103 40342 56115
rect 40394 56103 40400 56155
rect 40720 56103 40726 56155
rect 40778 56143 40784 56155
rect 42658 56143 42686 56180
rect 43408 56177 43414 56189
rect 43466 56177 43472 56229
rect 43888 56217 43894 56229
rect 43849 56189 43894 56217
rect 43888 56177 43894 56189
rect 43946 56217 43952 56229
rect 44179 56220 44237 56226
rect 44179 56217 44191 56220
rect 43946 56189 44191 56217
rect 43946 56177 43952 56189
rect 44179 56186 44191 56189
rect 44225 56186 44237 56220
rect 44752 56217 44758 56229
rect 44713 56189 44758 56217
rect 44179 56180 44237 56186
rect 44752 56177 44758 56189
rect 44810 56217 44816 56229
rect 45139 56220 45197 56226
rect 45139 56217 45151 56220
rect 44810 56189 45151 56217
rect 44810 56177 44816 56189
rect 45139 56186 45151 56189
rect 45185 56186 45197 56220
rect 46768 56217 46774 56229
rect 46729 56189 46774 56217
rect 45139 56180 45197 56186
rect 46768 56177 46774 56189
rect 46826 56177 46832 56229
rect 47824 56217 47830 56229
rect 47785 56189 47830 56217
rect 47824 56177 47830 56189
rect 47882 56217 47888 56229
rect 48115 56220 48173 56226
rect 48115 56217 48127 56220
rect 47882 56189 48127 56217
rect 47882 56177 47888 56189
rect 48115 56186 48127 56189
rect 48161 56217 48173 56220
rect 48403 56220 48461 56226
rect 48403 56217 48415 56220
rect 48161 56189 48415 56217
rect 48161 56186 48173 56189
rect 48115 56180 48173 56186
rect 48403 56186 48415 56189
rect 48449 56186 48461 56220
rect 48592 56217 48598 56229
rect 48553 56189 48598 56217
rect 48403 56180 48461 56186
rect 48592 56177 48598 56189
rect 48650 56217 48656 56229
rect 48883 56220 48941 56226
rect 48883 56217 48895 56220
rect 48650 56189 48895 56217
rect 48650 56177 48656 56189
rect 48883 56186 48895 56189
rect 48929 56186 48941 56220
rect 50224 56217 50230 56229
rect 50185 56189 50230 56217
rect 48883 56180 48941 56186
rect 50224 56177 50230 56189
rect 50282 56217 50288 56229
rect 50515 56220 50573 56226
rect 50515 56217 50527 56220
rect 50282 56189 50527 56217
rect 50282 56177 50288 56189
rect 50515 56186 50527 56189
rect 50561 56186 50573 56220
rect 51664 56217 51670 56229
rect 51625 56189 51670 56217
rect 50515 56180 50573 56186
rect 51664 56177 51670 56189
rect 51722 56217 51728 56229
rect 51955 56220 52013 56226
rect 51955 56217 51967 56220
rect 51722 56189 51967 56217
rect 51722 56177 51728 56189
rect 51955 56186 51967 56189
rect 52001 56186 52013 56220
rect 51955 56180 52013 56186
rect 52051 56220 52109 56226
rect 52051 56186 52063 56220
rect 52097 56186 52109 56220
rect 53392 56217 53398 56229
rect 53353 56189 53398 56217
rect 52051 56180 52109 56186
rect 40778 56115 42686 56143
rect 40778 56103 40784 56115
rect 51184 56103 51190 56155
rect 51242 56143 51248 56155
rect 52066 56143 52094 56180
rect 53392 56177 53398 56189
rect 53450 56217 53456 56229
rect 53683 56220 53741 56226
rect 53683 56217 53695 56220
rect 53450 56189 53695 56217
rect 53450 56177 53456 56189
rect 53683 56186 53695 56189
rect 53729 56186 53741 56220
rect 57586 56217 57614 56263
rect 57811 56260 57823 56294
rect 57857 56291 57869 56294
rect 58576 56291 58582 56303
rect 57857 56263 58582 56291
rect 57857 56260 57869 56263
rect 57811 56254 57869 56260
rect 58576 56251 58582 56263
rect 58634 56251 58640 56303
rect 58192 56217 58198 56229
rect 57586 56189 58198 56217
rect 53683 56180 53741 56186
rect 58192 56177 58198 56189
rect 58250 56177 58256 56229
rect 51242 56115 52094 56143
rect 51242 56103 51248 56115
rect 1152 55970 58848 55992
rect 1152 55918 4294 55970
rect 4346 55918 4358 55970
rect 4410 55918 4422 55970
rect 4474 55918 4486 55970
rect 4538 55918 35014 55970
rect 35066 55918 35078 55970
rect 35130 55918 35142 55970
rect 35194 55918 35206 55970
rect 35258 55918 58848 55970
rect 1152 55896 58848 55918
rect 36112 55807 36118 55859
rect 36170 55847 36176 55859
rect 36170 55819 39950 55847
rect 36170 55807 36176 55819
rect 38896 55733 38902 55785
rect 38954 55733 38960 55785
rect 1168 55659 1174 55711
rect 1226 55699 1232 55711
rect 1651 55702 1709 55708
rect 1651 55699 1663 55702
rect 1226 55671 1663 55699
rect 1226 55659 1232 55671
rect 1651 55668 1663 55671
rect 1697 55668 1709 55702
rect 1651 55662 1709 55668
rect 4435 55702 4493 55708
rect 4435 55668 4447 55702
rect 4481 55699 4493 55702
rect 4624 55699 4630 55711
rect 4481 55671 4630 55699
rect 4481 55668 4493 55671
rect 4435 55662 4493 55668
rect 4624 55659 4630 55671
rect 4682 55659 4688 55711
rect 7504 55659 7510 55711
rect 7562 55699 7568 55711
rect 7603 55702 7661 55708
rect 7603 55699 7615 55702
rect 7562 55671 7615 55699
rect 7562 55659 7568 55671
rect 7603 55668 7615 55671
rect 7649 55668 7661 55702
rect 7603 55662 7661 55668
rect 9136 55659 9142 55711
rect 9194 55699 9200 55711
rect 9235 55702 9293 55708
rect 9235 55699 9247 55702
rect 9194 55671 9247 55699
rect 9194 55659 9200 55671
rect 9235 55668 9247 55671
rect 9281 55668 9293 55702
rect 9235 55662 9293 55668
rect 13840 55659 13846 55711
rect 13898 55699 13904 55711
rect 14035 55702 14093 55708
rect 14035 55699 14047 55702
rect 13898 55671 14047 55699
rect 13898 55659 13904 55671
rect 14035 55668 14047 55671
rect 14081 55668 14093 55702
rect 14035 55662 14093 55668
rect 20176 55659 20182 55711
rect 20234 55699 20240 55711
rect 20275 55702 20333 55708
rect 20275 55699 20287 55702
rect 20234 55671 20287 55699
rect 20234 55659 20240 55671
rect 20275 55668 20287 55671
rect 20321 55668 20333 55702
rect 20275 55662 20333 55668
rect 23344 55659 23350 55711
rect 23402 55699 23408 55711
rect 23539 55702 23597 55708
rect 23539 55699 23551 55702
rect 23402 55671 23551 55699
rect 23402 55659 23408 55671
rect 23539 55668 23551 55671
rect 23585 55668 23597 55702
rect 23539 55662 23597 55668
rect 24880 55659 24886 55711
rect 24938 55699 24944 55711
rect 24979 55702 25037 55708
rect 24979 55699 24991 55702
rect 24938 55671 24991 55699
rect 24938 55659 24944 55671
rect 24979 55668 24991 55671
rect 25025 55668 25037 55702
rect 39922 55685 39950 55819
rect 41776 55807 41782 55859
rect 41834 55807 41840 55859
rect 41794 55773 41822 55807
rect 41760 55745 41822 55773
rect 24979 55662 25037 55668
rect 42256 55659 42262 55711
rect 42314 55699 42320 55711
rect 42451 55702 42509 55708
rect 42451 55699 42463 55702
rect 42314 55671 42463 55699
rect 42314 55659 42320 55671
rect 42451 55668 42463 55671
rect 42497 55668 42509 55702
rect 42451 55662 42509 55668
rect 45424 55659 45430 55711
rect 45482 55699 45488 55711
rect 45619 55702 45677 55708
rect 45619 55699 45631 55702
rect 45482 55671 45631 55699
rect 45482 55659 45488 55671
rect 45619 55668 45631 55671
rect 45665 55668 45677 55702
rect 45619 55662 45677 55668
rect 46960 55659 46966 55711
rect 47018 55699 47024 55711
rect 47155 55702 47213 55708
rect 47155 55699 47167 55702
rect 47018 55671 47167 55699
rect 47018 55659 47024 55671
rect 47155 55668 47167 55671
rect 47201 55668 47213 55702
rect 47155 55662 47213 55668
rect 51760 55659 51766 55711
rect 51818 55699 51824 55711
rect 51859 55702 51917 55708
rect 51859 55699 51871 55702
rect 51818 55671 51871 55699
rect 51818 55659 51824 55671
rect 51859 55668 51871 55671
rect 51905 55668 51917 55702
rect 51859 55662 51917 55668
rect 56464 55659 56470 55711
rect 56522 55699 56528 55711
rect 56563 55702 56621 55708
rect 56563 55699 56575 55702
rect 56522 55671 56575 55699
rect 56522 55659 56528 55671
rect 56563 55668 56575 55671
rect 56609 55668 56621 55702
rect 56563 55662 56621 55668
rect 57520 55659 57526 55711
rect 57578 55699 57584 55711
rect 57715 55702 57773 55708
rect 57715 55699 57727 55702
rect 57578 55671 57727 55699
rect 57578 55659 57584 55671
rect 57715 55668 57727 55671
rect 57761 55668 57773 55702
rect 57715 55662 57773 55668
rect 1747 55554 1805 55560
rect 1747 55520 1759 55554
rect 1793 55520 1805 55554
rect 1747 55514 1805 55520
rect 4531 55554 4589 55560
rect 4531 55520 4543 55554
rect 4577 55551 4589 55554
rect 5392 55551 5398 55563
rect 4577 55523 5398 55551
rect 4577 55520 4589 55523
rect 4531 55514 4589 55520
rect 1762 55403 1790 55514
rect 5392 55511 5398 55523
rect 5450 55511 5456 55563
rect 7411 55554 7469 55560
rect 7411 55520 7423 55554
rect 7457 55551 7469 55554
rect 7696 55551 7702 55563
rect 7457 55523 7702 55551
rect 7457 55520 7469 55523
rect 7411 55514 7469 55520
rect 7696 55511 7702 55523
rect 7754 55511 7760 55563
rect 9328 55551 9334 55563
rect 9289 55523 9334 55551
rect 9328 55511 9334 55523
rect 9386 55511 9392 55563
rect 12115 55554 12173 55560
rect 12115 55520 12127 55554
rect 12161 55551 12173 55554
rect 12400 55551 12406 55563
rect 12161 55523 12406 55551
rect 12161 55520 12173 55523
rect 12115 55514 12173 55520
rect 12400 55511 12406 55523
rect 12458 55511 12464 55563
rect 13939 55554 13997 55560
rect 13939 55551 13951 55554
rect 13858 55523 13951 55551
rect 13858 55415 13886 55523
rect 13939 55520 13951 55523
rect 13985 55520 13997 55554
rect 13939 55514 13997 55520
rect 20371 55554 20429 55560
rect 20371 55520 20383 55554
rect 20417 55551 20429 55554
rect 20464 55551 20470 55563
rect 20417 55523 20470 55551
rect 20417 55520 20429 55523
rect 20371 55514 20429 55520
rect 20464 55511 20470 55523
rect 20522 55511 20528 55563
rect 23443 55554 23501 55560
rect 23443 55551 23455 55554
rect 23170 55523 23455 55551
rect 23170 55415 23198 55523
rect 23443 55520 23455 55523
rect 23489 55520 23501 55554
rect 23443 55514 23501 55520
rect 24787 55554 24845 55560
rect 24787 55520 24799 55554
rect 24833 55551 24845 55554
rect 25072 55551 25078 55563
rect 24833 55523 25078 55551
rect 24833 55520 24845 55523
rect 24787 55514 24845 55520
rect 25072 55511 25078 55523
rect 25130 55511 25136 55563
rect 42544 55551 42550 55563
rect 42505 55523 42550 55551
rect 42544 55511 42550 55523
rect 42602 55511 42608 55563
rect 45331 55554 45389 55560
rect 45331 55520 45343 55554
rect 45377 55551 45389 55554
rect 45520 55551 45526 55563
rect 45377 55523 45526 55551
rect 45377 55520 45389 55523
rect 45331 55514 45389 55520
rect 45520 55511 45526 55523
rect 45578 55511 45584 55563
rect 47059 55554 47117 55560
rect 47059 55551 47071 55554
rect 46978 55523 47071 55551
rect 46978 55415 47006 55523
rect 47059 55520 47071 55523
rect 47105 55551 47117 55554
rect 47347 55554 47405 55560
rect 47347 55551 47359 55554
rect 47105 55523 47359 55551
rect 47105 55520 47117 55523
rect 47059 55514 47117 55520
rect 47347 55520 47359 55523
rect 47393 55520 47405 55554
rect 47347 55514 47405 55520
rect 51955 55554 52013 55560
rect 51955 55520 51967 55554
rect 52001 55551 52013 55554
rect 52048 55551 52054 55563
rect 52001 55523 52054 55551
rect 52001 55520 52013 55523
rect 51955 55514 52013 55520
rect 52048 55511 52054 55523
rect 52106 55511 52112 55563
rect 55795 55554 55853 55560
rect 55795 55520 55807 55554
rect 55841 55520 55853 55554
rect 55795 55514 55853 55520
rect 2032 55403 2038 55415
rect 1762 55375 2038 55403
rect 2032 55363 2038 55375
rect 2090 55363 2096 55415
rect 13747 55406 13805 55412
rect 13747 55372 13759 55406
rect 13793 55403 13805 55406
rect 13840 55403 13846 55415
rect 13793 55375 13846 55403
rect 13793 55372 13805 55375
rect 13747 55366 13805 55372
rect 13840 55363 13846 55375
rect 13898 55363 13904 55415
rect 23152 55403 23158 55415
rect 23113 55375 23158 55403
rect 23152 55363 23158 55375
rect 23210 55363 23216 55415
rect 39760 55363 39766 55415
rect 39818 55363 39824 55415
rect 46867 55406 46925 55412
rect 46867 55372 46879 55406
rect 46913 55403 46925 55406
rect 46960 55403 46966 55415
rect 46913 55375 46966 55403
rect 46913 55372 46925 55375
rect 46867 55366 46925 55372
rect 46960 55363 46966 55375
rect 47018 55363 47024 55415
rect 55600 55403 55606 55415
rect 55561 55375 55606 55403
rect 55600 55363 55606 55375
rect 55658 55403 55664 55415
rect 55810 55403 55838 55514
rect 55888 55511 55894 55563
rect 55946 55551 55952 55563
rect 56659 55554 56717 55560
rect 56659 55551 56671 55554
rect 55946 55523 56671 55551
rect 55946 55511 55952 55523
rect 56659 55520 56671 55523
rect 56705 55520 56717 55554
rect 57619 55554 57677 55560
rect 57619 55551 57631 55554
rect 56659 55514 56717 55520
rect 57346 55523 57631 55551
rect 57346 55415 57374 55523
rect 57619 55520 57631 55523
rect 57665 55551 57677 55554
rect 57907 55554 57965 55560
rect 57907 55551 57919 55554
rect 57665 55523 57919 55551
rect 57665 55520 57677 55523
rect 57619 55514 57677 55520
rect 57907 55520 57919 55523
rect 57953 55520 57965 55554
rect 57907 55514 57965 55520
rect 57328 55403 57334 55415
rect 55658 55375 55838 55403
rect 57289 55375 57334 55403
rect 55658 55363 55664 55375
rect 57328 55363 57334 55375
rect 57386 55363 57392 55415
rect 1152 55304 58848 55326
rect 1152 55252 19654 55304
rect 19706 55252 19718 55304
rect 19770 55252 19782 55304
rect 19834 55252 19846 55304
rect 19898 55252 50374 55304
rect 50426 55252 50438 55304
rect 50490 55252 50502 55304
rect 50554 55252 50566 55304
rect 50618 55252 58848 55304
rect 1152 55230 58848 55252
rect 12400 55141 12406 55193
rect 12458 55181 12464 55193
rect 28336 55181 28342 55193
rect 12458 55153 28342 55181
rect 12458 55141 12464 55153
rect 28336 55141 28342 55153
rect 28394 55141 28400 55193
rect 39088 55141 39094 55193
rect 39146 55181 39152 55193
rect 39187 55184 39245 55190
rect 39187 55181 39199 55184
rect 39146 55153 39199 55181
rect 39146 55141 39152 55153
rect 39187 55150 39199 55153
rect 39233 55150 39245 55184
rect 39187 55144 39245 55150
rect 57811 55184 57869 55190
rect 57811 55150 57823 55184
rect 57857 55181 57869 55184
rect 59152 55181 59158 55193
rect 57857 55153 59158 55181
rect 57857 55150 57869 55153
rect 57811 55144 57869 55150
rect 59152 55141 59158 55153
rect 59210 55141 59216 55193
rect 2032 54993 2038 55045
rect 2090 55033 2096 55045
rect 55600 55033 55606 55045
rect 2090 55005 55606 55033
rect 2090 54993 2096 55005
rect 55600 54993 55606 55005
rect 55658 54993 55664 55045
rect 39280 54845 39286 54897
rect 39338 54885 39344 54897
rect 39338 54857 39383 54885
rect 39338 54845 39344 54857
rect 57904 54845 57910 54897
rect 57962 54885 57968 54897
rect 57962 54857 58007 54885
rect 57962 54845 57968 54857
rect 53968 54771 53974 54823
rect 54026 54811 54032 54823
rect 55603 54814 55661 54820
rect 55603 54811 55615 54814
rect 54026 54783 55615 54811
rect 54026 54771 54032 54783
rect 55603 54780 55615 54783
rect 55649 54811 55661 54814
rect 55795 54814 55853 54820
rect 55795 54811 55807 54814
rect 55649 54783 55807 54811
rect 55649 54780 55661 54783
rect 55603 54774 55661 54780
rect 55795 54780 55807 54783
rect 55841 54780 55853 54814
rect 55795 54774 55853 54780
rect 35824 54737 35830 54749
rect 35785 54709 35830 54737
rect 35824 54697 35830 54709
rect 35882 54737 35888 54749
rect 36019 54740 36077 54746
rect 36019 54737 36031 54740
rect 35882 54709 36031 54737
rect 35882 54697 35888 54709
rect 36019 54706 36031 54709
rect 36065 54706 36077 54740
rect 36019 54700 36077 54706
rect 39763 54740 39821 54746
rect 39763 54706 39775 54740
rect 39809 54737 39821 54740
rect 39856 54737 39862 54749
rect 39809 54709 39862 54737
rect 39809 54706 39821 54709
rect 39763 54700 39821 54706
rect 39856 54697 39862 54709
rect 39914 54697 39920 54749
rect 53872 54737 53878 54749
rect 53833 54709 53878 54737
rect 53872 54697 53878 54709
rect 53930 54737 53936 54749
rect 54067 54740 54125 54746
rect 54067 54737 54079 54740
rect 53930 54709 54079 54737
rect 53930 54697 53936 54709
rect 54067 54706 54079 54709
rect 54113 54706 54125 54740
rect 54067 54700 54125 54706
rect 1152 54638 58848 54660
rect 1152 54586 4294 54638
rect 4346 54586 4358 54638
rect 4410 54586 4422 54638
rect 4474 54586 4486 54638
rect 4538 54586 35014 54638
rect 35066 54586 35078 54638
rect 35130 54586 35142 54638
rect 35194 54586 35206 54638
rect 35258 54586 58848 54638
rect 1152 54564 58848 54586
rect 11152 54475 11158 54527
rect 11210 54515 11216 54527
rect 42643 54518 42701 54524
rect 42643 54515 42655 54518
rect 11210 54487 42655 54515
rect 11210 54475 11216 54487
rect 42643 54484 42655 54487
rect 42689 54484 42701 54518
rect 42643 54478 42701 54484
rect 57811 54370 57869 54376
rect 57811 54336 57823 54370
rect 57857 54367 57869 54370
rect 58096 54367 58102 54379
rect 57857 54339 58102 54367
rect 57857 54336 57869 54339
rect 57811 54330 57869 54336
rect 58096 54327 58102 54339
rect 58154 54327 58160 54379
rect 31216 54179 31222 54231
rect 31274 54219 31280 54231
rect 34498 54219 34526 54316
rect 31274 54191 34526 54219
rect 31274 54179 31280 54191
rect 35026 54145 35054 54316
rect 36499 54222 36557 54228
rect 36499 54219 36511 54222
rect 33922 54117 35054 54145
rect 36322 54191 36511 54219
rect 31120 54031 31126 54083
rect 31178 54071 31184 54083
rect 33922 54080 33950 54117
rect 36322 54083 36350 54191
rect 36499 54188 36511 54191
rect 36545 54188 36557 54222
rect 36499 54182 36557 54188
rect 57808 54179 57814 54231
rect 57866 54219 57872 54231
rect 57907 54222 57965 54228
rect 57907 54219 57919 54222
rect 57866 54191 57919 54219
rect 57866 54179 57872 54191
rect 57907 54188 57919 54191
rect 57953 54188 57965 54222
rect 57907 54182 57965 54188
rect 33907 54074 33965 54080
rect 33907 54071 33919 54074
rect 31178 54043 33919 54071
rect 31178 54031 31184 54043
rect 33907 54040 33919 54043
rect 33953 54040 33965 54074
rect 33907 54034 33965 54040
rect 34864 54031 34870 54083
rect 34922 54031 34928 54083
rect 36304 54071 36310 54083
rect 36265 54043 36310 54071
rect 36304 54031 36310 54043
rect 36362 54031 36368 54083
rect 1152 53972 58848 53994
rect 1152 53920 19654 53972
rect 19706 53920 19718 53972
rect 19770 53920 19782 53972
rect 19834 53920 19846 53972
rect 19898 53920 50374 53972
rect 50426 53920 50438 53972
rect 50490 53920 50502 53972
rect 50554 53920 50566 53972
rect 50618 53920 58848 53972
rect 1152 53898 58848 53920
rect 57907 53852 57965 53858
rect 57907 53818 57919 53852
rect 57953 53849 57965 53852
rect 59632 53849 59638 53861
rect 57953 53821 59638 53849
rect 57953 53818 57965 53821
rect 57907 53812 57965 53818
rect 59632 53809 59638 53821
rect 59690 53809 59696 53861
rect 25552 53513 25558 53565
rect 25610 53553 25616 53565
rect 57619 53556 57677 53562
rect 57619 53553 57631 53556
rect 25610 53525 57631 53553
rect 25610 53513 25616 53525
rect 57619 53522 57631 53525
rect 57665 53553 57677 53556
rect 57811 53556 57869 53562
rect 57811 53553 57823 53556
rect 57665 53525 57823 53553
rect 57665 53522 57677 53525
rect 57619 53516 57677 53522
rect 57811 53522 57823 53525
rect 57857 53522 57869 53556
rect 57811 53516 57869 53522
rect 22291 53408 22349 53414
rect 22291 53374 22303 53408
rect 22337 53405 22349 53408
rect 22579 53408 22637 53414
rect 22579 53405 22591 53408
rect 22337 53377 22591 53405
rect 22337 53374 22349 53377
rect 22291 53368 22349 53374
rect 22579 53374 22591 53377
rect 22625 53405 22637 53408
rect 26608 53405 26614 53417
rect 22625 53377 26614 53405
rect 22625 53374 22637 53377
rect 22579 53368 22637 53374
rect 26608 53365 26614 53377
rect 26666 53365 26672 53417
rect 44947 53408 45005 53414
rect 44947 53374 44959 53408
rect 44993 53405 45005 53408
rect 45235 53408 45293 53414
rect 45235 53405 45247 53408
rect 44993 53377 45247 53405
rect 44993 53374 45005 53377
rect 44947 53368 45005 53374
rect 45235 53374 45247 53377
rect 45281 53405 45293 53408
rect 49648 53405 49654 53417
rect 45281 53377 49654 53405
rect 45281 53374 45293 53377
rect 45235 53368 45293 53374
rect 49648 53365 49654 53377
rect 49706 53365 49712 53417
rect 1152 53306 58848 53328
rect 1152 53254 4294 53306
rect 4346 53254 4358 53306
rect 4410 53254 4422 53306
rect 4474 53254 4486 53306
rect 4538 53254 35014 53306
rect 35066 53254 35078 53306
rect 35130 53254 35142 53306
rect 35194 53254 35206 53306
rect 35258 53254 58848 53306
rect 1152 53232 58848 53254
rect 29395 52890 29453 52896
rect 29395 52856 29407 52890
rect 29441 52887 29453 52890
rect 29683 52890 29741 52896
rect 29683 52887 29695 52890
rect 29441 52859 29695 52887
rect 29441 52856 29453 52859
rect 29395 52850 29453 52856
rect 29683 52856 29695 52859
rect 29729 52856 29741 52890
rect 56179 52890 56237 52896
rect 56179 52887 56191 52890
rect 29683 52850 29741 52856
rect 37426 52859 56191 52887
rect 17008 52773 17014 52825
rect 17066 52813 17072 52825
rect 37426 52813 37454 52859
rect 56179 52856 56191 52859
rect 56225 52887 56237 52890
rect 56275 52890 56333 52896
rect 56275 52887 56287 52890
rect 56225 52859 56287 52887
rect 56225 52856 56237 52859
rect 56179 52850 56237 52856
rect 56275 52856 56287 52859
rect 56321 52856 56333 52890
rect 56275 52850 56333 52856
rect 17066 52785 37454 52813
rect 17066 52773 17072 52785
rect 16336 52699 16342 52751
rect 16394 52739 16400 52751
rect 29395 52742 29453 52748
rect 29395 52739 29407 52742
rect 16394 52711 29407 52739
rect 16394 52699 16400 52711
rect 29395 52708 29407 52711
rect 29441 52739 29453 52742
rect 29491 52742 29549 52748
rect 29491 52739 29503 52742
rect 29441 52711 29503 52739
rect 29441 52708 29453 52711
rect 29395 52702 29453 52708
rect 29491 52708 29503 52711
rect 29537 52708 29549 52742
rect 29491 52702 29549 52708
rect 1152 52640 58848 52662
rect 1152 52588 19654 52640
rect 19706 52588 19718 52640
rect 19770 52588 19782 52640
rect 19834 52588 19846 52640
rect 19898 52588 50374 52640
rect 50426 52588 50438 52640
rect 50490 52588 50502 52640
rect 50554 52588 50566 52640
rect 50618 52588 58848 52640
rect 1152 52566 58848 52588
rect 19987 52150 20045 52156
rect 19987 52147 19999 52150
rect 7186 52119 19999 52147
rect 2128 52033 2134 52085
rect 2186 52073 2192 52085
rect 7186 52073 7214 52119
rect 19987 52116 19999 52119
rect 20033 52147 20045 52150
rect 20179 52150 20237 52156
rect 20179 52147 20191 52150
rect 20033 52119 20191 52147
rect 20033 52116 20045 52119
rect 19987 52110 20045 52116
rect 20179 52116 20191 52119
rect 20225 52116 20237 52150
rect 20179 52110 20237 52116
rect 2186 52045 7214 52073
rect 17683 52076 17741 52082
rect 2186 52033 2192 52045
rect 17683 52042 17695 52076
rect 17729 52073 17741 52076
rect 17971 52076 18029 52082
rect 17971 52073 17983 52076
rect 17729 52045 17983 52073
rect 17729 52042 17741 52045
rect 17683 52036 17741 52042
rect 17971 52042 17983 52045
rect 18017 52073 18029 52076
rect 22192 52073 22198 52085
rect 18017 52045 22198 52073
rect 18017 52042 18029 52045
rect 17971 52036 18029 52042
rect 22192 52033 22198 52045
rect 22250 52033 22256 52085
rect 32371 52076 32429 52082
rect 32371 52042 32383 52076
rect 32417 52073 32429 52076
rect 32656 52073 32662 52085
rect 32417 52045 32662 52073
rect 32417 52042 32429 52045
rect 32371 52036 32429 52042
rect 32656 52033 32662 52045
rect 32714 52033 32720 52085
rect 1152 51974 58848 51996
rect 1152 51922 4294 51974
rect 4346 51922 4358 51974
rect 4410 51922 4422 51974
rect 4474 51922 4486 51974
rect 4538 51922 35014 51974
rect 35066 51922 35078 51974
rect 35130 51922 35142 51974
rect 35194 51922 35206 51974
rect 35258 51922 58848 51974
rect 1152 51900 58848 51922
rect 13459 51632 13517 51638
rect 13459 51598 13471 51632
rect 13505 51629 13517 51632
rect 30928 51629 30934 51641
rect 13505 51601 30934 51629
rect 13505 51598 13517 51601
rect 13459 51592 13517 51598
rect 30928 51589 30934 51601
rect 30986 51589 30992 51641
rect 4531 51558 4589 51564
rect 4531 51524 4543 51558
rect 4577 51555 4589 51558
rect 15859 51558 15917 51564
rect 4577 51527 7214 51555
rect 4577 51524 4589 51527
rect 4531 51518 4589 51524
rect 7186 51481 7214 51527
rect 15859 51524 15871 51558
rect 15905 51555 15917 51558
rect 16147 51558 16205 51564
rect 16147 51555 16159 51558
rect 15905 51527 16159 51555
rect 15905 51524 15917 51527
rect 15859 51518 15917 51524
rect 16147 51524 16159 51527
rect 16193 51555 16205 51558
rect 16243 51558 16301 51564
rect 16243 51555 16255 51558
rect 16193 51527 16255 51555
rect 16193 51524 16205 51527
rect 16147 51518 16205 51524
rect 16243 51524 16255 51527
rect 16289 51524 16301 51558
rect 23248 51555 23254 51567
rect 23209 51527 23254 51555
rect 16243 51518 16301 51524
rect 23248 51515 23254 51527
rect 23306 51555 23312 51567
rect 23443 51558 23501 51564
rect 23443 51555 23455 51558
rect 23306 51527 23455 51555
rect 23306 51515 23312 51527
rect 23443 51524 23455 51527
rect 23489 51524 23501 51558
rect 53392 51555 53398 51567
rect 23443 51518 23501 51524
rect 27346 51527 53398 51555
rect 27346 51481 27374 51527
rect 53392 51515 53398 51527
rect 53450 51515 53456 51567
rect 7186 51453 27374 51481
rect 16243 51410 16301 51416
rect 16243 51376 16255 51410
rect 16289 51407 16301 51410
rect 53200 51407 53206 51419
rect 16289 51379 53206 51407
rect 16289 51376 16301 51379
rect 16243 51370 16301 51376
rect 53200 51367 53206 51379
rect 53258 51367 53264 51419
rect 1152 51308 58848 51330
rect 1152 51256 19654 51308
rect 19706 51256 19718 51308
rect 19770 51256 19782 51308
rect 19834 51256 19846 51308
rect 19898 51256 50374 51308
rect 50426 51256 50438 51308
rect 50490 51256 50502 51308
rect 50554 51256 50566 51308
rect 50618 51256 58848 51308
rect 1152 51234 58848 51256
rect 20755 51188 20813 51194
rect 20755 51154 20767 51188
rect 20801 51185 20813 51188
rect 21424 51185 21430 51197
rect 20801 51157 21430 51185
rect 20801 51154 20813 51157
rect 20755 51148 20813 51154
rect 21424 51145 21430 51157
rect 21482 51145 21488 51197
rect 11040 50861 11102 50889
rect 11074 50827 11102 50861
rect 11266 50861 11328 50889
rect 11056 50775 11062 50827
rect 11114 50775 11120 50827
rect 10675 50744 10733 50750
rect 10675 50710 10687 50744
rect 10721 50741 10733 50744
rect 11155 50744 11213 50750
rect 11155 50741 11167 50744
rect 10721 50713 11167 50741
rect 10721 50710 10733 50713
rect 10675 50704 10733 50710
rect 11155 50710 11167 50713
rect 11201 50710 11213 50744
rect 11266 50741 11294 50861
rect 11539 50818 11597 50824
rect 11539 50815 11551 50818
rect 11424 50787 11551 50815
rect 11539 50784 11551 50787
rect 11585 50815 11597 50818
rect 14992 50815 14998 50827
rect 11585 50787 14998 50815
rect 11585 50784 11597 50787
rect 11539 50778 11597 50784
rect 14992 50775 14998 50787
rect 15050 50775 15056 50827
rect 14032 50741 14038 50753
rect 11266 50713 14038 50741
rect 11155 50704 11213 50710
rect 14032 50701 14038 50713
rect 14090 50701 14096 50753
rect 27187 50744 27245 50750
rect 27187 50710 27199 50744
rect 27233 50741 27245 50744
rect 27475 50744 27533 50750
rect 27475 50741 27487 50744
rect 27233 50713 27487 50741
rect 27233 50710 27245 50713
rect 27187 50704 27245 50710
rect 27475 50710 27487 50713
rect 27521 50741 27533 50744
rect 55024 50741 55030 50753
rect 27521 50713 55030 50741
rect 27521 50710 27533 50713
rect 27475 50704 27533 50710
rect 55024 50701 55030 50713
rect 55082 50701 55088 50753
rect 1152 50642 58848 50664
rect 1152 50590 4294 50642
rect 4346 50590 4358 50642
rect 4410 50590 4422 50642
rect 4474 50590 4486 50642
rect 4538 50590 35014 50642
rect 35066 50590 35078 50642
rect 35130 50590 35142 50642
rect 35194 50590 35206 50642
rect 35258 50590 58848 50642
rect 1152 50568 58848 50590
rect 47248 50405 47254 50457
rect 47306 50445 47312 50457
rect 47539 50448 47597 50454
rect 47539 50445 47551 50448
rect 47306 50417 47551 50445
rect 47306 50405 47312 50417
rect 47539 50414 47551 50417
rect 47585 50414 47597 50448
rect 47539 50408 47597 50414
rect 29971 50374 30029 50380
rect 29971 50340 29983 50374
rect 30017 50371 30029 50374
rect 34387 50374 34445 50380
rect 34387 50371 34399 50374
rect 30017 50343 34399 50371
rect 30017 50340 30029 50343
rect 29971 50334 30029 50340
rect 34387 50340 34399 50343
rect 34433 50340 34445 50374
rect 34387 50334 34445 50340
rect 25840 50257 25846 50309
rect 25898 50297 25904 50309
rect 55696 50297 55702 50309
rect 25898 50269 55702 50297
rect 25898 50257 25904 50269
rect 55696 50257 55702 50269
rect 55754 50257 55760 50309
rect 26323 50226 26381 50232
rect 26323 50192 26335 50226
rect 26369 50223 26381 50226
rect 26611 50226 26669 50232
rect 26611 50223 26623 50226
rect 26369 50195 26623 50223
rect 26369 50192 26381 50195
rect 26323 50186 26381 50192
rect 26611 50192 26623 50195
rect 26657 50223 26669 50226
rect 52432 50223 52438 50235
rect 26657 50195 52438 50223
rect 26657 50192 26669 50195
rect 26611 50186 26669 50192
rect 52432 50183 52438 50195
rect 52490 50183 52496 50235
rect 54451 50226 54509 50232
rect 54451 50192 54463 50226
rect 54497 50192 54509 50226
rect 54451 50186 54509 50192
rect 5584 50109 5590 50161
rect 5642 50149 5648 50161
rect 23347 50152 23405 50158
rect 23347 50149 23359 50152
rect 5642 50121 23359 50149
rect 5642 50109 5648 50121
rect 23347 50118 23359 50121
rect 23393 50118 23405 50152
rect 27760 50149 27766 50161
rect 23347 50112 23405 50118
rect 23458 50121 27766 50149
rect 6931 50078 6989 50084
rect 6931 50044 6943 50078
rect 6977 50075 6989 50078
rect 23458 50075 23486 50121
rect 27760 50109 27766 50121
rect 27818 50109 27824 50161
rect 29299 50152 29357 50158
rect 29299 50118 29311 50152
rect 29345 50149 29357 50152
rect 34387 50152 34445 50158
rect 29345 50121 34334 50149
rect 29345 50118 29357 50121
rect 29299 50112 29357 50118
rect 6977 50047 23486 50075
rect 34306 50075 34334 50121
rect 34387 50118 34399 50152
rect 34433 50149 34445 50152
rect 38800 50149 38806 50161
rect 34433 50121 38806 50149
rect 34433 50118 34445 50121
rect 34387 50112 34445 50118
rect 38800 50109 38806 50121
rect 38858 50109 38864 50161
rect 54466 50087 54494 50186
rect 46192 50075 46198 50087
rect 34306 50047 46198 50075
rect 6977 50044 6989 50047
rect 6931 50038 6989 50044
rect 46192 50035 46198 50047
rect 46250 50035 46256 50087
rect 47248 50035 47254 50087
rect 47306 50075 47312 50087
rect 47347 50078 47405 50084
rect 47347 50075 47359 50078
rect 47306 50047 47359 50075
rect 47306 50035 47312 50047
rect 47347 50044 47359 50047
rect 47393 50044 47405 50078
rect 47347 50038 47405 50044
rect 54355 50078 54413 50084
rect 54355 50044 54367 50078
rect 54401 50075 54413 50078
rect 54448 50075 54454 50087
rect 54401 50047 54454 50075
rect 54401 50044 54413 50047
rect 54355 50038 54413 50044
rect 54448 50035 54454 50047
rect 54506 50035 54512 50087
rect 1152 49976 58848 49998
rect 1152 49924 19654 49976
rect 19706 49924 19718 49976
rect 19770 49924 19782 49976
rect 19834 49924 19846 49976
rect 19898 49924 50374 49976
rect 50426 49924 50438 49976
rect 50490 49924 50502 49976
rect 50554 49924 50566 49976
rect 50618 49924 58848 49976
rect 1152 49902 58848 49924
rect 25558 49865 25610 49871
rect 25558 49807 25610 49813
rect 25840 49779 25846 49791
rect 25728 49751 25846 49779
rect 25840 49739 25846 49751
rect 25898 49739 25904 49791
rect 26016 49751 27374 49779
rect 27346 49705 27374 49751
rect 56944 49705 56950 49717
rect 27346 49677 56950 49705
rect 56944 49665 56950 49677
rect 57002 49665 57008 49717
rect 26707 49560 26765 49566
rect 26707 49526 26719 49560
rect 26753 49557 26765 49560
rect 46768 49557 46774 49569
rect 26753 49529 46774 49557
rect 26753 49526 26765 49529
rect 26707 49520 26765 49526
rect 46768 49517 46774 49529
rect 46826 49517 46832 49569
rect 22960 49443 22966 49495
rect 23018 49483 23024 49495
rect 23018 49455 23486 49483
rect 23018 49443 23024 49455
rect 12208 49409 12214 49421
rect 12169 49381 12214 49409
rect 12208 49369 12214 49381
rect 12266 49409 12272 49421
rect 12403 49412 12461 49418
rect 12403 49409 12415 49412
rect 12266 49381 12415 49409
rect 12266 49369 12272 49381
rect 12403 49378 12415 49381
rect 12449 49378 12461 49412
rect 23056 49409 23062 49421
rect 23017 49381 23062 49409
rect 12403 49372 12461 49378
rect 23056 49369 23062 49381
rect 23114 49409 23120 49421
rect 23155 49412 23213 49418
rect 23155 49409 23167 49412
rect 23114 49381 23167 49409
rect 23114 49369 23120 49381
rect 23155 49378 23167 49381
rect 23201 49378 23213 49412
rect 23458 49409 23486 49455
rect 31891 49412 31949 49418
rect 31891 49409 31903 49412
rect 23458 49381 31903 49409
rect 23155 49372 23213 49378
rect 31891 49378 31903 49381
rect 31937 49409 31949 49412
rect 32083 49412 32141 49418
rect 32083 49409 32095 49412
rect 31937 49381 32095 49409
rect 31937 49378 31949 49381
rect 31891 49372 31949 49378
rect 32083 49378 32095 49381
rect 32129 49378 32141 49412
rect 32083 49372 32141 49378
rect 1152 49310 58848 49332
rect 1152 49258 4294 49310
rect 4346 49258 4358 49310
rect 4410 49258 4422 49310
rect 4474 49258 4486 49310
rect 4538 49258 35014 49310
rect 35066 49258 35078 49310
rect 35130 49258 35142 49310
rect 35194 49258 35206 49310
rect 35258 49258 58848 49310
rect 1152 49236 58848 49258
rect 23155 49190 23213 49196
rect 23155 49156 23167 49190
rect 23201 49187 23213 49190
rect 26128 49187 26134 49199
rect 23201 49159 26134 49187
rect 23201 49156 23213 49159
rect 23155 49150 23213 49156
rect 26128 49147 26134 49159
rect 26186 49147 26192 49199
rect 55795 49190 55853 49196
rect 55795 49156 55807 49190
rect 55841 49187 55853 49190
rect 55888 49187 55894 49199
rect 55841 49159 55894 49187
rect 55841 49156 55853 49159
rect 55795 49150 55853 49156
rect 55888 49147 55894 49159
rect 55946 49147 55952 49199
rect 54355 48968 54413 48974
rect 54355 48934 54367 48968
rect 54401 48965 54413 48968
rect 54643 48968 54701 48974
rect 54643 48965 54655 48968
rect 54401 48937 54655 48965
rect 54401 48934 54413 48937
rect 54355 48928 54413 48934
rect 54643 48934 54655 48937
rect 54689 48965 54701 48968
rect 56272 48965 56278 48977
rect 54689 48937 56278 48965
rect 54689 48934 54701 48937
rect 54643 48928 54701 48934
rect 56272 48925 56278 48937
rect 56330 48925 56336 48977
rect 6931 48894 6989 48900
rect 6931 48860 6943 48894
rect 6977 48860 6989 48894
rect 6931 48854 6989 48860
rect 6946 48755 6974 48854
rect 6835 48746 6893 48752
rect 6835 48712 6847 48746
rect 6881 48743 6893 48746
rect 6928 48743 6934 48755
rect 6881 48715 6934 48743
rect 6881 48712 6893 48715
rect 6835 48706 6893 48712
rect 6928 48703 6934 48715
rect 6986 48703 6992 48755
rect 12691 48746 12749 48752
rect 12691 48712 12703 48746
rect 12737 48743 12749 48746
rect 46288 48743 46294 48755
rect 12737 48715 46294 48743
rect 12737 48712 12749 48715
rect 12691 48706 12749 48712
rect 46288 48703 46294 48715
rect 46346 48703 46352 48755
rect 1152 48644 58848 48666
rect 1152 48592 19654 48644
rect 19706 48592 19718 48644
rect 19770 48592 19782 48644
rect 19834 48592 19846 48644
rect 19898 48592 50374 48644
rect 50426 48592 50438 48644
rect 50490 48592 50502 48644
rect 50554 48592 50566 48644
rect 50618 48592 58848 48644
rect 1152 48570 58848 48592
rect 5392 48481 5398 48533
rect 5450 48521 5456 48533
rect 22864 48521 22870 48533
rect 5450 48493 6240 48521
rect 22368 48493 22870 48521
rect 5450 48481 5456 48493
rect 22864 48481 22870 48493
rect 22922 48481 22928 48533
rect 4816 48407 4822 48459
rect 4874 48447 4880 48459
rect 6064 48447 6070 48459
rect 4874 48419 5568 48447
rect 5856 48419 6070 48447
rect 4874 48407 4880 48419
rect 6064 48407 6070 48419
rect 6122 48407 6128 48459
rect 21952 48407 21958 48459
rect 22010 48407 22016 48459
rect 1152 47978 58848 48000
rect 1152 47926 4294 47978
rect 4346 47926 4358 47978
rect 4410 47926 4422 47978
rect 4474 47926 4486 47978
rect 4538 47926 35014 47978
rect 35066 47926 35078 47978
rect 35130 47926 35142 47978
rect 35194 47926 35206 47978
rect 35258 47926 58848 47978
rect 1152 47904 58848 47926
rect 27952 47519 27958 47571
rect 28010 47559 28016 47571
rect 31987 47562 32045 47568
rect 31987 47559 31999 47562
rect 28010 47531 31999 47559
rect 28010 47519 28016 47531
rect 31987 47528 31999 47531
rect 32033 47559 32045 47562
rect 32179 47562 32237 47568
rect 32179 47559 32191 47562
rect 32033 47531 32191 47559
rect 32033 47528 32045 47531
rect 31987 47522 32045 47528
rect 32179 47528 32191 47531
rect 32225 47528 32237 47562
rect 32179 47522 32237 47528
rect 1152 47312 58848 47334
rect 1152 47260 19654 47312
rect 19706 47260 19718 47312
rect 19770 47260 19782 47312
rect 19834 47260 19846 47312
rect 19898 47260 50374 47312
rect 50426 47260 50438 47312
rect 50490 47260 50502 47312
rect 50554 47260 50566 47312
rect 50618 47260 58848 47312
rect 1152 47238 58848 47260
rect 51568 46705 51574 46757
rect 51626 46745 51632 46757
rect 51667 46748 51725 46754
rect 51667 46745 51679 46748
rect 51626 46717 51679 46745
rect 51626 46705 51632 46717
rect 51667 46714 51679 46717
rect 51713 46745 51725 46748
rect 51859 46748 51917 46754
rect 51859 46745 51871 46748
rect 51713 46717 51871 46745
rect 51713 46714 51725 46717
rect 51667 46708 51725 46714
rect 51859 46714 51871 46717
rect 51905 46714 51917 46748
rect 51859 46708 51917 46714
rect 1152 46646 58848 46668
rect 1152 46594 4294 46646
rect 4346 46594 4358 46646
rect 4410 46594 4422 46646
rect 4474 46594 4486 46646
rect 4538 46594 35014 46646
rect 35066 46594 35078 46646
rect 35130 46594 35142 46646
rect 35194 46594 35206 46646
rect 35258 46594 58848 46646
rect 1152 46572 58848 46594
rect 29008 46335 29014 46387
rect 29066 46375 29072 46387
rect 35824 46375 35830 46387
rect 29066 46347 35830 46375
rect 29066 46335 29072 46347
rect 35824 46335 35830 46347
rect 35882 46335 35888 46387
rect 20464 46261 20470 46313
rect 20522 46301 20528 46313
rect 50899 46304 50957 46310
rect 50899 46301 50911 46304
rect 20522 46273 50911 46301
rect 20522 46261 20528 46273
rect 50899 46270 50911 46273
rect 50945 46270 50957 46304
rect 50899 46264 50957 46270
rect 12883 46230 12941 46236
rect 12883 46196 12895 46230
rect 12929 46196 12941 46230
rect 12883 46190 12941 46196
rect 13939 46230 13997 46236
rect 13939 46196 13951 46230
rect 13985 46196 13997 46230
rect 13939 46190 13997 46196
rect 23443 46230 23501 46236
rect 23443 46196 23455 46230
rect 23489 46196 23501 46230
rect 23443 46190 23501 46196
rect 26035 46230 26093 46236
rect 26035 46196 26047 46230
rect 26081 46227 26093 46230
rect 26323 46230 26381 46236
rect 26323 46227 26335 46230
rect 26081 46199 26335 46227
rect 26081 46196 26093 46199
rect 26035 46190 26093 46196
rect 26323 46196 26335 46199
rect 26369 46227 26381 46230
rect 30832 46227 30838 46239
rect 26369 46199 30838 46227
rect 26369 46196 26381 46199
rect 26323 46190 26381 46196
rect 12595 46156 12653 46162
rect 12595 46122 12607 46156
rect 12641 46153 12653 46156
rect 12784 46153 12790 46165
rect 12641 46125 12790 46153
rect 12641 46122 12653 46125
rect 12595 46116 12653 46122
rect 12784 46113 12790 46125
rect 12842 46153 12848 46165
rect 12898 46153 12926 46190
rect 13744 46153 13750 46165
rect 12842 46125 12926 46153
rect 13705 46125 13750 46153
rect 12842 46113 12848 46125
rect 13744 46113 13750 46125
rect 13802 46153 13808 46165
rect 13954 46153 13982 46190
rect 13802 46125 13982 46153
rect 23155 46156 23213 46162
rect 13802 46113 13808 46125
rect 23155 46122 23167 46156
rect 23201 46153 23213 46156
rect 23458 46153 23486 46190
rect 30832 46187 30838 46199
rect 30890 46187 30896 46239
rect 41008 46153 41014 46165
rect 23201 46125 41014 46153
rect 23201 46122 23213 46125
rect 23155 46116 23213 46122
rect 41008 46113 41014 46125
rect 41066 46113 41072 46165
rect 24400 46039 24406 46091
rect 24458 46079 24464 46091
rect 35635 46082 35693 46088
rect 35635 46079 35647 46082
rect 24458 46051 35647 46079
rect 24458 46039 24464 46051
rect 35635 46048 35647 46051
rect 35681 46048 35693 46082
rect 50032 46079 50038 46091
rect 49993 46051 50038 46079
rect 35635 46042 35693 46048
rect 50032 46039 50038 46051
rect 50090 46039 50096 46091
rect 1152 45980 58848 46002
rect 1152 45928 19654 45980
rect 19706 45928 19718 45980
rect 19770 45928 19782 45980
rect 19834 45928 19846 45980
rect 19898 45928 50374 45980
rect 50426 45928 50438 45980
rect 50490 45928 50502 45980
rect 50554 45928 50566 45980
rect 50618 45928 58848 45980
rect 1152 45906 58848 45928
rect 48304 45669 48310 45721
rect 48362 45709 48368 45721
rect 49075 45712 49133 45718
rect 49075 45709 49087 45712
rect 48362 45681 49087 45709
rect 48362 45669 48368 45681
rect 49075 45678 49087 45681
rect 49121 45678 49133 45712
rect 49075 45672 49133 45678
rect 27955 45416 28013 45422
rect 27955 45382 27967 45416
rect 28001 45413 28013 45416
rect 28240 45413 28246 45425
rect 28001 45385 28246 45413
rect 28001 45382 28013 45385
rect 27955 45376 28013 45382
rect 28240 45373 28246 45385
rect 28298 45373 28304 45425
rect 38896 45413 38902 45425
rect 38857 45385 38902 45413
rect 38896 45373 38902 45385
rect 38954 45413 38960 45425
rect 39091 45416 39149 45422
rect 39091 45413 39103 45416
rect 38954 45385 39103 45413
rect 38954 45373 38960 45385
rect 39091 45382 39103 45385
rect 39137 45382 39149 45416
rect 39091 45376 39149 45382
rect 1152 45314 58848 45336
rect 1152 45262 4294 45314
rect 4346 45262 4358 45314
rect 4410 45262 4422 45314
rect 4474 45262 4486 45314
rect 4538 45262 35014 45314
rect 35066 45262 35078 45314
rect 35130 45262 35142 45314
rect 35194 45262 35206 45314
rect 35258 45262 58848 45314
rect 1152 45240 58848 45262
rect 30160 45151 30166 45203
rect 30218 45191 30224 45203
rect 38896 45191 38902 45203
rect 30218 45163 38902 45191
rect 30218 45151 30224 45163
rect 38896 45151 38902 45163
rect 38954 45151 38960 45203
rect 28240 45077 28246 45129
rect 28298 45117 28304 45129
rect 48976 45117 48982 45129
rect 28298 45089 48982 45117
rect 28298 45077 28304 45089
rect 48976 45077 48982 45089
rect 49034 45077 49040 45129
rect 26323 44898 26381 44904
rect 26323 44864 26335 44898
rect 26369 44895 26381 44898
rect 26611 44898 26669 44904
rect 26611 44895 26623 44898
rect 26369 44867 26623 44895
rect 26369 44864 26381 44867
rect 26323 44858 26381 44864
rect 26611 44864 26623 44867
rect 26657 44895 26669 44898
rect 26657 44867 27374 44895
rect 26657 44864 26669 44867
rect 26611 44858 26669 44864
rect 27346 44747 27374 44867
rect 44464 44747 44470 44759
rect 27346 44719 44470 44747
rect 44464 44707 44470 44719
rect 44522 44707 44528 44759
rect 1152 44648 58848 44670
rect 1152 44596 19654 44648
rect 19706 44596 19718 44648
rect 19770 44596 19782 44648
rect 19834 44596 19846 44648
rect 19898 44596 50374 44648
rect 50426 44596 50438 44648
rect 50490 44596 50502 44648
rect 50554 44596 50566 44648
rect 50618 44596 58848 44648
rect 1152 44574 58848 44596
rect 7186 44127 37454 44155
rect 6352 44041 6358 44093
rect 6410 44081 6416 44093
rect 7186 44081 7214 44127
rect 6410 44053 7214 44081
rect 27091 44084 27149 44090
rect 6410 44041 6416 44053
rect 27091 44050 27103 44084
rect 27137 44081 27149 44084
rect 27379 44084 27437 44090
rect 27379 44081 27391 44084
rect 27137 44053 27391 44081
rect 27137 44050 27149 44053
rect 27091 44044 27149 44050
rect 27379 44050 27391 44053
rect 27425 44081 27437 44084
rect 30736 44081 30742 44093
rect 27425 44053 30742 44081
rect 27425 44050 27437 44053
rect 27379 44044 27437 44050
rect 30736 44041 30742 44053
rect 30794 44041 30800 44093
rect 32467 44084 32525 44090
rect 32467 44050 32479 44084
rect 32513 44081 32525 44084
rect 32752 44081 32758 44093
rect 32513 44053 32758 44081
rect 32513 44050 32525 44053
rect 32467 44044 32525 44050
rect 32752 44041 32758 44053
rect 32810 44041 32816 44093
rect 33136 44081 33142 44093
rect 33097 44053 33142 44081
rect 33136 44041 33142 44053
rect 33194 44081 33200 44093
rect 33331 44084 33389 44090
rect 33331 44081 33343 44084
rect 33194 44053 33343 44081
rect 33194 44041 33200 44053
rect 33331 44050 33343 44053
rect 33377 44050 33389 44084
rect 34768 44081 34774 44093
rect 34729 44053 34774 44081
rect 33331 44044 33389 44050
rect 34768 44041 34774 44053
rect 34826 44081 34832 44093
rect 34867 44084 34925 44090
rect 34867 44081 34879 44084
rect 34826 44053 34879 44081
rect 34826 44041 34832 44053
rect 34867 44050 34879 44053
rect 34913 44050 34925 44084
rect 37426 44081 37454 44127
rect 45619 44084 45677 44090
rect 45619 44081 45631 44084
rect 37426 44053 45631 44081
rect 34867 44044 34925 44050
rect 45619 44050 45631 44053
rect 45665 44050 45677 44084
rect 45619 44044 45677 44050
rect 55027 44084 55085 44090
rect 55027 44050 55039 44084
rect 55073 44081 55085 44084
rect 55312 44081 55318 44093
rect 55073 44053 55318 44081
rect 55073 44050 55085 44053
rect 55027 44044 55085 44050
rect 55312 44041 55318 44053
rect 55370 44041 55376 44093
rect 1152 43982 58848 44004
rect 1152 43930 4294 43982
rect 4346 43930 4358 43982
rect 4410 43930 4422 43982
rect 4474 43930 4486 43982
rect 4538 43930 35014 43982
rect 35066 43930 35078 43982
rect 35130 43930 35142 43982
rect 35194 43930 35206 43982
rect 35258 43930 58848 43982
rect 1152 43908 58848 43930
rect 30736 43819 30742 43871
rect 30794 43859 30800 43871
rect 55888 43859 55894 43871
rect 30794 43831 55894 43859
rect 30794 43819 30800 43831
rect 55888 43819 55894 43831
rect 55946 43819 55952 43871
rect 7600 43745 7606 43797
rect 7658 43785 7664 43797
rect 33136 43785 33142 43797
rect 7658 43757 33142 43785
rect 7658 43745 7664 43757
rect 33136 43745 33142 43757
rect 33194 43745 33200 43797
rect 32752 43671 32758 43723
rect 32810 43711 32816 43723
rect 49744 43711 49750 43723
rect 32810 43683 49750 43711
rect 32810 43671 32816 43683
rect 49744 43671 49750 43683
rect 49802 43671 49808 43723
rect 28243 43566 28301 43572
rect 28243 43563 28255 43566
rect 27346 43535 28255 43563
rect 26704 43375 26710 43427
rect 26762 43415 26768 43427
rect 27346 43415 27374 43535
rect 28243 43532 28255 43535
rect 28289 43563 28301 43566
rect 28339 43566 28397 43572
rect 28339 43563 28351 43566
rect 28289 43535 28351 43563
rect 28289 43532 28301 43535
rect 28243 43526 28301 43532
rect 28339 43532 28351 43535
rect 28385 43532 28397 43566
rect 28339 43526 28397 43532
rect 45907 43566 45965 43572
rect 45907 43532 45919 43566
rect 45953 43563 45965 43566
rect 46195 43566 46253 43572
rect 46195 43563 46207 43566
rect 45953 43535 46207 43563
rect 45953 43532 45965 43535
rect 45907 43526 45965 43532
rect 46195 43532 46207 43535
rect 46241 43563 46253 43566
rect 57136 43563 57142 43575
rect 46241 43535 57142 43563
rect 46241 43532 46253 43535
rect 46195 43526 46253 43532
rect 57136 43523 57142 43535
rect 57194 43523 57200 43575
rect 26762 43387 27374 43415
rect 26762 43375 26768 43387
rect 1152 43316 58848 43338
rect 1152 43264 19654 43316
rect 19706 43264 19718 43316
rect 19770 43264 19782 43316
rect 19834 43264 19846 43316
rect 19898 43264 50374 43316
rect 50426 43264 50438 43316
rect 50490 43264 50502 43316
rect 50554 43264 50566 43316
rect 50618 43264 58848 43316
rect 1152 43242 58848 43264
rect 50515 43048 50573 43054
rect 50515 43014 50527 43048
rect 50561 43045 50573 43048
rect 57808 43045 57814 43057
rect 50561 43017 57814 43045
rect 50561 43014 50573 43017
rect 50515 43008 50573 43014
rect 57808 43005 57814 43017
rect 57866 43005 57872 43057
rect 38128 42823 38134 42835
rect 27346 42795 38134 42823
rect 14803 42752 14861 42758
rect 14803 42718 14815 42752
rect 14849 42749 14861 42752
rect 15091 42752 15149 42758
rect 15091 42749 15103 42752
rect 14849 42721 15103 42749
rect 14849 42718 14861 42721
rect 14803 42712 14861 42718
rect 15091 42718 15103 42721
rect 15137 42749 15149 42752
rect 27346 42749 27374 42795
rect 38128 42783 38134 42795
rect 38186 42783 38192 42835
rect 34672 42749 34678 42761
rect 15137 42721 27374 42749
rect 34633 42721 34678 42749
rect 15137 42718 15149 42721
rect 15091 42712 15149 42718
rect 34672 42709 34678 42721
rect 34730 42749 34736 42761
rect 34867 42752 34925 42758
rect 34867 42749 34879 42752
rect 34730 42721 34879 42749
rect 34730 42709 34736 42721
rect 34867 42718 34879 42721
rect 34913 42718 34925 42752
rect 52528 42749 52534 42761
rect 52489 42721 52534 42749
rect 34867 42712 34925 42718
rect 52528 42709 52534 42721
rect 52586 42749 52592 42761
rect 52723 42752 52781 42758
rect 52723 42749 52735 42752
rect 52586 42721 52735 42749
rect 52586 42709 52592 42721
rect 52723 42718 52735 42721
rect 52769 42718 52781 42752
rect 52723 42712 52781 42718
rect 1152 42650 58848 42672
rect 1152 42598 4294 42650
rect 4346 42598 4358 42650
rect 4410 42598 4422 42650
rect 4474 42598 4486 42650
rect 4538 42598 35014 42650
rect 35066 42598 35078 42650
rect 35130 42598 35142 42650
rect 35194 42598 35206 42650
rect 35258 42598 58848 42650
rect 1152 42576 58848 42598
rect 17968 42487 17974 42539
rect 18026 42527 18032 42539
rect 34672 42527 34678 42539
rect 18026 42499 34678 42527
rect 18026 42487 18032 42499
rect 34672 42487 34678 42499
rect 34730 42487 34736 42539
rect 41104 42487 41110 42539
rect 41162 42527 41168 42539
rect 52528 42527 52534 42539
rect 41162 42499 52534 42527
rect 41162 42487 41168 42499
rect 52528 42487 52534 42499
rect 52586 42487 52592 42539
rect 30064 42191 30070 42243
rect 30122 42231 30128 42243
rect 30163 42234 30221 42240
rect 30163 42231 30175 42234
rect 30122 42203 30175 42231
rect 30122 42191 30128 42203
rect 30163 42200 30175 42203
rect 30209 42200 30221 42234
rect 30163 42194 30221 42200
rect 43696 42191 43702 42243
rect 43754 42231 43760 42243
rect 54931 42234 54989 42240
rect 54931 42231 54943 42234
rect 43754 42203 54943 42231
rect 43754 42191 43760 42203
rect 54931 42200 54943 42203
rect 54977 42231 54989 42234
rect 55123 42234 55181 42240
rect 55123 42231 55135 42234
rect 54977 42203 55135 42231
rect 54977 42200 54989 42203
rect 54931 42194 54989 42200
rect 55123 42200 55135 42203
rect 55169 42200 55181 42234
rect 55123 42194 55181 42200
rect 28051 42160 28109 42166
rect 28051 42126 28063 42160
rect 28097 42157 28109 42160
rect 28097 42129 37454 42157
rect 28097 42126 28109 42129
rect 28051 42120 28109 42126
rect 30064 42083 30070 42095
rect 30025 42055 30070 42083
rect 30064 42043 30070 42055
rect 30122 42043 30128 42095
rect 37426 42083 37454 42129
rect 40816 42083 40822 42095
rect 37426 42055 40822 42083
rect 40816 42043 40822 42055
rect 40874 42043 40880 42095
rect 1152 41984 58848 42006
rect 1152 41932 19654 41984
rect 19706 41932 19718 41984
rect 19770 41932 19782 41984
rect 19834 41932 19846 41984
rect 19898 41932 50374 41984
rect 50426 41932 50438 41984
rect 50490 41932 50502 41984
rect 50554 41932 50566 41984
rect 50618 41932 58848 41984
rect 1152 41910 58848 41932
rect 7312 41525 7318 41577
rect 7370 41565 7376 41577
rect 7370 41537 22176 41565
rect 22306 41537 22464 41565
rect 7370 41525 7376 41537
rect 9328 41451 9334 41503
rect 9386 41491 9392 41503
rect 22195 41494 22253 41500
rect 22195 41491 22207 41494
rect 9386 41463 22207 41491
rect 9386 41451 9392 41463
rect 22195 41460 22207 41463
rect 22241 41460 22253 41494
rect 22195 41454 22253 41460
rect 5200 41377 5206 41429
rect 5258 41417 5264 41429
rect 22306 41417 22334 41537
rect 5258 41389 22334 41417
rect 22387 41420 22445 41426
rect 5258 41377 5264 41389
rect 22387 41386 22399 41420
rect 22433 41417 22445 41420
rect 22834 41417 22862 41477
rect 22433 41389 22862 41417
rect 22433 41386 22445 41389
rect 22387 41380 22445 41386
rect 42064 41377 42070 41429
rect 42122 41417 42128 41429
rect 42259 41420 42317 41426
rect 42259 41417 42271 41420
rect 42122 41389 42271 41417
rect 42122 41377 42128 41389
rect 42259 41386 42271 41389
rect 42305 41417 42317 41420
rect 42451 41420 42509 41426
rect 42451 41417 42463 41420
rect 42305 41389 42463 41417
rect 42305 41386 42317 41389
rect 42259 41380 42317 41386
rect 42451 41386 42463 41389
rect 42497 41386 42509 41420
rect 42451 41380 42509 41386
rect 57139 41420 57197 41426
rect 57139 41386 57151 41420
rect 57185 41417 57197 41420
rect 57232 41417 57238 41429
rect 57185 41389 57238 41417
rect 57185 41386 57197 41389
rect 57139 41380 57197 41386
rect 57232 41377 57238 41389
rect 57290 41377 57296 41429
rect 1152 41318 58848 41340
rect 1152 41266 4294 41318
rect 4346 41266 4358 41318
rect 4410 41266 4422 41318
rect 4474 41266 4486 41318
rect 4538 41266 35014 41318
rect 35066 41266 35078 41318
rect 35130 41266 35142 41318
rect 35194 41266 35206 41318
rect 35258 41266 58848 41318
rect 1152 41244 58848 41266
rect 8560 40933 8566 40985
rect 8618 40973 8624 40985
rect 45715 40976 45773 40982
rect 45715 40973 45727 40976
rect 8618 40945 45727 40973
rect 8618 40933 8624 40945
rect 45715 40942 45727 40945
rect 45761 40942 45773 40976
rect 45715 40936 45773 40942
rect 23347 40902 23405 40908
rect 23347 40868 23359 40902
rect 23393 40868 23405 40902
rect 23347 40862 23405 40868
rect 23059 40828 23117 40834
rect 23059 40794 23071 40828
rect 23105 40825 23117 40828
rect 23362 40825 23390 40862
rect 26800 40859 26806 40911
rect 26858 40899 26864 40911
rect 30163 40902 30221 40908
rect 30163 40899 30175 40902
rect 26858 40871 30175 40899
rect 26858 40859 26864 40871
rect 30163 40868 30175 40871
rect 30209 40868 30221 40902
rect 30163 40862 30221 40868
rect 23105 40797 27374 40825
rect 23105 40794 23117 40797
rect 23059 40788 23117 40794
rect 27346 40751 27374 40797
rect 41200 40751 41206 40763
rect 27346 40723 41206 40751
rect 41200 40711 41206 40723
rect 41258 40711 41264 40763
rect 1152 40652 58848 40674
rect 1152 40600 19654 40652
rect 19706 40600 19718 40652
rect 19770 40600 19782 40652
rect 19834 40600 19846 40652
rect 19898 40600 50374 40652
rect 50426 40600 50438 40652
rect 50490 40600 50502 40652
rect 50554 40600 50566 40652
rect 50618 40600 58848 40652
rect 1152 40578 58848 40600
rect 7216 40341 7222 40393
rect 7274 40381 7280 40393
rect 49555 40384 49613 40390
rect 49555 40381 49567 40384
rect 7274 40353 49567 40381
rect 7274 40341 7280 40353
rect 49555 40350 49567 40353
rect 49601 40350 49613 40384
rect 49555 40344 49613 40350
rect 16723 40310 16781 40316
rect 16723 40276 16735 40310
rect 16769 40307 16781 40310
rect 18064 40307 18070 40319
rect 16769 40279 18070 40307
rect 16769 40276 16781 40279
rect 16723 40270 16781 40276
rect 18064 40267 18070 40279
rect 18122 40267 18128 40319
rect 52048 40307 52054 40319
rect 52009 40279 52054 40307
rect 52048 40267 52054 40279
rect 52106 40267 52112 40319
rect 1152 39986 58848 40008
rect 1152 39934 4294 39986
rect 4346 39934 4358 39986
rect 4410 39934 4422 39986
rect 4474 39934 4486 39986
rect 4538 39934 35014 39986
rect 35066 39934 35078 39986
rect 35130 39934 35142 39986
rect 35194 39934 35206 39986
rect 35258 39934 58848 39986
rect 1152 39912 58848 39934
rect 12115 39570 12173 39576
rect 12115 39536 12127 39570
rect 12161 39567 12173 39570
rect 12403 39570 12461 39576
rect 12403 39567 12415 39570
rect 12161 39539 12415 39567
rect 12161 39536 12173 39539
rect 12115 39530 12173 39536
rect 12403 39536 12415 39539
rect 12449 39567 12461 39570
rect 12449 39539 17294 39567
rect 12449 39536 12461 39539
rect 12403 39530 12461 39536
rect 17266 39419 17294 39539
rect 25168 39527 25174 39579
rect 25226 39567 25232 39579
rect 46672 39567 46678 39579
rect 25226 39539 46678 39567
rect 25226 39527 25232 39539
rect 46672 39527 46678 39539
rect 46730 39527 46736 39579
rect 25264 39453 25270 39505
rect 25322 39493 25328 39505
rect 47536 39493 47542 39505
rect 25322 39465 47542 39493
rect 25322 39453 25328 39465
rect 47536 39453 47542 39465
rect 47594 39453 47600 39505
rect 45328 39419 45334 39431
rect 17266 39391 45334 39419
rect 45328 39379 45334 39391
rect 45386 39379 45392 39431
rect 1152 39320 58848 39342
rect 1152 39268 19654 39320
rect 19706 39268 19718 39320
rect 19770 39268 19782 39320
rect 19834 39268 19846 39320
rect 19898 39268 50374 39320
rect 50426 39268 50438 39320
rect 50490 39268 50502 39320
rect 50554 39268 50566 39320
rect 50618 39268 58848 39320
rect 1152 39246 58848 39268
rect 47536 39197 47542 39209
rect 47122 39169 47542 39197
rect 46816 39083 46822 39135
rect 46874 39083 46880 39135
rect 47122 39109 47150 39169
rect 47536 39157 47542 39169
rect 47594 39157 47600 39209
rect 47362 38873 47424 38901
rect 36208 38827 36214 38839
rect 7186 38799 36214 38827
rect 5875 38756 5933 38762
rect 5875 38722 5887 38756
rect 5921 38753 5933 38756
rect 7186 38753 7214 38799
rect 36208 38787 36214 38799
rect 36266 38787 36272 38839
rect 5921 38725 7214 38753
rect 21235 38756 21293 38762
rect 5921 38722 5933 38725
rect 5875 38716 5933 38722
rect 21235 38722 21247 38756
rect 21281 38753 21293 38756
rect 21328 38753 21334 38765
rect 21281 38725 21334 38753
rect 21281 38722 21293 38725
rect 21235 38716 21293 38722
rect 21328 38713 21334 38725
rect 21386 38713 21392 38765
rect 26899 38756 26957 38762
rect 26899 38722 26911 38756
rect 26945 38753 26957 38756
rect 27184 38753 27190 38765
rect 26945 38725 27190 38753
rect 26945 38722 26957 38725
rect 26899 38716 26957 38722
rect 27184 38713 27190 38725
rect 27242 38713 27248 38765
rect 41296 38713 41302 38765
rect 41354 38753 41360 38765
rect 46387 38756 46445 38762
rect 46387 38753 46399 38756
rect 41354 38725 46399 38753
rect 41354 38713 41360 38725
rect 46387 38722 46399 38725
rect 46433 38753 46445 38756
rect 46690 38753 46718 38813
rect 46433 38725 46718 38753
rect 46433 38722 46445 38725
rect 46387 38716 46445 38722
rect 46864 38713 46870 38765
rect 46922 38753 46928 38765
rect 47362 38753 47390 38873
rect 46922 38725 47390 38753
rect 46922 38713 46928 38725
rect 1152 38654 58848 38676
rect 1152 38602 4294 38654
rect 4346 38602 4358 38654
rect 4410 38602 4422 38654
rect 4474 38602 4486 38654
rect 4538 38602 35014 38654
rect 35066 38602 35078 38654
rect 35130 38602 35142 38654
rect 35194 38602 35206 38654
rect 35258 38602 58848 38654
rect 1152 38580 58848 38602
rect 27184 38491 27190 38543
rect 27242 38531 27248 38543
rect 39184 38531 39190 38543
rect 27242 38503 39190 38531
rect 27242 38491 27248 38503
rect 39184 38491 39190 38503
rect 39242 38491 39248 38543
rect 13552 38343 13558 38395
rect 13610 38383 13616 38395
rect 15955 38386 16013 38392
rect 15955 38383 15967 38386
rect 13610 38355 15967 38383
rect 13610 38343 13616 38355
rect 15955 38352 15967 38355
rect 16001 38352 16013 38386
rect 15955 38346 16013 38352
rect 27346 38281 30686 38309
rect 24688 38195 24694 38247
rect 24746 38235 24752 38247
rect 27346 38235 27374 38281
rect 30256 38235 30262 38247
rect 24746 38207 27374 38235
rect 30169 38207 30262 38235
rect 24746 38195 24752 38207
rect 30256 38195 30262 38207
rect 30314 38235 30320 38247
rect 30547 38238 30605 38244
rect 30547 38235 30559 38238
rect 30314 38207 30559 38235
rect 30314 38195 30320 38207
rect 30547 38204 30559 38207
rect 30593 38204 30605 38238
rect 30658 38235 30686 38281
rect 32464 38269 32470 38321
rect 32522 38309 32528 38321
rect 52051 38312 52109 38318
rect 52051 38309 52063 38312
rect 32522 38281 52063 38309
rect 32522 38269 32528 38281
rect 52051 38278 52063 38281
rect 52097 38278 52109 38312
rect 52051 38272 52109 38278
rect 57715 38238 57773 38244
rect 57715 38235 57727 38238
rect 30658 38207 43214 38235
rect 30547 38198 30605 38204
rect 15184 38121 15190 38173
rect 15242 38161 15248 38173
rect 32368 38161 32374 38173
rect 15242 38133 32374 38161
rect 15242 38121 15248 38133
rect 32368 38121 32374 38133
rect 32426 38121 32432 38173
rect 43186 38161 43214 38207
rect 57586 38207 57727 38235
rect 57586 38161 57614 38207
rect 57715 38204 57727 38207
rect 57761 38235 57773 38238
rect 57811 38238 57869 38244
rect 57811 38235 57823 38238
rect 57761 38207 57823 38235
rect 57761 38204 57773 38207
rect 57715 38198 57773 38204
rect 57811 38204 57823 38207
rect 57857 38204 57869 38238
rect 57811 38198 57869 38204
rect 43186 38133 57614 38161
rect 1152 37988 58848 38010
rect 1152 37936 19654 37988
rect 19706 37936 19718 37988
rect 19770 37936 19782 37988
rect 19834 37936 19846 37988
rect 19898 37936 50374 37988
rect 50426 37936 50438 37988
rect 50490 37936 50502 37988
rect 50554 37936 50566 37988
rect 50618 37936 58848 37988
rect 1152 37914 58848 37936
rect 41491 37498 41549 37504
rect 41491 37464 41503 37498
rect 41537 37495 41549 37498
rect 41537 37467 41822 37495
rect 41537 37464 41549 37467
rect 41491 37458 41549 37464
rect 41794 37433 41822 37467
rect 42928 37455 42934 37507
rect 42986 37495 42992 37507
rect 43027 37498 43085 37504
rect 43027 37495 43039 37498
rect 42986 37467 43039 37495
rect 42986 37455 42992 37467
rect 43027 37464 43039 37467
rect 43073 37464 43085 37498
rect 43027 37458 43085 37464
rect 16339 37424 16397 37430
rect 16339 37390 16351 37424
rect 16385 37421 16397 37424
rect 16432 37421 16438 37433
rect 16385 37393 16438 37421
rect 16385 37390 16397 37393
rect 16339 37384 16397 37390
rect 16432 37381 16438 37393
rect 16490 37381 16496 37433
rect 41776 37421 41782 37433
rect 41689 37393 41782 37421
rect 41776 37381 41782 37393
rect 41834 37381 41840 37433
rect 43042 37421 43070 37458
rect 43219 37424 43277 37430
rect 43219 37421 43231 37424
rect 43042 37393 43231 37421
rect 43219 37390 43231 37393
rect 43265 37390 43277 37424
rect 43219 37384 43277 37390
rect 53776 37381 53782 37433
rect 53834 37421 53840 37433
rect 53875 37424 53933 37430
rect 53875 37421 53887 37424
rect 53834 37393 53887 37421
rect 53834 37381 53840 37393
rect 53875 37390 53887 37393
rect 53921 37421 53933 37424
rect 54067 37424 54125 37430
rect 54067 37421 54079 37424
rect 53921 37393 54079 37421
rect 53921 37390 53933 37393
rect 53875 37384 53933 37390
rect 54067 37390 54079 37393
rect 54113 37390 54125 37424
rect 54067 37384 54125 37390
rect 1152 37322 58848 37344
rect 1152 37270 4294 37322
rect 4346 37270 4358 37322
rect 4410 37270 4422 37322
rect 4474 37270 4486 37322
rect 4538 37270 35014 37322
rect 35066 37270 35078 37322
rect 35130 37270 35142 37322
rect 35194 37270 35206 37322
rect 35258 37270 58848 37322
rect 1152 37248 58848 37270
rect 41776 37159 41782 37211
rect 41834 37199 41840 37211
rect 53104 37199 53110 37211
rect 41834 37171 53110 37199
rect 41834 37159 41840 37171
rect 53104 37159 53110 37171
rect 53162 37159 53168 37211
rect 32752 37085 32758 37137
rect 32810 37125 32816 37137
rect 53776 37125 53782 37137
rect 32810 37097 53782 37125
rect 32810 37085 32816 37097
rect 53776 37085 53782 37097
rect 53834 37085 53840 37137
rect 25360 36715 25366 36767
rect 25418 36755 25424 36767
rect 42928 36755 42934 36767
rect 25418 36727 42934 36755
rect 25418 36715 25424 36727
rect 42928 36715 42934 36727
rect 42986 36715 42992 36767
rect 1152 36656 58848 36678
rect 1152 36604 19654 36656
rect 19706 36604 19718 36656
rect 19770 36604 19782 36656
rect 19834 36604 19846 36656
rect 19898 36604 50374 36656
rect 50426 36604 50438 36656
rect 50490 36604 50502 36656
rect 50554 36604 50566 36656
rect 50618 36604 58848 36656
rect 1152 36582 58848 36604
rect 2707 36240 2765 36246
rect 2707 36206 2719 36240
rect 2753 36237 2765 36240
rect 20368 36237 20374 36249
rect 2753 36209 20374 36237
rect 2753 36206 2765 36209
rect 2707 36200 2765 36206
rect 20368 36197 20374 36209
rect 20426 36197 20432 36249
rect 1651 36092 1709 36098
rect 1651 36058 1663 36092
rect 1697 36089 1709 36092
rect 1936 36089 1942 36101
rect 1697 36061 1942 36089
rect 1697 36058 1709 36061
rect 1651 36052 1709 36058
rect 1936 36049 1942 36061
rect 1994 36049 2000 36101
rect 7984 36049 7990 36101
rect 8042 36089 8048 36101
rect 22387 36092 22445 36098
rect 22387 36089 22399 36092
rect 8042 36061 22399 36089
rect 8042 36049 8048 36061
rect 22387 36058 22399 36061
rect 22433 36089 22445 36092
rect 22579 36092 22637 36098
rect 22579 36089 22591 36092
rect 22433 36061 22591 36089
rect 22433 36058 22445 36061
rect 22387 36052 22445 36058
rect 22579 36058 22591 36061
rect 22625 36058 22637 36092
rect 38512 36089 38518 36101
rect 38473 36061 38518 36089
rect 22579 36052 22637 36058
rect 38512 36049 38518 36061
rect 38570 36049 38576 36101
rect 54736 36089 54742 36101
rect 54697 36061 54742 36089
rect 54736 36049 54742 36061
rect 54794 36089 54800 36101
rect 54835 36092 54893 36098
rect 54835 36089 54847 36092
rect 54794 36061 54847 36089
rect 54794 36049 54800 36061
rect 54835 36058 54847 36061
rect 54881 36058 54893 36092
rect 54835 36052 54893 36058
rect 1152 35990 58848 36012
rect 1152 35938 4294 35990
rect 4346 35938 4358 35990
rect 4410 35938 4422 35990
rect 4474 35938 4486 35990
rect 4538 35938 35014 35990
rect 35066 35938 35078 35990
rect 35130 35938 35142 35990
rect 35194 35938 35206 35990
rect 35258 35938 58848 35990
rect 1152 35916 58848 35938
rect 22672 35719 22678 35731
rect 7186 35691 22678 35719
rect 4528 35605 4534 35657
rect 4586 35645 4592 35657
rect 7186 35645 7214 35691
rect 22672 35679 22678 35691
rect 22730 35679 22736 35731
rect 4586 35617 7214 35645
rect 20290 35617 27374 35645
rect 4586 35605 4592 35617
rect 2323 35574 2381 35580
rect 2323 35540 2335 35574
rect 2369 35571 2381 35574
rect 2611 35574 2669 35580
rect 2611 35571 2623 35574
rect 2369 35543 2623 35571
rect 2369 35540 2381 35543
rect 2323 35534 2381 35540
rect 2611 35540 2623 35543
rect 2657 35571 2669 35574
rect 20290 35571 20318 35617
rect 20464 35571 20470 35583
rect 2657 35543 20318 35571
rect 20425 35543 20470 35571
rect 2657 35540 2669 35543
rect 2611 35534 2669 35540
rect 20464 35531 20470 35543
rect 20522 35531 20528 35583
rect 21331 35574 21389 35580
rect 21331 35540 21343 35574
rect 21377 35571 21389 35574
rect 21619 35574 21677 35580
rect 21619 35571 21631 35574
rect 21377 35543 21631 35571
rect 21377 35540 21389 35543
rect 21331 35534 21389 35540
rect 21619 35540 21631 35543
rect 21665 35540 21677 35574
rect 27346 35571 27374 35617
rect 39952 35571 39958 35583
rect 27346 35543 39958 35571
rect 21619 35534 21677 35540
rect 9427 35500 9485 35506
rect 9427 35466 9439 35500
rect 9473 35497 9485 35500
rect 21634 35497 21662 35534
rect 39952 35531 39958 35543
rect 40010 35531 40016 35583
rect 45043 35574 45101 35580
rect 45043 35540 45055 35574
rect 45089 35540 45101 35574
rect 49171 35574 49229 35580
rect 49171 35571 49183 35574
rect 45043 35534 45101 35540
rect 48994 35543 49183 35571
rect 35920 35497 35926 35509
rect 9473 35469 21374 35497
rect 21634 35469 35926 35497
rect 9473 35466 9485 35469
rect 9427 35460 9485 35466
rect 21346 35423 21374 35469
rect 35920 35457 35926 35469
rect 35978 35457 35984 35509
rect 32560 35423 32566 35435
rect 21346 35395 32566 35423
rect 32560 35383 32566 35395
rect 32618 35383 32624 35435
rect 44368 35383 44374 35435
rect 44426 35423 44432 35435
rect 44851 35426 44909 35432
rect 44851 35423 44863 35426
rect 44426 35395 44863 35423
rect 44426 35383 44432 35395
rect 44851 35392 44863 35395
rect 44897 35423 44909 35426
rect 45058 35423 45086 35534
rect 44897 35395 45086 35423
rect 44897 35392 44909 35395
rect 44851 35386 44909 35392
rect 47920 35383 47926 35435
rect 47978 35423 47984 35435
rect 48994 35432 49022 35543
rect 49171 35540 49183 35543
rect 49217 35540 49229 35574
rect 49171 35534 49229 35540
rect 51379 35574 51437 35580
rect 51379 35540 51391 35574
rect 51425 35540 51437 35574
rect 51379 35534 51437 35540
rect 48979 35426 49037 35432
rect 48979 35423 48991 35426
rect 47978 35395 48991 35423
rect 47978 35383 47984 35395
rect 48979 35392 48991 35395
rect 49025 35392 49037 35426
rect 51184 35423 51190 35435
rect 51145 35395 51190 35423
rect 48979 35386 49037 35392
rect 51184 35383 51190 35395
rect 51242 35423 51248 35435
rect 51394 35423 51422 35534
rect 51242 35395 51422 35423
rect 51242 35383 51248 35395
rect 1152 35324 58848 35346
rect 1152 35272 19654 35324
rect 19706 35272 19718 35324
rect 19770 35272 19782 35324
rect 19834 35272 19846 35324
rect 19898 35272 50374 35324
rect 50426 35272 50438 35324
rect 50490 35272 50502 35324
rect 50554 35272 50566 35324
rect 50618 35272 58848 35324
rect 1152 35250 58848 35272
rect 29392 35161 29398 35213
rect 29450 35201 29456 35213
rect 51184 35201 51190 35213
rect 29450 35173 51190 35201
rect 29450 35161 29456 35173
rect 51184 35161 51190 35173
rect 51242 35161 51248 35213
rect 21616 35087 21622 35139
rect 21674 35127 21680 35139
rect 21674 35099 21888 35127
rect 21674 35087 21680 35099
rect 4528 35053 4534 35065
rect 4489 35025 4534 35053
rect 4528 35013 4534 35025
rect 4586 35013 4592 35065
rect 19120 34865 19126 34917
rect 19178 34905 19184 34917
rect 21043 34908 21101 34914
rect 21043 34905 21055 34908
rect 19178 34877 21055 34905
rect 19178 34865 19184 34877
rect 21043 34874 21055 34877
rect 21089 34874 21101 34908
rect 21043 34868 21101 34874
rect 21331 34908 21389 34914
rect 21331 34874 21343 34908
rect 21377 34905 21389 34908
rect 21377 34877 21600 34905
rect 21377 34874 21389 34877
rect 21331 34868 21389 34874
rect 19984 34791 19990 34843
rect 20042 34831 20048 34843
rect 21043 34834 21101 34840
rect 21043 34831 21055 34834
rect 20042 34803 21055 34831
rect 20042 34791 20048 34803
rect 21043 34800 21055 34803
rect 21089 34800 21101 34834
rect 21331 34834 21389 34840
rect 21043 34794 21101 34800
rect 17776 34757 17782 34769
rect 17737 34729 17782 34757
rect 17776 34717 17782 34729
rect 17834 34717 17840 34769
rect 20368 34717 20374 34769
rect 20426 34757 20432 34769
rect 20851 34760 20909 34766
rect 20851 34757 20863 34760
rect 20426 34729 20863 34757
rect 20426 34717 20432 34729
rect 20851 34726 20863 34729
rect 20897 34757 20909 34760
rect 21202 34757 21230 34817
rect 21331 34800 21343 34834
rect 21377 34831 21389 34834
rect 21377 34803 27374 34831
rect 21377 34800 21389 34803
rect 21331 34794 21389 34800
rect 20897 34729 21230 34757
rect 27346 34757 27374 34803
rect 50035 34760 50093 34766
rect 50035 34757 50047 34760
rect 27346 34729 50047 34757
rect 20897 34726 20909 34729
rect 20851 34720 20909 34726
rect 50035 34726 50047 34729
rect 50081 34757 50093 34760
rect 50227 34760 50285 34766
rect 50227 34757 50239 34760
rect 50081 34729 50239 34757
rect 50081 34726 50093 34729
rect 50035 34720 50093 34726
rect 50227 34726 50239 34729
rect 50273 34726 50285 34760
rect 50227 34720 50285 34726
rect 1152 34658 58848 34680
rect 1152 34606 4294 34658
rect 4346 34606 4358 34658
rect 4410 34606 4422 34658
rect 4474 34606 4486 34658
rect 4538 34606 35014 34658
rect 35066 34606 35078 34658
rect 35130 34606 35142 34658
rect 35194 34606 35206 34658
rect 35258 34606 58848 34658
rect 1152 34584 58848 34606
rect 21331 34242 21389 34248
rect 21331 34208 21343 34242
rect 21377 34239 21389 34242
rect 33808 34239 33814 34251
rect 21377 34211 33814 34239
rect 21377 34208 21389 34211
rect 21331 34202 21389 34208
rect 33808 34199 33814 34211
rect 33866 34199 33872 34251
rect 36688 34239 36694 34251
rect 36649 34211 36694 34239
rect 36688 34199 36694 34211
rect 36746 34199 36752 34251
rect 17776 34051 17782 34103
rect 17834 34091 17840 34103
rect 32464 34091 32470 34103
rect 17834 34063 32470 34091
rect 17834 34051 17840 34063
rect 32464 34051 32470 34063
rect 32522 34051 32528 34103
rect 1152 33992 58848 34014
rect 1152 33940 19654 33992
rect 19706 33940 19718 33992
rect 19770 33940 19782 33992
rect 19834 33940 19846 33992
rect 19898 33940 50374 33992
rect 50426 33940 50438 33992
rect 50490 33940 50502 33992
rect 50554 33940 50566 33992
rect 50618 33940 58848 33992
rect 1152 33918 58848 33940
rect 9328 33829 9334 33881
rect 9386 33869 9392 33881
rect 57232 33869 57238 33881
rect 9386 33841 57238 33869
rect 9386 33829 9392 33841
rect 57232 33829 57238 33841
rect 57290 33829 57296 33881
rect 41392 33459 41398 33511
rect 41450 33499 41456 33511
rect 52531 33502 52589 33508
rect 52531 33499 52543 33502
rect 41450 33471 52543 33499
rect 41450 33459 41456 33471
rect 52531 33468 52543 33471
rect 52577 33499 52589 33502
rect 52723 33502 52781 33508
rect 52723 33499 52735 33502
rect 52577 33471 52735 33499
rect 52577 33468 52589 33471
rect 52531 33462 52589 33468
rect 52723 33468 52735 33471
rect 52769 33468 52781 33502
rect 52723 33462 52781 33468
rect 45619 33428 45677 33434
rect 45619 33394 45631 33428
rect 45665 33425 45677 33428
rect 45712 33425 45718 33437
rect 45665 33397 45718 33425
rect 45665 33394 45677 33397
rect 45619 33388 45677 33394
rect 45712 33385 45718 33397
rect 45770 33385 45776 33437
rect 1152 33326 58848 33348
rect 1152 33274 4294 33326
rect 4346 33274 4358 33326
rect 4410 33274 4422 33326
rect 4474 33274 4486 33326
rect 4538 33274 35014 33326
rect 35066 33274 35078 33326
rect 35130 33274 35142 33326
rect 35194 33274 35206 33326
rect 35258 33274 58848 33326
rect 1152 33252 58848 33274
rect 57331 33206 57389 33212
rect 57331 33172 57343 33206
rect 57377 33203 57389 33206
rect 57904 33203 57910 33215
rect 57377 33175 57910 33203
rect 57377 33172 57389 33175
rect 57331 33166 57389 33172
rect 57904 33163 57910 33175
rect 57962 33163 57968 33215
rect 10000 33129 10006 33141
rect 8434 33101 10006 33129
rect 8434 33041 8462 33101
rect 10000 33089 10006 33101
rect 10058 33089 10064 33141
rect 8851 33058 8909 33064
rect 8851 33055 8863 33058
rect 8736 33027 8863 33055
rect 8851 33024 8863 33027
rect 8897 33024 8909 33058
rect 8851 33018 8909 33024
rect 8992 33015 8998 33067
rect 9050 33015 9056 33067
rect 9139 33058 9197 33064
rect 9139 33024 9151 33058
rect 9185 33055 9197 33058
rect 13072 33055 13078 33067
rect 9185 33027 13078 33055
rect 9185 33024 9197 33027
rect 9139 33018 9197 33024
rect 13072 33015 13078 33027
rect 13130 33015 13136 33067
rect 8848 32719 8854 32771
rect 8906 32719 8912 32771
rect 1152 32660 58848 32682
rect 1152 32608 19654 32660
rect 19706 32608 19718 32660
rect 19770 32608 19782 32660
rect 19834 32608 19846 32660
rect 19898 32608 50374 32660
rect 50426 32608 50438 32660
rect 50490 32608 50502 32660
rect 50554 32608 50566 32660
rect 50618 32608 58848 32660
rect 1152 32586 58848 32608
rect 6832 32497 6838 32549
rect 6890 32497 6896 32549
rect 8848 32497 8854 32549
rect 8906 32537 8912 32549
rect 15280 32537 15286 32549
rect 8906 32509 15286 32537
rect 8906 32497 8912 32509
rect 15280 32497 15286 32509
rect 15338 32497 15344 32549
rect 6544 32389 6550 32401
rect 6432 32361 6550 32389
rect 6544 32349 6550 32361
rect 6602 32349 6608 32401
rect 50896 32241 50902 32253
rect 7296 32213 50902 32241
rect 50896 32201 50902 32213
rect 50954 32201 50960 32253
rect 42832 32167 42838 32179
rect 6912 32139 42838 32167
rect 42832 32127 42838 32139
rect 42890 32127 42896 32179
rect 13072 32093 13078 32105
rect 13033 32065 13078 32093
rect 13072 32053 13078 32065
rect 13130 32053 13136 32105
rect 1152 31994 58848 32016
rect 1152 31942 4294 31994
rect 4346 31942 4358 31994
rect 4410 31942 4422 31994
rect 4474 31942 4486 31994
rect 4538 31942 35014 31994
rect 35066 31942 35078 31994
rect 35130 31942 35142 31994
rect 35194 31942 35206 31994
rect 35258 31942 58848 31994
rect 1152 31920 58848 31942
rect 6544 31831 6550 31883
rect 6602 31871 6608 31883
rect 52816 31871 52822 31883
rect 6602 31843 52822 31871
rect 6602 31831 6608 31843
rect 52816 31831 52822 31843
rect 52874 31831 52880 31883
rect 6832 31757 6838 31809
rect 6890 31797 6896 31809
rect 48880 31797 48886 31809
rect 6890 31769 48886 31797
rect 6890 31757 6896 31769
rect 48880 31757 48886 31769
rect 48938 31757 48944 31809
rect 26512 31723 26518 31735
rect 26473 31695 26518 31723
rect 26512 31683 26518 31695
rect 26570 31683 26576 31735
rect 57331 31726 57389 31732
rect 57331 31692 57343 31726
rect 57377 31723 57389 31726
rect 57424 31723 57430 31735
rect 57377 31695 57430 31723
rect 57377 31692 57389 31695
rect 57331 31686 57389 31692
rect 57424 31683 57430 31695
rect 57482 31683 57488 31735
rect 1152 31328 58848 31350
rect 1152 31276 19654 31328
rect 19706 31276 19718 31328
rect 19770 31276 19782 31328
rect 19834 31276 19846 31328
rect 19898 31276 50374 31328
rect 50426 31276 50438 31328
rect 50490 31276 50502 31328
rect 50554 31276 50566 31328
rect 50618 31276 58848 31328
rect 1152 31254 58848 31276
rect 1744 30869 1750 30921
rect 1802 30909 1808 30921
rect 23059 30912 23117 30918
rect 23059 30909 23071 30912
rect 1802 30881 23071 30909
rect 1802 30869 1808 30881
rect 23059 30878 23071 30881
rect 23105 30878 23117 30912
rect 23059 30872 23117 30878
rect 18832 30795 18838 30847
rect 18890 30835 18896 30847
rect 40912 30835 40918 30847
rect 18890 30807 40918 30835
rect 18890 30795 18896 30807
rect 40912 30795 40918 30807
rect 40970 30795 40976 30847
rect 1152 30662 58848 30684
rect 1152 30610 4294 30662
rect 4346 30610 4358 30662
rect 4410 30610 4422 30662
rect 4474 30610 4486 30662
rect 4538 30610 35014 30662
rect 35066 30610 35078 30662
rect 35130 30610 35142 30662
rect 35194 30610 35206 30662
rect 35258 30610 58848 30662
rect 1152 30588 58848 30610
rect 38224 30499 38230 30551
rect 38282 30539 38288 30551
rect 45184 30539 45190 30551
rect 38282 30511 45190 30539
rect 38282 30499 38288 30511
rect 45184 30499 45190 30511
rect 45242 30499 45248 30551
rect 39280 30465 39286 30477
rect 30096 30437 39286 30465
rect 39280 30425 39286 30437
rect 39338 30425 39344 30477
rect 40912 30425 40918 30477
rect 40970 30465 40976 30477
rect 40970 30437 44702 30465
rect 40970 30425 40976 30437
rect 44674 30430 44702 30437
rect 2992 30351 2998 30403
rect 3050 30391 3056 30403
rect 20851 30394 20909 30400
rect 20851 30391 20863 30394
rect 3050 30363 20863 30391
rect 3050 30351 3056 30363
rect 20851 30360 20863 30363
rect 20897 30360 20909 30394
rect 36880 30391 36886 30403
rect 30240 30363 36886 30391
rect 20851 30354 20909 30360
rect 36880 30351 36886 30363
rect 36938 30351 36944 30403
rect 45190 30366 45242 30372
rect 38320 30277 38326 30329
rect 38378 30317 38384 30329
rect 38378 30289 44510 30317
rect 45190 30308 45242 30314
rect 46771 30320 46829 30326
rect 38378 30277 38384 30289
rect 44482 30095 44510 30289
rect 46771 30286 46783 30320
rect 46817 30317 46829 30320
rect 51088 30317 51094 30329
rect 46817 30289 51094 30317
rect 46817 30286 46829 30289
rect 46771 30280 46829 30286
rect 51088 30277 51094 30289
rect 51146 30277 51152 30329
rect 44608 30129 44614 30181
rect 44666 30129 44672 30181
rect 44896 30129 44902 30181
rect 44954 30129 44960 30181
rect 45490 30095 45518 30155
rect 44482 30067 45518 30095
rect 1152 29996 58848 30018
rect 1152 29944 19654 29996
rect 19706 29944 19718 29996
rect 19770 29944 19782 29996
rect 19834 29944 19846 29996
rect 19898 29944 50374 29996
rect 50426 29944 50438 29996
rect 50490 29944 50502 29996
rect 50554 29944 50566 29996
rect 50618 29944 58848 29996
rect 1152 29922 58848 29944
rect 44368 29833 44374 29885
rect 44426 29873 44432 29885
rect 44560 29873 44566 29885
rect 44426 29845 44566 29873
rect 44426 29833 44432 29845
rect 44560 29833 44566 29845
rect 44618 29833 44624 29885
rect 3568 29463 3574 29515
rect 3626 29503 3632 29515
rect 54736 29503 54742 29515
rect 3626 29475 54742 29503
rect 3626 29463 3632 29475
rect 54736 29463 54742 29475
rect 54794 29463 54800 29515
rect 27955 29432 28013 29438
rect 27955 29398 27967 29432
rect 28001 29429 28013 29432
rect 28243 29432 28301 29438
rect 28243 29429 28255 29432
rect 28001 29401 28255 29429
rect 28001 29398 28013 29401
rect 27955 29392 28013 29398
rect 28243 29398 28255 29401
rect 28289 29429 28301 29432
rect 41584 29429 41590 29441
rect 28289 29401 41590 29429
rect 28289 29398 28301 29401
rect 28243 29392 28301 29398
rect 41584 29389 41590 29401
rect 41642 29389 41648 29441
rect 1152 29330 58848 29352
rect 1152 29278 4294 29330
rect 4346 29278 4358 29330
rect 4410 29278 4422 29330
rect 4474 29278 4486 29330
rect 4538 29278 35014 29330
rect 35066 29278 35078 29330
rect 35130 29278 35142 29330
rect 35194 29278 35206 29330
rect 35258 29278 58848 29330
rect 1152 29256 58848 29278
rect 9331 28914 9389 28920
rect 9331 28880 9343 28914
rect 9377 28880 9389 28914
rect 9331 28874 9389 28880
rect 9043 28840 9101 28846
rect 9043 28806 9055 28840
rect 9089 28837 9101 28840
rect 9346 28837 9374 28874
rect 25456 28871 25462 28923
rect 25514 28911 25520 28923
rect 28915 28914 28973 28920
rect 28915 28911 28927 28914
rect 25514 28883 28927 28911
rect 25514 28871 25520 28883
rect 28915 28880 28927 28883
rect 28961 28880 28973 28914
rect 28915 28874 28973 28880
rect 52336 28837 52342 28849
rect 9089 28809 52342 28837
rect 9089 28806 9101 28809
rect 9043 28800 9101 28806
rect 52336 28797 52342 28809
rect 52394 28797 52400 28849
rect 1152 28664 58848 28686
rect 1152 28612 19654 28664
rect 19706 28612 19718 28664
rect 19770 28612 19782 28664
rect 19834 28612 19846 28664
rect 19898 28612 50374 28664
rect 50426 28612 50438 28664
rect 50490 28612 50502 28664
rect 50554 28612 50566 28664
rect 50618 28612 58848 28664
rect 1152 28590 58848 28612
rect 37744 28501 37750 28553
rect 37802 28541 37808 28553
rect 46387 28544 46445 28550
rect 46387 28541 46399 28544
rect 37802 28513 46399 28541
rect 37802 28501 37808 28513
rect 46387 28510 46399 28513
rect 46433 28541 46445 28544
rect 46433 28513 46622 28541
rect 46433 28510 46445 28513
rect 46387 28504 46445 28510
rect 46594 28402 46622 28513
rect 46579 28396 46637 28402
rect 46579 28362 46591 28396
rect 46625 28362 46637 28396
rect 46579 28356 46637 28362
rect 3664 28279 3670 28331
rect 3722 28319 3728 28331
rect 53872 28319 53878 28331
rect 3722 28291 53878 28319
rect 3722 28279 3728 28291
rect 53872 28279 53878 28291
rect 53930 28279 53936 28331
rect 13648 28205 13654 28257
rect 13706 28245 13712 28257
rect 38035 28248 38093 28254
rect 38035 28245 38047 28248
rect 13706 28217 38047 28245
rect 13706 28205 13712 28217
rect 38035 28214 38047 28217
rect 38081 28245 38093 28248
rect 38131 28248 38189 28254
rect 38131 28245 38143 28248
rect 38081 28217 38143 28245
rect 38081 28214 38093 28217
rect 38035 28208 38093 28214
rect 38131 28214 38143 28217
rect 38177 28214 38189 28248
rect 38131 28208 38189 28214
rect 6256 28097 6262 28109
rect 6217 28069 6262 28097
rect 6256 28057 6262 28069
rect 6314 28057 6320 28109
rect 15184 28057 15190 28109
rect 15242 28097 15248 28109
rect 26800 28097 26806 28109
rect 15242 28069 26806 28097
rect 15242 28057 15248 28069
rect 26800 28057 26806 28069
rect 26858 28057 26864 28109
rect 55984 28057 55990 28109
rect 56042 28097 56048 28109
rect 57331 28100 57389 28106
rect 57331 28097 57343 28100
rect 56042 28069 57343 28097
rect 56042 28057 56048 28069
rect 57331 28066 57343 28069
rect 57377 28066 57389 28100
rect 58000 28097 58006 28109
rect 57961 28069 58006 28097
rect 57331 28060 57389 28066
rect 58000 28057 58006 28069
rect 58058 28057 58064 28109
rect 1152 27998 58848 28020
rect 1152 27946 4294 27998
rect 4346 27946 4358 27998
rect 4410 27946 4422 27998
rect 4474 27946 4486 27998
rect 4538 27946 35014 27998
rect 35066 27946 35078 27998
rect 35130 27946 35142 27998
rect 35194 27946 35206 27998
rect 35258 27946 58848 27998
rect 1152 27924 58848 27946
rect 27184 27835 27190 27887
rect 27242 27875 27248 27887
rect 58000 27875 58006 27887
rect 27242 27847 58006 27875
rect 27242 27835 27248 27847
rect 58000 27835 58006 27847
rect 58058 27835 58064 27887
rect 1152 27332 58848 27354
rect 1152 27280 19654 27332
rect 19706 27280 19718 27332
rect 19770 27280 19782 27332
rect 19834 27280 19846 27332
rect 19898 27280 50374 27332
rect 50426 27280 50438 27332
rect 50490 27280 50502 27332
rect 50554 27280 50566 27332
rect 50618 27280 58848 27332
rect 1152 27258 58848 27280
rect 37747 27064 37805 27070
rect 37747 27030 37759 27064
rect 37793 27061 37805 27064
rect 38035 27064 38093 27070
rect 38035 27061 38047 27064
rect 37793 27033 38047 27061
rect 37793 27030 37805 27033
rect 37747 27024 37805 27030
rect 38035 27030 38047 27033
rect 38081 27061 38093 27064
rect 43888 27061 43894 27073
rect 38081 27033 43894 27061
rect 38081 27030 38093 27033
rect 38035 27024 38093 27030
rect 43888 27021 43894 27033
rect 43946 27021 43952 27073
rect 26512 26873 26518 26925
rect 26570 26913 26576 26925
rect 46384 26913 46390 26925
rect 26570 26885 46390 26913
rect 26570 26873 26576 26885
rect 46384 26873 46390 26885
rect 46442 26873 46448 26925
rect 6544 26799 6550 26851
rect 6602 26839 6608 26851
rect 32752 26839 32758 26851
rect 6602 26811 32758 26839
rect 6602 26799 6608 26811
rect 32752 26799 32758 26811
rect 32810 26799 32816 26851
rect 48208 26839 48214 26851
rect 37426 26811 48214 26839
rect 12499 26768 12557 26774
rect 12499 26734 12511 26768
rect 12545 26765 12557 26768
rect 37426 26765 37454 26811
rect 48208 26799 48214 26811
rect 48266 26799 48272 26851
rect 12545 26737 37454 26765
rect 12545 26734 12557 26737
rect 12499 26728 12557 26734
rect 1152 26666 58848 26688
rect 1152 26614 4294 26666
rect 4346 26614 4358 26666
rect 4410 26614 4422 26666
rect 4474 26614 4486 26666
rect 4538 26614 35014 26666
rect 35066 26614 35078 26666
rect 35130 26614 35142 26666
rect 35194 26614 35206 26666
rect 35258 26614 58848 26666
rect 1152 26592 58848 26614
rect 40144 26247 40150 26259
rect 40105 26219 40150 26247
rect 40144 26207 40150 26219
rect 40202 26207 40208 26259
rect 47728 26247 47734 26259
rect 47689 26219 47734 26247
rect 47728 26207 47734 26219
rect 47786 26207 47792 26259
rect 54256 26207 54262 26259
rect 54314 26247 54320 26259
rect 54643 26250 54701 26256
rect 54643 26247 54655 26250
rect 54314 26219 54655 26247
rect 54314 26207 54320 26219
rect 54643 26216 54655 26219
rect 54689 26216 54701 26250
rect 54643 26210 54701 26216
rect 1152 26000 58848 26022
rect 1152 25948 19654 26000
rect 19706 25948 19718 26000
rect 19770 25948 19782 26000
rect 19834 25948 19846 26000
rect 19898 25948 50374 26000
rect 50426 25948 50438 26000
rect 50490 25948 50502 26000
rect 50554 25948 50566 26000
rect 50618 25948 58848 26000
rect 1152 25926 58848 25948
rect 13555 25732 13613 25738
rect 13555 25698 13567 25732
rect 13601 25729 13613 25732
rect 13840 25729 13846 25741
rect 13601 25701 13846 25729
rect 13601 25698 13613 25701
rect 13555 25692 13613 25698
rect 13840 25689 13846 25701
rect 13898 25689 13904 25741
rect 10864 25541 10870 25593
rect 10922 25581 10928 25593
rect 30064 25581 30070 25593
rect 10922 25553 30070 25581
rect 10922 25541 10928 25553
rect 30064 25541 30070 25553
rect 30122 25541 30128 25593
rect 4435 25510 4493 25516
rect 4435 25476 4447 25510
rect 4481 25507 4493 25510
rect 4723 25510 4781 25516
rect 4723 25507 4735 25510
rect 4481 25479 4735 25507
rect 4481 25476 4493 25479
rect 4435 25470 4493 25476
rect 4723 25476 4735 25479
rect 4769 25507 4781 25510
rect 22096 25507 22102 25519
rect 4769 25479 22102 25507
rect 4769 25476 4781 25479
rect 4723 25470 4781 25476
rect 22096 25467 22102 25479
rect 22154 25467 22160 25519
rect 5392 25433 5398 25445
rect 5353 25405 5398 25433
rect 5392 25393 5398 25405
rect 5450 25393 5456 25445
rect 36976 25393 36982 25445
rect 37034 25433 37040 25445
rect 39763 25436 39821 25442
rect 39763 25433 39775 25436
rect 37034 25405 39775 25433
rect 37034 25393 37040 25405
rect 39763 25402 39775 25405
rect 39809 25402 39821 25436
rect 39763 25396 39821 25402
rect 1152 25334 58848 25356
rect 1152 25282 4294 25334
rect 4346 25282 4358 25334
rect 4410 25282 4422 25334
rect 4474 25282 4486 25334
rect 4538 25282 35014 25334
rect 35066 25282 35078 25334
rect 35130 25282 35142 25334
rect 35194 25282 35206 25334
rect 35258 25282 58848 25334
rect 1152 25260 58848 25282
rect 13552 25171 13558 25223
rect 13610 25211 13616 25223
rect 36304 25211 36310 25223
rect 13610 25183 36310 25211
rect 13610 25171 13616 25183
rect 36304 25171 36310 25183
rect 36362 25171 36368 25223
rect 40144 25171 40150 25223
rect 40202 25211 40208 25223
rect 51472 25211 51478 25223
rect 40202 25183 51478 25211
rect 40202 25171 40208 25183
rect 51472 25171 51478 25183
rect 51530 25171 51536 25223
rect 5392 25097 5398 25149
rect 5450 25137 5456 25149
rect 45232 25137 45238 25149
rect 5450 25109 45238 25137
rect 5450 25097 5456 25109
rect 45232 25097 45238 25109
rect 45290 25097 45296 25149
rect 15667 24992 15725 24998
rect 15667 24958 15679 24992
rect 15713 24989 15725 24992
rect 30640 24989 30646 25001
rect 15713 24961 30646 24989
rect 15713 24958 15725 24961
rect 15667 24952 15725 24958
rect 30640 24949 30646 24961
rect 30698 24949 30704 25001
rect 26611 24918 26669 24924
rect 26611 24884 26623 24918
rect 26657 24915 26669 24918
rect 26899 24918 26957 24924
rect 26899 24915 26911 24918
rect 26657 24887 26911 24915
rect 26657 24884 26669 24887
rect 26611 24878 26669 24884
rect 26899 24884 26911 24887
rect 26945 24884 26957 24918
rect 26899 24878 26957 24884
rect 26914 24767 26942 24878
rect 31696 24875 31702 24927
rect 31754 24915 31760 24927
rect 36691 24918 36749 24924
rect 36691 24915 36703 24918
rect 31754 24887 36703 24915
rect 31754 24875 31760 24887
rect 36691 24884 36703 24887
rect 36737 24884 36749 24918
rect 36691 24878 36749 24884
rect 38704 24767 38710 24779
rect 26914 24739 38710 24767
rect 38704 24727 38710 24739
rect 38762 24727 38768 24779
rect 1152 24668 58848 24690
rect 1152 24616 19654 24668
rect 19706 24616 19718 24668
rect 19770 24616 19782 24668
rect 19834 24616 19846 24668
rect 19898 24616 50374 24668
rect 50426 24616 50438 24668
rect 50490 24616 50502 24668
rect 50554 24616 50566 24668
rect 50618 24616 58848 24668
rect 1152 24594 58848 24616
rect 1152 24002 58848 24024
rect 1152 23950 4294 24002
rect 4346 23950 4358 24002
rect 4410 23950 4422 24002
rect 4474 23950 4486 24002
rect 4538 23950 35014 24002
rect 35066 23950 35078 24002
rect 35130 23950 35142 24002
rect 35194 23950 35206 24002
rect 35258 23950 58848 24002
rect 1152 23928 58848 23950
rect 1936 23691 1942 23743
rect 1994 23731 2000 23743
rect 36880 23731 36886 23743
rect 1994 23703 36886 23731
rect 1994 23691 2000 23703
rect 36880 23691 36886 23703
rect 36938 23691 36944 23743
rect 8560 23583 8566 23595
rect 8521 23555 8566 23583
rect 8560 23543 8566 23555
rect 8618 23543 8624 23595
rect 13648 23583 13654 23595
rect 13609 23555 13654 23583
rect 13648 23543 13654 23555
rect 13706 23543 13712 23595
rect 41875 23586 41933 23592
rect 41875 23583 41887 23586
rect 27346 23555 41887 23583
rect 26992 23469 26998 23521
rect 27050 23509 27056 23521
rect 27346 23509 27374 23555
rect 41875 23552 41887 23555
rect 41921 23552 41933 23586
rect 41875 23546 41933 23552
rect 45523 23586 45581 23592
rect 45523 23552 45535 23586
rect 45569 23552 45581 23586
rect 45523 23546 45581 23552
rect 27050 23481 27374 23509
rect 27050 23469 27056 23481
rect 7120 23395 7126 23447
rect 7178 23435 7184 23447
rect 45538 23435 45566 23546
rect 7178 23407 45566 23435
rect 7178 23395 7184 23407
rect 1152 23336 58848 23358
rect 1152 23284 19654 23336
rect 19706 23284 19718 23336
rect 19770 23284 19782 23336
rect 19834 23284 19846 23336
rect 19898 23284 50374 23336
rect 50426 23284 50438 23336
rect 50490 23284 50502 23336
rect 50554 23284 50566 23336
rect 50618 23284 58848 23336
rect 1152 23262 58848 23284
rect 20467 23068 20525 23074
rect 20467 23034 20479 23068
rect 20513 23065 20525 23068
rect 20755 23068 20813 23074
rect 20755 23065 20767 23068
rect 20513 23037 20767 23065
rect 20513 23034 20525 23037
rect 20467 23028 20525 23034
rect 20755 23034 20767 23037
rect 20801 23065 20813 23068
rect 57328 23065 57334 23077
rect 20801 23037 57334 23065
rect 20801 23034 20813 23037
rect 20755 23028 20813 23034
rect 57328 23025 57334 23037
rect 57386 23025 57392 23077
rect 33808 22951 33814 23003
rect 33866 22991 33872 23003
rect 38800 22991 38806 23003
rect 33866 22963 38806 22991
rect 33866 22951 33872 22963
rect 38800 22951 38806 22963
rect 38858 22951 38864 23003
rect 8659 22772 8717 22778
rect 8659 22738 8671 22772
rect 8705 22769 8717 22772
rect 8752 22769 8758 22781
rect 8705 22741 8758 22769
rect 8705 22738 8717 22741
rect 8659 22732 8717 22738
rect 8752 22729 8758 22741
rect 8810 22729 8816 22781
rect 19408 22729 19414 22781
rect 19466 22769 19472 22781
rect 24019 22772 24077 22778
rect 24019 22769 24031 22772
rect 19466 22741 24031 22769
rect 19466 22729 19472 22741
rect 24019 22738 24031 22741
rect 24065 22738 24077 22772
rect 36304 22769 36310 22781
rect 36265 22741 36310 22769
rect 24019 22732 24077 22738
rect 36304 22729 36310 22741
rect 36362 22729 36368 22781
rect 49360 22729 49366 22781
rect 49418 22769 49424 22781
rect 57331 22772 57389 22778
rect 57331 22769 57343 22772
rect 49418 22741 57343 22769
rect 49418 22729 49424 22741
rect 57331 22738 57343 22741
rect 57377 22738 57389 22772
rect 57331 22732 57389 22738
rect 1152 22670 58848 22692
rect 1152 22618 4294 22670
rect 4346 22618 4358 22670
rect 4410 22618 4422 22670
rect 4474 22618 4486 22670
rect 4538 22618 35014 22670
rect 35066 22618 35078 22670
rect 35130 22618 35142 22670
rect 35194 22618 35206 22670
rect 35258 22618 58848 22670
rect 1152 22596 58848 22618
rect 8560 22433 8566 22485
rect 8618 22473 8624 22485
rect 33232 22473 33238 22485
rect 8618 22445 33238 22473
rect 8618 22433 8624 22445
rect 33232 22433 33238 22445
rect 33290 22433 33296 22485
rect 13648 22359 13654 22411
rect 13706 22399 13712 22411
rect 40048 22399 40054 22411
rect 13706 22371 40054 22399
rect 13706 22359 13712 22371
rect 40048 22359 40054 22371
rect 40106 22359 40112 22411
rect 7888 22285 7894 22337
rect 7946 22325 7952 22337
rect 54928 22325 54934 22337
rect 7946 22297 54934 22325
rect 7946 22285 7952 22297
rect 54928 22285 54934 22297
rect 54986 22285 54992 22337
rect 15088 22251 15094 22263
rect 15049 22223 15094 22251
rect 15088 22211 15094 22223
rect 15146 22211 15152 22263
rect 20563 22254 20621 22260
rect 20563 22220 20575 22254
rect 20609 22251 20621 22254
rect 22864 22251 22870 22263
rect 20609 22223 22870 22251
rect 20609 22220 20621 22223
rect 20563 22214 20621 22220
rect 22864 22211 22870 22223
rect 22922 22211 22928 22263
rect 25552 22211 25558 22263
rect 25610 22251 25616 22263
rect 34963 22254 35021 22260
rect 34963 22251 34975 22254
rect 25610 22223 34975 22251
rect 25610 22211 25616 22223
rect 34963 22220 34975 22223
rect 35009 22220 35021 22254
rect 34963 22214 35021 22220
rect 1152 22004 58848 22026
rect 1152 21952 19654 22004
rect 19706 21952 19718 22004
rect 19770 21952 19782 22004
rect 19834 21952 19846 22004
rect 19898 21952 50374 22004
rect 50426 21952 50438 22004
rect 50490 21952 50502 22004
rect 50554 21952 50566 22004
rect 50618 21952 58848 22004
rect 1152 21930 58848 21952
rect 26608 21619 26614 21671
rect 26666 21659 26672 21671
rect 28144 21659 28150 21671
rect 26666 21631 28150 21659
rect 26666 21619 26672 21631
rect 28144 21619 28150 21631
rect 28202 21619 28208 21671
rect 38128 21545 38134 21597
rect 38186 21585 38192 21597
rect 39472 21585 39478 21597
rect 38186 21557 39478 21585
rect 38186 21545 38192 21557
rect 39472 21545 39478 21557
rect 39530 21545 39536 21597
rect 5107 21440 5165 21446
rect 5107 21406 5119 21440
rect 5153 21437 5165 21440
rect 9424 21437 9430 21449
rect 5153 21409 9430 21437
rect 5153 21406 5165 21409
rect 5107 21400 5165 21406
rect 9424 21397 9430 21409
rect 9482 21397 9488 21449
rect 15091 21440 15149 21446
rect 15091 21406 15103 21440
rect 15137 21437 15149 21440
rect 38416 21437 38422 21449
rect 15137 21409 38422 21437
rect 15137 21406 15149 21409
rect 15091 21400 15149 21406
rect 38416 21397 38422 21409
rect 38474 21397 38480 21449
rect 1152 21338 58848 21360
rect 1152 21286 4294 21338
rect 4346 21286 4358 21338
rect 4410 21286 4422 21338
rect 4474 21286 4486 21338
rect 4538 21286 35014 21338
rect 35066 21286 35078 21338
rect 35130 21286 35142 21338
rect 35194 21286 35206 21338
rect 35258 21286 58848 21338
rect 1152 21264 58848 21286
rect 23026 21113 37454 21141
rect 13072 20953 13078 21005
rect 13130 20993 13136 21005
rect 23026 20993 23054 21113
rect 25072 21027 25078 21079
rect 25130 21067 25136 21079
rect 25130 21039 37310 21067
rect 25130 21027 25136 21039
rect 13130 20965 23054 20993
rect 13130 20953 13136 20965
rect 26224 20879 26230 20931
rect 26282 20919 26288 20931
rect 37075 20922 37133 20928
rect 37075 20919 37087 20922
rect 26282 20891 37087 20919
rect 26282 20879 26288 20891
rect 37075 20888 37087 20891
rect 37121 20888 37133 20922
rect 37282 20919 37310 21039
rect 37426 20993 37454 21113
rect 46768 20993 46774 21005
rect 37426 20965 46774 20993
rect 46768 20953 46774 20965
rect 46826 20953 46832 21005
rect 47635 20922 47693 20928
rect 47635 20919 47647 20922
rect 37282 20891 47647 20919
rect 37075 20882 37133 20888
rect 47635 20888 47647 20891
rect 47681 20919 47693 20922
rect 47731 20922 47789 20928
rect 47731 20919 47743 20922
rect 47681 20891 47743 20919
rect 47681 20888 47693 20891
rect 47635 20882 47693 20888
rect 47731 20888 47743 20891
rect 47777 20888 47789 20922
rect 47731 20882 47789 20888
rect 1152 20672 58848 20694
rect 1152 20620 19654 20672
rect 19706 20620 19718 20672
rect 19770 20620 19782 20672
rect 19834 20620 19846 20672
rect 19898 20620 50374 20672
rect 50426 20620 50438 20672
rect 50490 20620 50502 20672
rect 50554 20620 50566 20672
rect 50618 20620 58848 20672
rect 1152 20598 58848 20620
rect 24496 20139 24502 20191
rect 24554 20179 24560 20191
rect 26704 20179 26710 20191
rect 24554 20151 26710 20179
rect 24554 20139 24560 20151
rect 26704 20139 26710 20151
rect 26762 20139 26768 20191
rect 5968 20065 5974 20117
rect 6026 20105 6032 20117
rect 23152 20105 23158 20117
rect 6026 20077 23158 20105
rect 6026 20065 6032 20077
rect 23152 20065 23158 20077
rect 23210 20065 23216 20117
rect 1152 20006 58848 20028
rect 1152 19954 4294 20006
rect 4346 19954 4358 20006
rect 4410 19954 4422 20006
rect 4474 19954 4486 20006
rect 4538 19954 35014 20006
rect 35066 19954 35078 20006
rect 35130 19954 35142 20006
rect 35194 19954 35206 20006
rect 35258 19954 58848 20006
rect 1152 19932 58848 19954
rect 7987 19812 8045 19818
rect 7987 19778 7999 19812
rect 8033 19809 8045 19812
rect 19216 19809 19222 19821
rect 8033 19781 19222 19809
rect 8033 19778 8045 19781
rect 7987 19772 8045 19778
rect 19216 19769 19222 19781
rect 19274 19769 19280 19821
rect 6160 19695 6166 19747
rect 6218 19735 6224 19747
rect 20848 19735 20854 19747
rect 6218 19707 20854 19735
rect 6218 19695 6224 19707
rect 20848 19695 20854 19707
rect 20906 19695 20912 19747
rect 25648 19621 25654 19673
rect 25706 19661 25712 19673
rect 25706 19633 37454 19661
rect 25706 19621 25712 19633
rect 1747 19590 1805 19596
rect 1747 19556 1759 19590
rect 1793 19587 1805 19590
rect 4144 19587 4150 19599
rect 1793 19559 4150 19587
rect 1793 19556 1805 19559
rect 1747 19550 1805 19556
rect 4144 19547 4150 19559
rect 4202 19547 4208 19599
rect 8467 19590 8525 19596
rect 8467 19556 8479 19590
rect 8513 19556 8525 19590
rect 13936 19587 13942 19599
rect 13897 19559 13942 19587
rect 8467 19550 8525 19556
rect 6448 19473 6454 19525
rect 6506 19513 6512 19525
rect 8482 19513 8510 19550
rect 13936 19547 13942 19559
rect 13994 19547 14000 19599
rect 28240 19587 28246 19599
rect 28201 19559 28246 19587
rect 28240 19547 28246 19559
rect 28298 19547 28304 19599
rect 37426 19587 37454 19633
rect 38899 19590 38957 19596
rect 38899 19587 38911 19590
rect 37426 19559 38911 19587
rect 38899 19556 38911 19559
rect 38945 19556 38957 19590
rect 38899 19550 38957 19556
rect 36784 19513 36790 19525
rect 6506 19485 8414 19513
rect 8482 19485 36790 19513
rect 6506 19473 6512 19485
rect 5872 19399 5878 19451
rect 5930 19439 5936 19451
rect 7987 19442 8045 19448
rect 7987 19439 7999 19442
rect 5930 19411 7999 19439
rect 5930 19399 5936 19411
rect 7987 19408 7999 19411
rect 8033 19408 8045 19442
rect 8386 19439 8414 19485
rect 36784 19473 36790 19485
rect 36842 19473 36848 19525
rect 17872 19439 17878 19451
rect 8386 19411 17878 19439
rect 7987 19402 8045 19408
rect 17872 19399 17878 19411
rect 17930 19399 17936 19451
rect 22864 19399 22870 19451
rect 22922 19439 22928 19451
rect 49072 19439 49078 19451
rect 22922 19411 49078 19439
rect 22922 19399 22928 19411
rect 49072 19399 49078 19411
rect 49130 19399 49136 19451
rect 1152 19340 58848 19362
rect 1152 19288 19654 19340
rect 19706 19288 19718 19340
rect 19770 19288 19782 19340
rect 19834 19288 19846 19340
rect 19898 19288 50374 19340
rect 50426 19288 50438 19340
rect 50490 19288 50502 19340
rect 50554 19288 50566 19340
rect 50618 19288 58848 19340
rect 1152 19266 58848 19288
rect 5968 19177 5974 19229
rect 6026 19177 6032 19229
rect 5824 19103 5830 19155
rect 5882 19103 5888 19155
rect 5491 18850 5549 18856
rect 5491 18816 5503 18850
rect 5537 18847 5549 18850
rect 5986 18847 6014 19177
rect 6112 19103 6118 19155
rect 6170 19103 6176 19155
rect 6400 19103 6406 19155
rect 6458 19103 6464 19155
rect 16048 19143 16054 19155
rect 6720 19115 16054 19143
rect 16048 19103 16054 19115
rect 16106 19103 16112 19155
rect 47728 18955 47734 19007
rect 47786 18995 47792 19007
rect 49936 18995 49942 19007
rect 47786 18967 49942 18995
rect 47786 18955 47792 18967
rect 49936 18955 49942 18967
rect 49994 18955 50000 19007
rect 5537 18819 6014 18847
rect 5537 18816 5549 18819
rect 5491 18810 5549 18816
rect 30256 18733 30262 18785
rect 30314 18773 30320 18785
rect 37648 18773 37654 18785
rect 30314 18745 37654 18773
rect 30314 18733 30320 18745
rect 37648 18733 37654 18745
rect 37706 18733 37712 18785
rect 1152 18674 58848 18696
rect 1152 18622 4294 18674
rect 4346 18622 4358 18674
rect 4410 18622 4422 18674
rect 4474 18622 4486 18674
rect 4538 18622 35014 18674
rect 35066 18622 35078 18674
rect 35130 18622 35142 18674
rect 35194 18622 35206 18674
rect 35258 18622 58848 18674
rect 1152 18600 58848 18622
rect 28816 18215 28822 18267
rect 28874 18255 28880 18267
rect 34003 18258 34061 18264
rect 34003 18255 34015 18258
rect 28874 18227 34015 18255
rect 28874 18215 28880 18227
rect 34003 18224 34015 18227
rect 34049 18224 34061 18258
rect 34003 18218 34061 18224
rect 13936 18067 13942 18119
rect 13994 18107 14000 18119
rect 46576 18107 46582 18119
rect 13994 18079 46582 18107
rect 13994 18067 14000 18079
rect 46576 18067 46582 18079
rect 46634 18067 46640 18119
rect 1152 18008 58848 18030
rect 1152 17956 19654 18008
rect 19706 17956 19718 18008
rect 19770 17956 19782 18008
rect 19834 17956 19846 18008
rect 19898 17956 50374 18008
rect 50426 17956 50438 18008
rect 50490 17956 50502 18008
rect 50554 17956 50566 18008
rect 50618 17956 58848 18008
rect 1152 17934 58848 17956
rect 20752 17771 20758 17823
rect 20810 17811 20816 17823
rect 23248 17811 23254 17823
rect 20810 17783 23254 17811
rect 20810 17771 20816 17783
rect 23248 17771 23254 17783
rect 23306 17771 23312 17823
rect 11920 17549 11926 17601
rect 11978 17589 11984 17601
rect 27091 17592 27149 17598
rect 27091 17589 27103 17592
rect 11978 17561 27103 17589
rect 11978 17549 11984 17561
rect 27091 17558 27103 17561
rect 27137 17589 27149 17592
rect 27283 17592 27341 17598
rect 27283 17589 27295 17592
rect 27137 17561 27295 17589
rect 27137 17558 27149 17561
rect 27091 17552 27149 17558
rect 27283 17558 27295 17561
rect 27329 17558 27341 17592
rect 27283 17552 27341 17558
rect 37456 17475 37462 17527
rect 37514 17515 37520 17527
rect 54067 17518 54125 17524
rect 54067 17515 54079 17518
rect 37514 17487 54079 17515
rect 37514 17475 37520 17487
rect 54067 17484 54079 17487
rect 54113 17484 54125 17518
rect 54067 17478 54125 17484
rect 23152 17441 23158 17453
rect 23113 17413 23158 17441
rect 23152 17401 23158 17413
rect 23210 17401 23216 17453
rect 41488 17401 41494 17453
rect 41546 17441 41552 17453
rect 46771 17444 46829 17450
rect 46771 17441 46783 17444
rect 41546 17413 46783 17441
rect 41546 17401 41552 17413
rect 46771 17410 46783 17413
rect 46817 17410 46829 17444
rect 46771 17404 46829 17410
rect 1152 17342 58848 17364
rect 1152 17290 4294 17342
rect 4346 17290 4358 17342
rect 4410 17290 4422 17342
rect 4474 17290 4486 17342
rect 4538 17290 35014 17342
rect 35066 17290 35078 17342
rect 35130 17290 35142 17342
rect 35194 17290 35206 17342
rect 35258 17290 58848 17342
rect 1152 17268 58848 17290
rect 2803 17000 2861 17006
rect 2803 16966 2815 17000
rect 2849 16997 2861 17000
rect 3091 17000 3149 17006
rect 3091 16997 3103 17000
rect 2849 16969 3103 16997
rect 2849 16966 2861 16969
rect 2803 16960 2861 16966
rect 3091 16966 3103 16969
rect 3137 16997 3149 17000
rect 34384 16997 34390 17009
rect 3137 16969 34390 16997
rect 3137 16966 3149 16969
rect 3091 16960 3149 16966
rect 34384 16957 34390 16969
rect 34442 16957 34448 17009
rect 10483 16926 10541 16932
rect 10483 16892 10495 16926
rect 10529 16923 10541 16926
rect 16528 16923 16534 16935
rect 10529 16895 16534 16923
rect 10529 16892 10541 16895
rect 10483 16886 10541 16892
rect 16528 16883 16534 16895
rect 16586 16883 16592 16935
rect 31504 16883 31510 16935
rect 31562 16923 31568 16935
rect 35539 16926 35597 16932
rect 35539 16923 35551 16926
rect 31562 16895 35551 16923
rect 31562 16883 31568 16895
rect 35539 16892 35551 16895
rect 35585 16892 35597 16926
rect 46099 16926 46157 16932
rect 46099 16923 46111 16926
rect 35539 16886 35597 16892
rect 37426 16895 46111 16923
rect 29488 16809 29494 16861
rect 29546 16849 29552 16861
rect 37426 16849 37454 16895
rect 46099 16892 46111 16895
rect 46145 16892 46157 16926
rect 54640 16923 54646 16935
rect 54601 16895 54646 16923
rect 46099 16886 46157 16892
rect 54640 16883 54646 16895
rect 54698 16883 54704 16935
rect 29546 16821 37454 16849
rect 29546 16809 29552 16821
rect 10192 16735 10198 16787
rect 10250 16775 10256 16787
rect 28816 16775 28822 16787
rect 10250 16747 28822 16775
rect 10250 16735 10256 16747
rect 28816 16735 28822 16747
rect 28874 16735 28880 16787
rect 38896 16735 38902 16787
rect 38954 16775 38960 16787
rect 54448 16775 54454 16787
rect 38954 16747 54454 16775
rect 38954 16735 38960 16747
rect 54448 16735 54454 16747
rect 54506 16735 54512 16787
rect 1152 16676 58848 16698
rect 1152 16624 19654 16676
rect 19706 16624 19718 16676
rect 19770 16624 19782 16676
rect 19834 16624 19846 16676
rect 19898 16624 50374 16676
rect 50426 16624 50438 16676
rect 50490 16624 50502 16676
rect 50554 16624 50566 16676
rect 50618 16624 58848 16676
rect 1152 16602 58848 16624
rect 19024 16513 19030 16565
rect 19082 16553 19088 16565
rect 39856 16553 39862 16565
rect 19082 16525 39862 16553
rect 19082 16513 19088 16525
rect 39856 16513 39862 16525
rect 39914 16513 39920 16565
rect 53491 16260 53549 16266
rect 53491 16226 53503 16260
rect 53537 16226 53549 16260
rect 53491 16220 53549 16226
rect 21712 16069 21718 16121
rect 21770 16109 21776 16121
rect 53299 16112 53357 16118
rect 53299 16109 53311 16112
rect 21770 16081 53311 16109
rect 21770 16069 21776 16081
rect 53299 16078 53311 16081
rect 53345 16109 53357 16112
rect 53506 16109 53534 16220
rect 53345 16081 53534 16109
rect 53345 16078 53357 16081
rect 53299 16072 53357 16078
rect 1152 16010 58848 16032
rect 1152 15958 4294 16010
rect 4346 15958 4358 16010
rect 4410 15958 4422 16010
rect 4474 15958 4486 16010
rect 4538 15958 35014 16010
rect 35066 15958 35078 16010
rect 35130 15958 35142 16010
rect 35194 15958 35206 16010
rect 35258 15958 58848 16010
rect 1152 15936 58848 15958
rect 9811 15890 9869 15896
rect 9811 15856 9823 15890
rect 9857 15887 9869 15890
rect 15856 15887 15862 15899
rect 9857 15859 15862 15887
rect 9857 15856 9869 15859
rect 9811 15850 9869 15856
rect 15856 15847 15862 15859
rect 15914 15847 15920 15899
rect 15088 15699 15094 15751
rect 15146 15739 15152 15751
rect 26416 15739 26422 15751
rect 15146 15711 26422 15739
rect 15146 15699 15152 15711
rect 26416 15699 26422 15711
rect 26474 15699 26480 15751
rect 22480 15625 22486 15677
rect 22538 15665 22544 15677
rect 34864 15665 34870 15677
rect 22538 15637 34870 15665
rect 22538 15625 22544 15637
rect 34864 15625 34870 15637
rect 34922 15625 34928 15677
rect 18928 15551 18934 15603
rect 18986 15591 18992 15603
rect 44656 15591 44662 15603
rect 18986 15563 44662 15591
rect 18986 15551 18992 15563
rect 44656 15551 44662 15563
rect 44714 15551 44720 15603
rect 15472 15477 15478 15529
rect 15530 15517 15536 15529
rect 41296 15517 41302 15529
rect 15530 15489 41302 15517
rect 15530 15477 15536 15489
rect 41296 15477 41302 15489
rect 41354 15477 41360 15529
rect 18544 15403 18550 15455
rect 18602 15443 18608 15455
rect 44944 15443 44950 15455
rect 18602 15415 44950 15443
rect 18602 15403 18608 15415
rect 44944 15403 44950 15415
rect 45002 15403 45008 15455
rect 1152 15344 58848 15366
rect 1152 15292 19654 15344
rect 19706 15292 19718 15344
rect 19770 15292 19782 15344
rect 19834 15292 19846 15344
rect 19898 15292 50374 15344
rect 50426 15292 50438 15344
rect 50490 15292 50502 15344
rect 50554 15292 50566 15344
rect 50618 15292 58848 15344
rect 1152 15270 58848 15292
rect 18064 15181 18070 15233
rect 18122 15221 18128 15233
rect 53968 15221 53974 15233
rect 18122 15193 53974 15221
rect 18122 15181 18128 15193
rect 53968 15181 53974 15193
rect 54026 15181 54032 15233
rect 15856 15107 15862 15159
rect 15914 15147 15920 15159
rect 52624 15147 52630 15159
rect 15914 15119 52630 15147
rect 15914 15107 15920 15119
rect 52624 15107 52630 15119
rect 52682 15107 52688 15159
rect 32272 14777 32278 14789
rect 32233 14749 32278 14777
rect 32272 14737 32278 14749
rect 32330 14737 32336 14789
rect 1152 14678 58848 14700
rect 1152 14626 4294 14678
rect 4346 14626 4358 14678
rect 4410 14626 4422 14678
rect 4474 14626 4486 14678
rect 4538 14626 35014 14678
rect 35066 14626 35078 14678
rect 35130 14626 35142 14678
rect 35194 14626 35206 14678
rect 35258 14626 58848 14678
rect 1152 14604 58848 14626
rect 11536 14515 11542 14567
rect 11594 14555 11600 14567
rect 17968 14555 17974 14567
rect 11594 14527 17974 14555
rect 11594 14515 11600 14527
rect 17968 14515 17974 14527
rect 18026 14515 18032 14567
rect 41200 14515 41206 14567
rect 41258 14555 41264 14567
rect 42256 14555 42262 14567
rect 41258 14527 42262 14555
rect 41258 14515 41264 14527
rect 42256 14515 42262 14527
rect 42314 14515 42320 14567
rect 44752 14515 44758 14567
rect 44810 14555 44816 14567
rect 48979 14558 49037 14564
rect 48979 14555 48991 14558
rect 44810 14527 48991 14555
rect 44810 14515 44816 14527
rect 48979 14524 48991 14527
rect 49025 14555 49037 14558
rect 49171 14558 49229 14564
rect 49171 14555 49183 14558
rect 49025 14527 49183 14555
rect 49025 14524 49037 14527
rect 48979 14518 49037 14524
rect 49171 14524 49183 14527
rect 49217 14524 49229 14558
rect 49171 14518 49229 14524
rect 12976 14441 12982 14493
rect 13034 14481 13040 14493
rect 46579 14484 46637 14490
rect 46579 14481 46591 14484
rect 13034 14453 46591 14481
rect 13034 14441 13040 14453
rect 46579 14450 46591 14453
rect 46625 14450 46637 14484
rect 46579 14444 46637 14450
rect 12592 14219 12598 14271
rect 12650 14259 12656 14271
rect 34096 14259 34102 14271
rect 12650 14231 34102 14259
rect 12650 14219 12656 14231
rect 34096 14219 34102 14231
rect 34154 14219 34160 14271
rect 9424 14145 9430 14197
rect 9482 14185 9488 14197
rect 24208 14185 24214 14197
rect 9482 14157 24214 14185
rect 9482 14145 9488 14157
rect 24208 14145 24214 14157
rect 24266 14145 24272 14197
rect 34576 14145 34582 14197
rect 34634 14185 34640 14197
rect 41104 14185 41110 14197
rect 34634 14157 41110 14185
rect 34634 14145 34640 14157
rect 41104 14145 41110 14157
rect 41162 14145 41168 14197
rect 10096 14071 10102 14123
rect 10154 14111 10160 14123
rect 44659 14114 44717 14120
rect 44659 14111 44671 14114
rect 10154 14083 44671 14111
rect 10154 14071 10160 14083
rect 44659 14080 44671 14083
rect 44705 14111 44717 14114
rect 44851 14114 44909 14120
rect 44851 14111 44863 14114
rect 44705 14083 44863 14111
rect 44705 14080 44717 14083
rect 44659 14074 44717 14080
rect 44851 14080 44863 14083
rect 44897 14080 44909 14114
rect 44851 14074 44909 14080
rect 1152 14012 58848 14034
rect 1152 13960 19654 14012
rect 19706 13960 19718 14012
rect 19770 13960 19782 14012
rect 19834 13960 19846 14012
rect 19898 13960 50374 14012
rect 50426 13960 50438 14012
rect 50490 13960 50502 14012
rect 50554 13960 50566 14012
rect 50618 13960 58848 14012
rect 1152 13938 58848 13960
rect 33136 13849 33142 13901
rect 33194 13889 33200 13901
rect 41392 13889 41398 13901
rect 33194 13861 41398 13889
rect 33194 13849 33200 13861
rect 41392 13849 41398 13861
rect 41450 13849 41456 13901
rect 12592 13775 12598 13827
rect 12650 13815 12656 13827
rect 12650 13787 12768 13815
rect 12650 13775 12656 13787
rect 38416 13775 38422 13827
rect 38474 13815 38480 13827
rect 52048 13815 52054 13827
rect 38474 13787 52054 13815
rect 38474 13775 38480 13787
rect 52048 13775 52054 13787
rect 52106 13775 52112 13827
rect 34000 13701 34006 13753
rect 34058 13741 34064 13753
rect 54640 13741 54646 13753
rect 34058 13713 54646 13741
rect 34058 13701 34064 13713
rect 54640 13701 54646 13713
rect 54698 13701 54704 13753
rect 17968 13627 17974 13679
rect 18026 13667 18032 13679
rect 18026 13639 23054 13667
rect 18026 13627 18032 13639
rect 23026 13593 23054 13639
rect 47824 13593 47830 13605
rect 23026 13565 47830 13593
rect 47824 13553 47830 13565
rect 47882 13553 47888 13605
rect 12403 13522 12461 13528
rect 12403 13488 12415 13522
rect 12449 13519 12461 13522
rect 36592 13519 36598 13531
rect 12449 13491 36598 13519
rect 12449 13488 12461 13491
rect 12403 13482 12461 13488
rect 36592 13479 36598 13491
rect 36650 13479 36656 13531
rect 4144 13405 4150 13457
rect 4202 13445 4208 13457
rect 5299 13448 5357 13454
rect 5299 13445 5311 13448
rect 4202 13417 5311 13445
rect 4202 13405 4208 13417
rect 5299 13414 5311 13417
rect 5345 13414 5357 13448
rect 5299 13408 5357 13414
rect 1152 13346 58848 13368
rect 1152 13294 4294 13346
rect 4346 13294 4358 13346
rect 4410 13294 4422 13346
rect 4474 13294 4486 13346
rect 4538 13294 35014 13346
rect 35066 13294 35078 13346
rect 35130 13294 35142 13346
rect 35194 13294 35206 13346
rect 35258 13294 58848 13346
rect 1152 13272 58848 13294
rect 57715 13226 57773 13232
rect 57715 13192 57727 13226
rect 57761 13223 57773 13226
rect 57811 13226 57869 13232
rect 57811 13223 57823 13226
rect 57761 13195 57823 13223
rect 57761 13192 57773 13195
rect 57715 13186 57773 13192
rect 57811 13192 57823 13195
rect 57857 13223 57869 13226
rect 58192 13223 58198 13235
rect 57857 13195 58198 13223
rect 57857 13192 57869 13195
rect 57811 13186 57869 13192
rect 58192 13183 58198 13195
rect 58250 13183 58256 13235
rect 25456 13149 25462 13161
rect 23026 13121 25462 13149
rect 21904 13035 21910 13087
rect 21962 13075 21968 13087
rect 23026 13075 23054 13121
rect 25456 13109 25462 13121
rect 25514 13109 25520 13161
rect 44080 13149 44086 13161
rect 37426 13121 44086 13149
rect 21962 13047 23054 13075
rect 25282 13047 33134 13075
rect 21962 13035 21968 13047
rect 9715 13004 9773 13010
rect 9715 12970 9727 13004
rect 9761 13001 9773 13004
rect 25282 13001 25310 13047
rect 9761 12973 25310 13001
rect 9761 12970 9773 12973
rect 9715 12964 9773 12970
rect 25936 12961 25942 13013
rect 25994 13001 26000 13013
rect 29875 13004 29933 13010
rect 29875 13001 29887 13004
rect 25994 12973 29887 13001
rect 25994 12961 26000 12973
rect 29875 12970 29887 12973
rect 29921 12970 29933 13004
rect 33106 13001 33134 13047
rect 37426 13001 37454 13121
rect 44080 13109 44086 13121
rect 44138 13109 44144 13161
rect 41872 13035 41878 13087
rect 41930 13075 41936 13087
rect 45616 13075 45622 13087
rect 41930 13047 45622 13075
rect 41930 13035 41936 13047
rect 45616 13035 45622 13047
rect 45674 13035 45680 13087
rect 33106 12973 37454 13001
rect 29875 12964 29933 12970
rect 41008 12961 41014 13013
rect 41066 13001 41072 13013
rect 42928 13001 42934 13013
rect 41066 12973 42934 13001
rect 41066 12961 41072 12973
rect 42928 12961 42934 12973
rect 42986 12961 42992 13013
rect 49363 13004 49421 13010
rect 49363 12970 49375 13004
rect 49409 13001 49421 13004
rect 50128 13001 50134 13013
rect 49409 12973 50134 13001
rect 49409 12970 49421 12973
rect 49363 12964 49421 12970
rect 50128 12961 50134 12973
rect 50186 12961 50192 13013
rect 23440 12887 23446 12939
rect 23498 12927 23504 12939
rect 45520 12927 45526 12939
rect 23498 12899 45526 12927
rect 23498 12887 23504 12899
rect 45520 12887 45526 12899
rect 45578 12887 45584 12939
rect 1152 12680 58848 12702
rect 1152 12628 19654 12680
rect 19706 12628 19718 12680
rect 19770 12628 19782 12680
rect 19834 12628 19846 12680
rect 19898 12628 50374 12680
rect 50426 12628 50438 12680
rect 50490 12628 50502 12680
rect 50554 12628 50566 12680
rect 50618 12628 58848 12680
rect 1152 12606 58848 12628
rect 57136 12517 57142 12569
rect 57194 12557 57200 12569
rect 57331 12560 57389 12566
rect 57331 12557 57343 12560
rect 57194 12529 57343 12557
rect 57194 12517 57200 12529
rect 57331 12526 57343 12529
rect 57377 12526 57389 12560
rect 57331 12520 57389 12526
rect 13936 12443 13942 12495
rect 13994 12483 14000 12495
rect 21811 12486 21869 12492
rect 21811 12483 21823 12486
rect 13994 12455 21823 12483
rect 13994 12443 14000 12455
rect 21811 12452 21823 12455
rect 21857 12452 21869 12486
rect 21811 12446 21869 12452
rect 6064 12369 6070 12421
rect 6122 12409 6128 12421
rect 29296 12409 29302 12421
rect 6122 12381 29302 12409
rect 6122 12369 6128 12381
rect 29296 12369 29302 12381
rect 29354 12369 29360 12421
rect 57346 12409 57374 12520
rect 57619 12412 57677 12418
rect 57619 12409 57631 12412
rect 57346 12381 57631 12409
rect 57619 12378 57631 12381
rect 57665 12378 57677 12412
rect 57619 12372 57677 12378
rect 6256 12295 6262 12347
rect 6314 12335 6320 12347
rect 56176 12335 56182 12347
rect 6314 12307 56182 12335
rect 6314 12295 6320 12307
rect 56176 12295 56182 12307
rect 56234 12295 56240 12347
rect 20755 12264 20813 12270
rect 20755 12230 20767 12264
rect 20801 12261 20813 12264
rect 21043 12264 21101 12270
rect 21043 12261 21055 12264
rect 20801 12233 21055 12261
rect 20801 12230 20813 12233
rect 20755 12224 20813 12230
rect 21043 12230 21055 12233
rect 21089 12261 21101 12264
rect 21811 12264 21869 12270
rect 21089 12233 21374 12261
rect 21089 12230 21101 12233
rect 21043 12224 21101 12230
rect 21346 12187 21374 12233
rect 21811 12230 21823 12264
rect 21857 12261 21869 12264
rect 29779 12264 29837 12270
rect 29779 12261 29791 12264
rect 21857 12233 29791 12261
rect 21857 12230 21869 12233
rect 21811 12224 21869 12230
rect 29779 12230 29791 12233
rect 29825 12230 29837 12264
rect 29779 12224 29837 12230
rect 57715 12264 57773 12270
rect 57715 12230 57727 12264
rect 57761 12230 57773 12264
rect 57715 12224 57773 12230
rect 12946 12159 21182 12187
rect 21346 12159 33134 12187
rect 9619 12116 9677 12122
rect 9619 12082 9631 12116
rect 9665 12113 9677 12116
rect 9907 12116 9965 12122
rect 9907 12113 9919 12116
rect 9665 12085 9919 12113
rect 9665 12082 9677 12085
rect 9619 12076 9677 12082
rect 9907 12082 9919 12085
rect 9953 12113 9965 12116
rect 12946 12113 12974 12159
rect 9953 12085 12974 12113
rect 21154 12113 21182 12159
rect 29584 12113 29590 12125
rect 21154 12085 29590 12113
rect 9953 12082 9965 12085
rect 9907 12076 9965 12082
rect 29584 12073 29590 12085
rect 29642 12073 29648 12125
rect 33106 12113 33134 12159
rect 42640 12147 42646 12199
rect 42698 12187 42704 12199
rect 51568 12187 51574 12199
rect 42698 12159 51574 12187
rect 42698 12147 42704 12159
rect 51568 12147 51574 12159
rect 51626 12147 51632 12199
rect 57520 12147 57526 12199
rect 57578 12187 57584 12199
rect 57730 12187 57758 12224
rect 57578 12159 57758 12187
rect 57578 12147 57584 12159
rect 50224 12113 50230 12125
rect 33106 12085 50230 12113
rect 50224 12073 50230 12085
rect 50282 12073 50288 12125
rect 1152 12014 58848 12036
rect 1152 11962 4294 12014
rect 4346 11962 4358 12014
rect 4410 11962 4422 12014
rect 4474 11962 4486 12014
rect 4538 11962 35014 12014
rect 35066 11962 35078 12014
rect 35130 11962 35142 12014
rect 35194 11962 35206 12014
rect 35258 11962 58848 12014
rect 1152 11940 58848 11962
rect 7696 11851 7702 11903
rect 7754 11891 7760 11903
rect 39859 11894 39917 11900
rect 39859 11891 39871 11894
rect 7754 11863 39871 11891
rect 7754 11851 7760 11863
rect 39859 11860 39871 11863
rect 39905 11891 39917 11894
rect 40051 11894 40109 11900
rect 40051 11891 40063 11894
rect 39905 11863 40063 11891
rect 39905 11860 39917 11863
rect 39859 11854 39917 11860
rect 40051 11860 40063 11863
rect 40097 11860 40109 11894
rect 56176 11891 56182 11903
rect 56137 11863 56182 11891
rect 40051 11854 40109 11860
rect 56176 11851 56182 11863
rect 56234 11891 56240 11903
rect 56234 11863 56510 11891
rect 56234 11851 56240 11863
rect 22675 11820 22733 11826
rect 22675 11786 22687 11820
rect 22721 11817 22733 11820
rect 23440 11817 23446 11829
rect 22721 11789 23446 11817
rect 22721 11786 22733 11789
rect 22675 11780 22733 11786
rect 23440 11777 23446 11789
rect 23498 11777 23504 11829
rect 29296 11817 29302 11829
rect 29257 11789 29302 11817
rect 29296 11777 29302 11789
rect 29354 11777 29360 11829
rect 23536 11703 23542 11755
rect 23594 11743 23600 11755
rect 43024 11743 43030 11755
rect 23594 11715 43030 11743
rect 23594 11703 23600 11715
rect 43024 11703 43030 11715
rect 43082 11703 43088 11755
rect 56482 11752 56510 11863
rect 58192 11817 58198 11829
rect 57586 11789 58198 11817
rect 56467 11746 56525 11752
rect 56467 11712 56479 11746
rect 56513 11712 56525 11746
rect 56467 11706 56525 11712
rect 56563 11746 56621 11752
rect 56563 11712 56575 11746
rect 56609 11743 56621 11746
rect 57586 11743 57614 11789
rect 58192 11777 58198 11789
rect 58250 11777 58256 11829
rect 56609 11715 57614 11743
rect 56609 11712 56621 11715
rect 56563 11706 56621 11712
rect 39475 11672 39533 11678
rect 39475 11638 39487 11672
rect 39521 11669 39533 11672
rect 48112 11669 48118 11681
rect 39521 11641 48118 11669
rect 39521 11638 39533 11641
rect 39475 11632 39533 11638
rect 48112 11629 48118 11641
rect 48170 11629 48176 11681
rect 55312 11629 55318 11681
rect 55370 11669 55376 11681
rect 56947 11672 57005 11678
rect 56947 11669 56959 11672
rect 55370 11641 56959 11669
rect 55370 11629 55376 11641
rect 56947 11638 56959 11641
rect 56993 11669 57005 11672
rect 57235 11672 57293 11678
rect 57235 11669 57247 11672
rect 56993 11641 57247 11669
rect 56993 11638 57005 11641
rect 56947 11632 57005 11638
rect 57235 11638 57247 11641
rect 57281 11638 57293 11672
rect 57235 11632 57293 11638
rect 14608 11595 14614 11607
rect 14569 11567 14614 11595
rect 14608 11555 14614 11567
rect 14666 11555 14672 11607
rect 56848 11555 56854 11607
rect 56906 11595 56912 11607
rect 57315 11598 57373 11604
rect 57315 11595 57327 11598
rect 56906 11567 57327 11595
rect 56906 11555 56912 11567
rect 57315 11564 57327 11567
rect 57361 11564 57373 11598
rect 57315 11558 57373 11564
rect 23248 11481 23254 11533
rect 23306 11481 23312 11533
rect 1152 11348 58848 11370
rect 1152 11296 19654 11348
rect 19706 11296 19718 11348
rect 19770 11296 19782 11348
rect 19834 11296 19846 11348
rect 19898 11296 50374 11348
rect 50426 11296 50438 11348
rect 50490 11296 50502 11348
rect 50554 11296 50566 11348
rect 50618 11296 58848 11348
rect 1152 11274 58848 11296
rect 21520 11185 21526 11237
rect 21578 11225 21584 11237
rect 25360 11225 25366 11237
rect 21578 11197 25366 11225
rect 21578 11185 21584 11197
rect 25360 11185 25366 11197
rect 25418 11185 25424 11237
rect 31123 11228 31181 11234
rect 31123 11194 31135 11228
rect 31169 11225 31181 11228
rect 31411 11228 31469 11234
rect 31411 11225 31423 11228
rect 31169 11197 31423 11225
rect 31169 11194 31181 11197
rect 31123 11188 31181 11194
rect 31411 11194 31423 11197
rect 31457 11225 31469 11228
rect 43408 11225 43414 11237
rect 31457 11197 43414 11225
rect 31457 11194 31469 11197
rect 31411 11188 31469 11194
rect 43408 11185 43414 11197
rect 43466 11185 43472 11237
rect 13840 11111 13846 11163
rect 13898 11151 13904 11163
rect 25168 11151 25174 11163
rect 13898 11123 25174 11151
rect 13898 11111 13904 11123
rect 25168 11111 25174 11123
rect 25226 11111 25232 11163
rect 23920 11037 23926 11089
rect 23978 11077 23984 11089
rect 37456 11077 37462 11089
rect 23978 11049 37462 11077
rect 23978 11037 23984 11049
rect 37456 11037 37462 11049
rect 37514 11037 37520 11089
rect 57331 11080 57389 11086
rect 57331 11077 57343 11080
rect 43186 11049 57343 11077
rect 17584 10963 17590 11015
rect 17642 11003 17648 11015
rect 38320 11003 38326 11015
rect 17642 10975 38326 11003
rect 17642 10963 17648 10975
rect 38320 10963 38326 10975
rect 38378 10963 38384 11015
rect 38512 10963 38518 11015
rect 38570 11003 38576 11015
rect 43186 11003 43214 11049
rect 57331 11046 57343 11049
rect 57377 11046 57389 11080
rect 57331 11040 57389 11046
rect 56083 11006 56141 11012
rect 56083 11003 56095 11006
rect 38570 10975 43214 11003
rect 53266 10975 56095 11003
rect 38570 10963 38576 10975
rect 4048 10889 4054 10941
rect 4106 10929 4112 10941
rect 23248 10929 23254 10941
rect 4106 10901 23254 10929
rect 4106 10889 4112 10901
rect 23248 10889 23254 10901
rect 23306 10889 23312 10941
rect 36688 10889 36694 10941
rect 36746 10929 36752 10941
rect 53266 10929 53294 10975
rect 56083 10972 56095 10975
rect 56129 10972 56141 11006
rect 56083 10966 56141 10972
rect 36746 10901 53294 10929
rect 55987 10932 56045 10938
rect 36746 10889 36752 10901
rect 55987 10898 55999 10932
rect 56033 10898 56045 10932
rect 55987 10892 56045 10898
rect 17776 10815 17782 10867
rect 17834 10855 17840 10867
rect 38224 10855 38230 10867
rect 17834 10827 38230 10855
rect 17834 10815 17840 10827
rect 38224 10815 38230 10827
rect 38282 10815 38288 10867
rect 56002 10855 56030 10892
rect 56368 10889 56374 10941
rect 56426 10929 56432 10941
rect 57235 10932 57293 10938
rect 57235 10929 57247 10932
rect 56426 10901 57247 10929
rect 56426 10889 56432 10901
rect 57235 10898 57247 10901
rect 57281 10898 57293 10932
rect 57235 10892 57293 10898
rect 57136 10855 57142 10867
rect 56002 10827 57142 10855
rect 57136 10815 57142 10827
rect 57194 10815 57200 10867
rect 6928 10781 6934 10793
rect 6889 10753 6934 10781
rect 6928 10741 6934 10753
rect 6986 10741 6992 10793
rect 15667 10784 15725 10790
rect 15667 10750 15679 10784
rect 15713 10781 15725 10784
rect 32080 10781 32086 10793
rect 15713 10753 32086 10781
rect 15713 10750 15725 10753
rect 15667 10744 15725 10750
rect 32080 10741 32086 10753
rect 32138 10741 32144 10793
rect 41104 10741 41110 10793
rect 41162 10781 41168 10793
rect 42643 10784 42701 10790
rect 42643 10781 42655 10784
rect 41162 10753 42655 10781
rect 41162 10741 41168 10753
rect 42643 10750 42655 10753
rect 42689 10750 42701 10784
rect 54352 10781 54358 10793
rect 54313 10753 54358 10781
rect 42643 10744 42701 10750
rect 54352 10741 54358 10753
rect 54410 10741 54416 10793
rect 1152 10682 58848 10704
rect 1152 10630 4294 10682
rect 4346 10630 4358 10682
rect 4410 10630 4422 10682
rect 4474 10630 4486 10682
rect 4538 10630 35014 10682
rect 35066 10630 35078 10682
rect 35130 10630 35142 10682
rect 35194 10630 35206 10682
rect 35258 10630 58848 10682
rect 1152 10608 58848 10630
rect 56272 10559 56278 10571
rect 56233 10531 56278 10559
rect 56272 10519 56278 10531
rect 56330 10519 56336 10571
rect 6928 10445 6934 10497
rect 6986 10485 6992 10497
rect 16144 10485 16150 10497
rect 6986 10457 16150 10485
rect 6986 10445 6992 10457
rect 16144 10445 16150 10457
rect 16202 10445 16208 10497
rect 23155 10488 23213 10494
rect 23155 10454 23167 10488
rect 23201 10485 23213 10488
rect 31504 10485 31510 10497
rect 23201 10457 31510 10485
rect 23201 10454 23213 10457
rect 23155 10448 23213 10454
rect 31504 10445 31510 10457
rect 31562 10445 31568 10497
rect 14224 10371 14230 10423
rect 14282 10411 14288 10423
rect 25264 10411 25270 10423
rect 14282 10383 25270 10411
rect 14282 10371 14288 10383
rect 25264 10371 25270 10383
rect 25322 10371 25328 10423
rect 35344 10371 35350 10423
rect 35402 10411 35408 10423
rect 36976 10411 36982 10423
rect 35402 10383 36982 10411
rect 35402 10371 35408 10383
rect 36976 10371 36982 10383
rect 37034 10371 37040 10423
rect 54835 10414 54893 10420
rect 54835 10380 54847 10414
rect 54881 10411 54893 10414
rect 55024 10411 55030 10423
rect 54881 10383 55030 10411
rect 54881 10380 54893 10383
rect 54835 10374 54893 10380
rect 55024 10371 55030 10383
rect 55082 10411 55088 10423
rect 55315 10414 55373 10420
rect 55315 10411 55327 10414
rect 55082 10383 55327 10411
rect 55082 10371 55088 10383
rect 55315 10380 55327 10383
rect 55361 10380 55373 10414
rect 55315 10374 55373 10380
rect 55891 10414 55949 10420
rect 55891 10380 55903 10414
rect 55937 10411 55949 10414
rect 55984 10411 55990 10423
rect 55937 10383 55990 10411
rect 55937 10380 55949 10383
rect 55891 10374 55949 10380
rect 55984 10371 55990 10383
rect 56042 10371 56048 10423
rect 56290 10411 56318 10519
rect 56563 10414 56621 10420
rect 56563 10411 56575 10414
rect 56290 10383 56575 10411
rect 56563 10380 56575 10383
rect 56609 10380 56621 10414
rect 57424 10411 57430 10423
rect 57385 10383 57430 10411
rect 56563 10374 56621 10380
rect 57424 10371 57430 10383
rect 57482 10371 57488 10423
rect 20656 10297 20662 10349
rect 20714 10337 20720 10349
rect 31216 10337 31222 10349
rect 20714 10309 31222 10337
rect 20714 10297 20720 10309
rect 31216 10297 31222 10309
rect 31274 10297 31280 10349
rect 52912 10337 52918 10349
rect 33106 10309 52918 10337
rect 12595 10266 12653 10272
rect 12595 10232 12607 10266
rect 12641 10263 12653 10266
rect 33106 10263 33134 10309
rect 52912 10297 52918 10309
rect 52970 10297 52976 10349
rect 12641 10235 33134 10263
rect 38803 10266 38861 10272
rect 12641 10232 12653 10235
rect 12595 10226 12653 10232
rect 38803 10232 38815 10266
rect 38849 10263 38861 10266
rect 47824 10263 47830 10275
rect 38849 10235 47830 10263
rect 38849 10232 38861 10235
rect 38803 10226 38861 10232
rect 47824 10223 47830 10235
rect 47882 10223 47888 10275
rect 17296 10149 17302 10201
rect 17354 10189 17360 10201
rect 23155 10192 23213 10198
rect 23155 10189 23167 10192
rect 17354 10161 23167 10189
rect 17354 10149 17360 10161
rect 23155 10158 23167 10161
rect 23201 10158 23213 10192
rect 31120 10189 31126 10201
rect 23155 10152 23213 10158
rect 23362 10161 31126 10189
rect 10768 10075 10774 10127
rect 10826 10115 10832 10127
rect 12976 10115 12982 10127
rect 10826 10087 12982 10115
rect 10826 10075 10832 10087
rect 12976 10075 12982 10087
rect 13034 10075 13040 10127
rect 18448 10075 18454 10127
rect 18506 10115 18512 10127
rect 19408 10115 19414 10127
rect 18506 10087 19414 10115
rect 18506 10075 18512 10087
rect 19408 10075 19414 10087
rect 19466 10075 19472 10127
rect 21040 10075 21046 10127
rect 21098 10115 21104 10127
rect 23362 10115 23390 10161
rect 31120 10149 31126 10161
rect 31178 10149 31184 10201
rect 58576 10189 58582 10201
rect 55138 10161 58582 10189
rect 21098 10087 23390 10115
rect 21098 10075 21104 10087
rect 23440 10075 23446 10127
rect 23498 10115 23504 10127
rect 25552 10115 25558 10127
rect 23498 10087 25558 10115
rect 23498 10075 23504 10087
rect 25552 10075 25558 10087
rect 25610 10075 25616 10127
rect 45328 10075 45334 10127
rect 45386 10115 45392 10127
rect 47152 10115 47158 10127
rect 45386 10087 47158 10115
rect 45386 10075 45392 10087
rect 47152 10075 47158 10087
rect 47210 10075 47216 10127
rect 49648 10075 49654 10127
rect 49706 10115 49712 10127
rect 50704 10115 50710 10127
rect 49706 10087 50710 10115
rect 49706 10075 49712 10087
rect 50704 10075 50710 10087
rect 50762 10075 50768 10127
rect 55138 10124 55166 10161
rect 58576 10149 58582 10161
rect 58634 10149 58640 10201
rect 55123 10118 55181 10124
rect 55123 10084 55135 10118
rect 55169 10084 55181 10118
rect 55123 10078 55181 10084
rect 55696 10075 55702 10127
rect 55754 10115 55760 10127
rect 55795 10118 55853 10124
rect 55795 10115 55807 10118
rect 55754 10087 55807 10115
rect 55754 10075 55760 10087
rect 55795 10084 55807 10087
rect 55841 10084 55853 10118
rect 55795 10078 55853 10084
rect 56080 10075 56086 10127
rect 56138 10115 56144 10127
rect 56659 10118 56717 10124
rect 56659 10115 56671 10118
rect 56138 10087 56671 10115
rect 56138 10075 56144 10087
rect 56659 10084 56671 10087
rect 56705 10084 56717 10118
rect 56659 10078 56717 10084
rect 56752 10075 56758 10127
rect 56810 10115 56816 10127
rect 57331 10118 57389 10124
rect 57331 10115 57343 10118
rect 56810 10087 57343 10115
rect 56810 10075 56816 10087
rect 57331 10084 57343 10087
rect 57377 10084 57389 10118
rect 57331 10078 57389 10084
rect 1152 10016 58848 10038
rect 1152 9964 19654 10016
rect 19706 9964 19718 10016
rect 19770 9964 19782 10016
rect 19834 9964 19846 10016
rect 19898 9964 50374 10016
rect 50426 9964 50438 10016
rect 50490 9964 50502 10016
rect 50554 9964 50566 10016
rect 50618 9964 58848 10016
rect 1152 9942 58848 9964
rect 12403 9896 12461 9902
rect 12403 9862 12415 9896
rect 12449 9893 12461 9896
rect 48592 9893 48598 9905
rect 12449 9865 48598 9893
rect 12449 9862 12461 9865
rect 12403 9856 12461 9862
rect 48592 9853 48598 9865
rect 48650 9853 48656 9905
rect 14608 9779 14614 9831
rect 14666 9819 14672 9831
rect 54160 9819 54166 9831
rect 14666 9791 54166 9819
rect 14666 9779 14672 9791
rect 54160 9779 54166 9791
rect 54218 9779 54224 9831
rect 5488 9705 5494 9757
rect 5546 9705 5552 9757
rect 16816 9705 16822 9757
rect 16874 9745 16880 9757
rect 26227 9748 26285 9754
rect 26227 9745 26239 9748
rect 16874 9717 26239 9745
rect 16874 9705 16880 9717
rect 26227 9714 26239 9717
rect 26273 9745 26285 9748
rect 26419 9748 26477 9754
rect 26419 9745 26431 9748
rect 26273 9717 26431 9745
rect 26273 9714 26285 9717
rect 26227 9708 26285 9714
rect 26419 9714 26431 9717
rect 26465 9714 26477 9748
rect 26419 9708 26477 9714
rect 28144 9705 28150 9757
rect 28202 9745 28208 9757
rect 28528 9745 28534 9757
rect 28202 9717 28534 9745
rect 28202 9705 28208 9717
rect 28528 9705 28534 9717
rect 28586 9705 28592 9757
rect 32656 9705 32662 9757
rect 32714 9745 32720 9757
rect 54835 9748 54893 9754
rect 54835 9745 54847 9748
rect 32714 9717 54847 9745
rect 32714 9705 32720 9717
rect 54835 9714 54847 9717
rect 54881 9745 54893 9748
rect 55123 9748 55181 9754
rect 55123 9745 55135 9748
rect 54881 9717 55135 9745
rect 54881 9714 54893 9717
rect 54835 9708 54893 9714
rect 55123 9714 55135 9717
rect 55169 9714 55181 9748
rect 55123 9708 55181 9714
rect 55699 9748 55757 9754
rect 55699 9714 55711 9748
rect 55745 9745 55757 9748
rect 55888 9745 55894 9757
rect 55745 9717 55894 9745
rect 55745 9714 55757 9717
rect 55699 9708 55757 9714
rect 55888 9705 55894 9717
rect 55946 9745 55952 9757
rect 56179 9748 56237 9754
rect 56179 9745 56191 9748
rect 55946 9717 56191 9745
rect 55946 9705 55952 9717
rect 56179 9714 56191 9717
rect 56225 9714 56237 9748
rect 56179 9708 56237 9714
rect 5506 9620 5534 9705
rect 39664 9671 39670 9683
rect 12946 9643 39670 9671
rect 12946 9597 12974 9643
rect 39664 9631 39670 9643
rect 39722 9631 39728 9683
rect 57616 9631 57622 9683
rect 57674 9671 57680 9683
rect 57674 9643 57719 9671
rect 57674 9631 57680 9643
rect 42544 9597 42550 9609
rect 9888 9569 12974 9597
rect 23026 9569 42550 9597
rect 4435 9526 4493 9532
rect 4435 9492 4447 9526
rect 4481 9523 4493 9526
rect 23026 9523 23054 9569
rect 42544 9557 42550 9569
rect 42602 9557 42608 9609
rect 54256 9557 54262 9609
rect 54314 9597 54320 9609
rect 54355 9600 54413 9606
rect 54355 9597 54367 9600
rect 54314 9569 54367 9597
rect 54314 9557 54320 9569
rect 54355 9566 54367 9569
rect 54401 9566 54413 9600
rect 54355 9560 54413 9566
rect 54451 9600 54509 9606
rect 54451 9566 54463 9600
rect 54497 9597 54509 9600
rect 54832 9597 54838 9609
rect 54497 9569 54838 9597
rect 54497 9566 54509 9569
rect 54451 9560 54509 9566
rect 54832 9557 54838 9569
rect 54890 9557 54896 9609
rect 55219 9600 55277 9606
rect 55219 9566 55231 9600
rect 55265 9566 55277 9600
rect 55219 9560 55277 9566
rect 55987 9600 56045 9606
rect 55987 9566 55999 9600
rect 56033 9566 56045 9600
rect 55987 9560 56045 9566
rect 53395 9526 53453 9532
rect 53395 9523 53407 9526
rect 4481 9495 7214 9523
rect 9744 9495 23054 9523
rect 25666 9495 53407 9523
rect 4481 9492 4493 9495
rect 4435 9486 4493 9492
rect 7186 9449 7214 9495
rect 12403 9452 12461 9458
rect 12403 9449 12415 9452
rect 7186 9421 12415 9449
rect 12403 9418 12415 9421
rect 12449 9418 12461 9452
rect 12403 9412 12461 9418
rect 12496 9409 12502 9461
rect 12554 9449 12560 9461
rect 25666 9449 25694 9495
rect 53395 9492 53407 9495
rect 53441 9523 53453 9526
rect 53587 9526 53645 9532
rect 53587 9523 53599 9526
rect 53441 9495 53599 9523
rect 53441 9492 53453 9495
rect 53395 9486 53453 9492
rect 53587 9492 53599 9495
rect 53633 9492 53645 9526
rect 53587 9486 53645 9492
rect 55024 9483 55030 9535
rect 55082 9523 55088 9535
rect 55234 9523 55262 9560
rect 55082 9495 55262 9523
rect 55082 9483 55088 9495
rect 55312 9483 55318 9535
rect 55370 9523 55376 9535
rect 56002 9523 56030 9560
rect 55370 9495 56030 9523
rect 55370 9483 55376 9495
rect 45616 9449 45622 9461
rect 12554 9421 25694 9449
rect 45577 9421 45622 9449
rect 12554 9409 12560 9421
rect 45616 9409 45622 9421
rect 45674 9409 45680 9461
rect 46768 9449 46774 9461
rect 46729 9421 46774 9449
rect 46768 9409 46774 9421
rect 46826 9409 46832 9461
rect 1152 9350 58848 9372
rect 1152 9298 4294 9350
rect 4346 9298 4358 9350
rect 4410 9298 4422 9350
rect 4474 9298 4486 9350
rect 4538 9298 35014 9350
rect 35066 9298 35078 9350
rect 35130 9298 35142 9350
rect 35194 9298 35206 9350
rect 35258 9298 58848 9350
rect 1152 9276 58848 9298
rect 28240 9187 28246 9239
rect 28298 9227 28304 9239
rect 46768 9227 46774 9239
rect 28298 9199 46774 9227
rect 28298 9187 28304 9199
rect 46768 9187 46774 9199
rect 46826 9187 46832 9239
rect 54160 9187 54166 9239
rect 54218 9227 54224 9239
rect 54259 9230 54317 9236
rect 54259 9227 54271 9230
rect 54218 9199 54271 9227
rect 54218 9187 54224 9199
rect 54259 9196 54271 9199
rect 54305 9196 54317 9230
rect 54259 9190 54317 9196
rect 5488 9113 5494 9165
rect 5546 9153 5552 9165
rect 46096 9153 46102 9165
rect 5546 9125 46102 9153
rect 5546 9113 5552 9125
rect 46096 9113 46102 9125
rect 46154 9113 46160 9165
rect 55984 9153 55990 9165
rect 53410 9125 55990 9153
rect 12304 9039 12310 9091
rect 12362 9079 12368 9091
rect 38803 9082 38861 9088
rect 38803 9079 38815 9082
rect 12362 9051 38815 9079
rect 12362 9039 12368 9051
rect 38803 9048 38815 9051
rect 38849 9048 38861 9082
rect 53104 9079 53110 9091
rect 53017 9051 53110 9079
rect 38803 9042 38861 9048
rect 53104 9039 53110 9051
rect 53162 9079 53168 9091
rect 53410 9088 53438 9125
rect 55984 9113 55990 9125
rect 56042 9113 56048 9165
rect 53299 9082 53357 9088
rect 53299 9079 53311 9082
rect 53162 9051 53311 9079
rect 53162 9039 53168 9051
rect 53299 9048 53311 9051
rect 53345 9048 53357 9082
rect 53299 9042 53357 9048
rect 53395 9082 53453 9088
rect 53395 9048 53407 9082
rect 53441 9048 53453 9082
rect 53395 9042 53453 9048
rect 53872 9039 53878 9091
rect 53930 9079 53936 9091
rect 54643 9082 54701 9088
rect 54643 9079 54655 9082
rect 53930 9051 54655 9079
rect 53930 9039 53936 9051
rect 54643 9048 54655 9051
rect 54689 9048 54701 9082
rect 54643 9042 54701 9048
rect 20464 8965 20470 9017
rect 20522 9005 20528 9017
rect 55027 9008 55085 9014
rect 55027 9005 55039 9008
rect 20522 8977 55039 9005
rect 20522 8965 20528 8977
rect 55027 8974 55039 8977
rect 55073 9005 55085 9008
rect 55315 9008 55373 9014
rect 55315 9005 55327 9008
rect 55073 8977 55327 9005
rect 55073 8974 55085 8977
rect 55027 8968 55085 8974
rect 55315 8974 55327 8977
rect 55361 8974 55373 9008
rect 56560 9005 56566 9017
rect 56521 8977 56566 9005
rect 55315 8968 55373 8974
rect 56560 8965 56566 8977
rect 56618 8965 56624 9017
rect 57232 9005 57238 9017
rect 57193 8977 57238 9005
rect 57232 8965 57238 8977
rect 57290 8965 57296 9017
rect 1747 8934 1805 8940
rect 1747 8900 1759 8934
rect 1793 8900 1805 8934
rect 1747 8894 1805 8900
rect 3475 8934 3533 8940
rect 3475 8900 3487 8934
rect 3521 8931 3533 8934
rect 14704 8931 14710 8943
rect 3521 8903 14710 8931
rect 3521 8900 3533 8903
rect 3475 8894 3533 8900
rect 1762 8857 1790 8894
rect 14704 8891 14710 8903
rect 14762 8891 14768 8943
rect 49168 8891 49174 8943
rect 49226 8931 49232 8943
rect 52723 8934 52781 8940
rect 52723 8931 52735 8934
rect 49226 8903 52735 8931
rect 49226 8891 49232 8903
rect 52723 8900 52735 8903
rect 52769 8900 52781 8934
rect 52723 8894 52781 8900
rect 54160 8891 54166 8943
rect 54218 8931 54224 8943
rect 54547 8934 54605 8940
rect 54547 8931 54559 8934
rect 54218 8903 54559 8931
rect 54218 8891 54224 8903
rect 54547 8900 54559 8903
rect 54593 8900 54605 8934
rect 54547 8894 54605 8900
rect 56368 8891 56374 8943
rect 56426 8931 56432 8943
rect 56848 8931 56854 8943
rect 56426 8903 56854 8931
rect 56426 8891 56432 8903
rect 56848 8891 56854 8903
rect 56906 8891 56912 8943
rect 36688 8857 36694 8869
rect 1762 8829 36694 8857
rect 36688 8817 36694 8829
rect 36746 8817 36752 8869
rect 54562 8829 55454 8857
rect 54562 8795 54590 8829
rect 10963 8786 11021 8792
rect 10963 8752 10975 8786
rect 11009 8783 11021 8786
rect 11251 8786 11309 8792
rect 11251 8783 11263 8786
rect 11009 8755 11263 8783
rect 11009 8752 11021 8755
rect 10963 8746 11021 8752
rect 11251 8752 11263 8755
rect 11297 8783 11309 8786
rect 51664 8783 51670 8795
rect 11297 8755 51670 8783
rect 11297 8752 11309 8755
rect 11251 8746 11309 8752
rect 51664 8743 51670 8755
rect 51722 8743 51728 8795
rect 54544 8743 54550 8795
rect 54602 8743 54608 8795
rect 55426 8792 55454 8829
rect 55411 8786 55469 8792
rect 55411 8752 55423 8786
rect 55457 8752 55469 8786
rect 55411 8746 55469 8752
rect 1152 8684 58848 8706
rect 1152 8632 19654 8684
rect 19706 8632 19718 8684
rect 19770 8632 19782 8684
rect 19834 8632 19846 8684
rect 19898 8632 50374 8684
rect 50426 8632 50438 8684
rect 50490 8632 50502 8684
rect 50554 8632 50566 8684
rect 50618 8632 58848 8684
rect 1152 8610 58848 8632
rect 2128 8561 2134 8573
rect 2089 8533 2134 8561
rect 2128 8521 2134 8533
rect 2186 8521 2192 8573
rect 39091 8564 39149 8570
rect 39091 8530 39103 8564
rect 39137 8561 39149 8564
rect 39184 8561 39190 8573
rect 39137 8533 39190 8561
rect 39137 8530 39149 8533
rect 39091 8524 39149 8530
rect 39184 8521 39190 8533
rect 39242 8521 39248 8573
rect 42256 8561 42262 8573
rect 42217 8533 42262 8561
rect 42256 8521 42262 8533
rect 42314 8521 42320 8573
rect 44080 8561 44086 8573
rect 44041 8533 44086 8561
rect 44080 8521 44086 8533
rect 44138 8521 44144 8573
rect 48208 8561 48214 8573
rect 48169 8533 48214 8561
rect 48208 8521 48214 8533
rect 48266 8561 48272 8573
rect 52243 8564 52301 8570
rect 48266 8533 48542 8561
rect 48266 8521 48272 8533
rect 2146 8413 2174 8521
rect 2515 8416 2573 8422
rect 2515 8413 2527 8416
rect 2146 8385 2527 8413
rect 2515 8382 2527 8385
rect 2561 8382 2573 8416
rect 2515 8376 2573 8382
rect 4243 8416 4301 8422
rect 4243 8382 4255 8416
rect 4289 8413 4301 8416
rect 4531 8416 4589 8422
rect 4531 8413 4543 8416
rect 4289 8385 4543 8413
rect 4289 8382 4301 8385
rect 4243 8376 4301 8382
rect 4531 8382 4543 8385
rect 4577 8413 4589 8416
rect 9328 8413 9334 8425
rect 4577 8385 9334 8413
rect 4577 8382 4589 8385
rect 4531 8376 4589 8382
rect 9328 8373 9334 8385
rect 9386 8373 9392 8425
rect 10768 8413 10774 8425
rect 10729 8385 10774 8413
rect 10768 8373 10774 8385
rect 10826 8373 10832 8425
rect 11251 8416 11309 8422
rect 11251 8382 11263 8416
rect 11297 8413 11309 8416
rect 11536 8413 11542 8425
rect 11297 8385 11542 8413
rect 11297 8382 11309 8385
rect 11251 8376 11309 8382
rect 11536 8373 11542 8385
rect 11594 8373 11600 8425
rect 12304 8413 12310 8425
rect 12265 8385 12310 8413
rect 12304 8373 12310 8385
rect 12362 8373 12368 8425
rect 16144 8373 16150 8425
rect 16202 8413 16208 8425
rect 16243 8416 16301 8422
rect 16243 8413 16255 8416
rect 16202 8385 16255 8413
rect 16202 8373 16208 8385
rect 16243 8382 16255 8385
rect 16289 8382 16301 8416
rect 16243 8376 16301 8382
rect 16723 8416 16781 8422
rect 16723 8382 16735 8416
rect 16769 8413 16781 8416
rect 17008 8413 17014 8425
rect 16769 8385 17014 8413
rect 16769 8382 16781 8385
rect 16723 8376 16781 8382
rect 17008 8373 17014 8385
rect 17066 8373 17072 8425
rect 39202 8413 39230 8521
rect 39283 8416 39341 8422
rect 39283 8413 39295 8416
rect 39202 8385 39295 8413
rect 39283 8382 39295 8385
rect 39329 8382 39341 8416
rect 42274 8413 42302 8521
rect 42547 8416 42605 8422
rect 42547 8413 42559 8416
rect 42274 8385 42559 8413
rect 39283 8376 39341 8382
rect 42547 8382 42559 8385
rect 42593 8382 42605 8416
rect 44098 8413 44126 8521
rect 44371 8416 44429 8422
rect 44371 8413 44383 8416
rect 44098 8385 44383 8413
rect 42547 8376 42605 8382
rect 44371 8382 44383 8385
rect 44417 8382 44429 8416
rect 44371 8376 44429 8382
rect 47539 8416 47597 8422
rect 47539 8382 47551 8416
rect 47585 8413 47597 8416
rect 47827 8416 47885 8422
rect 47827 8413 47839 8416
rect 47585 8385 47839 8413
rect 47585 8382 47597 8385
rect 47539 8376 47597 8382
rect 47827 8382 47839 8385
rect 47873 8413 47885 8416
rect 47920 8413 47926 8425
rect 47873 8385 47926 8413
rect 47873 8382 47885 8385
rect 47827 8376 47885 8382
rect 47920 8373 47926 8385
rect 47978 8373 47984 8425
rect 48514 8422 48542 8533
rect 52243 8530 52255 8564
rect 52289 8561 52301 8564
rect 52336 8561 52342 8573
rect 52289 8533 52342 8561
rect 52289 8530 52301 8533
rect 52243 8524 52301 8530
rect 52336 8521 52342 8533
rect 52394 8521 52400 8573
rect 52912 8561 52918 8573
rect 52873 8533 52918 8561
rect 52912 8521 52918 8533
rect 52970 8521 52976 8573
rect 48499 8416 48557 8422
rect 48499 8382 48511 8416
rect 48545 8382 48557 8416
rect 49360 8413 49366 8425
rect 49321 8385 49366 8413
rect 48499 8376 48557 8382
rect 49360 8373 49366 8385
rect 49418 8373 49424 8425
rect 50128 8413 50134 8425
rect 50089 8385 50134 8413
rect 50128 8373 50134 8385
rect 50186 8373 50192 8425
rect 52354 8413 52382 8521
rect 52435 8416 52493 8422
rect 52435 8413 52447 8416
rect 52354 8385 52447 8413
rect 52435 8382 52447 8385
rect 52481 8382 52493 8416
rect 52930 8413 52958 8521
rect 53203 8416 53261 8422
rect 53203 8413 53215 8416
rect 52930 8385 53215 8413
rect 52435 8376 52493 8382
rect 53203 8382 53215 8385
rect 53249 8382 53261 8416
rect 53203 8376 53261 8382
rect 54067 8416 54125 8422
rect 54067 8382 54079 8416
rect 54113 8413 54125 8416
rect 54352 8413 54358 8425
rect 54113 8385 54358 8413
rect 54113 8382 54125 8385
rect 54067 8376 54125 8382
rect 54352 8373 54358 8385
rect 54410 8373 54416 8425
rect 2899 8342 2957 8348
rect 2899 8308 2911 8342
rect 2945 8339 2957 8342
rect 3283 8342 3341 8348
rect 3283 8339 3295 8342
rect 2945 8311 3295 8339
rect 2945 8308 2957 8311
rect 2899 8302 2957 8308
rect 3283 8308 3295 8311
rect 3329 8339 3341 8342
rect 21328 8339 21334 8351
rect 3329 8311 21334 8339
rect 3329 8308 3341 8311
rect 3283 8302 3341 8308
rect 21328 8299 21334 8311
rect 21386 8299 21392 8351
rect 53104 8299 53110 8351
rect 53162 8339 53168 8351
rect 55219 8342 55277 8348
rect 53162 8311 53246 8339
rect 53162 8299 53168 8311
rect 1648 8265 1654 8277
rect 1609 8237 1654 8265
rect 1648 8225 1654 8237
rect 1706 8225 1712 8277
rect 1747 8268 1805 8274
rect 1747 8234 1759 8268
rect 1793 8234 1805 8268
rect 1747 8228 1805 8234
rect 1762 8191 1790 8228
rect 2128 8225 2134 8277
rect 2186 8265 2192 8277
rect 2419 8268 2477 8274
rect 2419 8265 2431 8268
rect 2186 8237 2431 8265
rect 2186 8225 2192 8237
rect 2419 8234 2431 8237
rect 2465 8234 2477 8268
rect 2419 8228 2477 8234
rect 2992 8225 2998 8277
rect 3050 8265 3056 8277
rect 3187 8268 3245 8274
rect 3187 8265 3199 8268
rect 3050 8237 3199 8265
rect 3050 8225 3056 8237
rect 3187 8234 3199 8237
rect 3233 8234 3245 8268
rect 3187 8228 3245 8234
rect 4435 8268 4493 8274
rect 4435 8234 4447 8268
rect 4481 8265 4493 8268
rect 4816 8265 4822 8277
rect 4481 8237 4822 8265
rect 4481 8234 4493 8237
rect 4435 8228 4493 8234
rect 4816 8225 4822 8237
rect 4874 8225 4880 8277
rect 10576 8225 10582 8277
rect 10634 8265 10640 8277
rect 10675 8268 10733 8274
rect 10675 8265 10687 8268
rect 10634 8237 10687 8265
rect 10634 8225 10640 8237
rect 10675 8234 10687 8237
rect 10721 8234 10733 8268
rect 10675 8228 10733 8234
rect 10960 8225 10966 8277
rect 11018 8265 11024 8277
rect 11443 8268 11501 8274
rect 11443 8265 11455 8268
rect 11018 8237 11455 8265
rect 11018 8225 11024 8237
rect 11443 8234 11455 8237
rect 11489 8234 11501 8268
rect 11443 8228 11501 8234
rect 11728 8225 11734 8277
rect 11786 8265 11792 8277
rect 12211 8268 12269 8274
rect 12211 8265 12223 8268
rect 11786 8237 12223 8265
rect 11786 8225 11792 8237
rect 12211 8234 12223 8237
rect 12257 8234 12269 8268
rect 12211 8228 12269 8234
rect 12496 8225 12502 8277
rect 12554 8265 12560 8277
rect 12979 8268 13037 8274
rect 12979 8265 12991 8268
rect 12554 8237 12991 8265
rect 12554 8225 12560 8237
rect 12979 8234 12991 8237
rect 13025 8234 13037 8268
rect 12979 8228 13037 8234
rect 13075 8268 13133 8274
rect 13075 8234 13087 8268
rect 13121 8234 13133 8268
rect 13075 8228 13133 8234
rect 2035 8194 2093 8200
rect 2035 8191 2047 8194
rect 1762 8163 2047 8191
rect 2035 8160 2047 8163
rect 2081 8191 2093 8194
rect 3664 8191 3670 8203
rect 2081 8163 3670 8191
rect 2081 8160 2093 8163
rect 2035 8154 2093 8160
rect 3664 8151 3670 8163
rect 3722 8151 3728 8203
rect 13090 8191 13118 8228
rect 16048 8225 16054 8277
rect 16106 8265 16112 8277
rect 16147 8268 16205 8274
rect 16147 8265 16159 8268
rect 16106 8237 16159 8265
rect 16106 8225 16112 8237
rect 16147 8234 16159 8237
rect 16193 8234 16205 8268
rect 16147 8228 16205 8234
rect 16336 8225 16342 8277
rect 16394 8265 16400 8277
rect 16915 8268 16973 8274
rect 16915 8265 16927 8268
rect 16394 8237 16927 8265
rect 16394 8225 16400 8237
rect 16915 8234 16927 8237
rect 16961 8234 16973 8268
rect 16915 8228 16973 8234
rect 39184 8225 39190 8277
rect 39242 8265 39248 8277
rect 39379 8268 39437 8274
rect 39379 8265 39391 8268
rect 39242 8237 39391 8265
rect 39242 8225 39248 8237
rect 39379 8234 39391 8237
rect 39425 8234 39437 8268
rect 39379 8228 39437 8234
rect 42352 8225 42358 8277
rect 42410 8265 42416 8277
rect 42643 8268 42701 8274
rect 42643 8265 42655 8268
rect 42410 8237 42655 8265
rect 42410 8225 42416 8237
rect 42643 8234 42655 8237
rect 42689 8234 42701 8268
rect 42643 8228 42701 8234
rect 44272 8225 44278 8277
rect 44330 8265 44336 8277
rect 44467 8268 44525 8274
rect 44467 8265 44479 8268
rect 44330 8237 44479 8265
rect 44330 8225 44336 8237
rect 44467 8234 44479 8237
rect 44513 8234 44525 8268
rect 44467 8228 44525 8234
rect 47632 8225 47638 8277
rect 47690 8265 47696 8277
rect 47731 8268 47789 8274
rect 47731 8265 47743 8268
rect 47690 8237 47743 8265
rect 47690 8225 47696 8237
rect 47731 8234 47743 8237
rect 47777 8234 47789 8268
rect 47731 8228 47789 8234
rect 48016 8225 48022 8277
rect 48074 8265 48080 8277
rect 48595 8268 48653 8274
rect 48595 8265 48607 8268
rect 48074 8237 48607 8265
rect 48074 8225 48080 8237
rect 48595 8234 48607 8237
rect 48641 8234 48653 8268
rect 48595 8228 48653 8234
rect 48688 8225 48694 8277
rect 48746 8265 48752 8277
rect 49267 8268 49325 8274
rect 49267 8265 49279 8268
rect 48746 8237 49279 8265
rect 48746 8225 48752 8237
rect 49267 8234 49279 8237
rect 49313 8234 49325 8268
rect 49267 8228 49325 8234
rect 49456 8225 49462 8277
rect 49514 8265 49520 8277
rect 50035 8268 50093 8274
rect 50035 8265 50047 8268
rect 49514 8237 50047 8265
rect 49514 8225 49520 8237
rect 50035 8234 50047 8237
rect 50081 8234 50093 8268
rect 50035 8228 50093 8234
rect 52531 8268 52589 8274
rect 52531 8234 52543 8268
rect 52577 8265 52589 8268
rect 52577 8237 53150 8265
rect 52577 8234 52589 8237
rect 52531 8228 52589 8234
rect 40147 8194 40205 8200
rect 40147 8191 40159 8194
rect 13090 8163 40159 8191
rect 40147 8160 40159 8163
rect 40193 8160 40205 8194
rect 40147 8154 40205 8160
rect 7504 8117 7510 8129
rect 7465 8089 7510 8117
rect 7504 8077 7510 8089
rect 7562 8077 7568 8129
rect 12400 8077 12406 8129
rect 12458 8117 12464 8129
rect 13744 8117 13750 8129
rect 12458 8089 13750 8117
rect 12458 8077 12464 8089
rect 13744 8077 13750 8089
rect 13802 8077 13808 8129
rect 13843 8120 13901 8126
rect 13843 8086 13855 8120
rect 13889 8117 13901 8120
rect 15760 8117 15766 8129
rect 13889 8089 15766 8117
rect 13889 8086 13901 8089
rect 13843 8080 13901 8086
rect 15760 8077 15766 8089
rect 15818 8077 15824 8129
rect 43411 8120 43469 8126
rect 43411 8086 43423 8120
rect 43457 8117 43469 8120
rect 51088 8117 51094 8129
rect 43457 8089 51094 8117
rect 43457 8086 43469 8089
rect 43411 8080 43469 8086
rect 51088 8077 51094 8089
rect 51146 8077 51152 8129
rect 53122 8117 53150 8237
rect 53218 8191 53246 8311
rect 55219 8308 55231 8342
rect 55265 8339 55277 8342
rect 55987 8342 56045 8348
rect 55265 8311 55934 8339
rect 55265 8308 55277 8311
rect 55219 8302 55277 8308
rect 53299 8268 53357 8274
rect 53299 8234 53311 8268
rect 53345 8234 53357 8268
rect 53299 8228 53357 8234
rect 53314 8191 53342 8228
rect 53488 8225 53494 8277
rect 53546 8265 53552 8277
rect 53971 8268 54029 8274
rect 53971 8265 53983 8268
rect 53546 8237 53983 8265
rect 53546 8225 53552 8237
rect 53971 8234 53983 8237
rect 54017 8234 54029 8268
rect 53971 8228 54029 8234
rect 53218 8163 53342 8191
rect 55906 8191 55934 8311
rect 55987 8308 55999 8342
rect 56033 8308 56045 8342
rect 55987 8302 56045 8308
rect 56002 8265 56030 8302
rect 56944 8299 56950 8351
rect 57002 8339 57008 8351
rect 57139 8342 57197 8348
rect 57139 8339 57151 8342
rect 57002 8311 57151 8339
rect 57002 8299 57008 8311
rect 57139 8308 57151 8311
rect 57185 8308 57197 8342
rect 57139 8302 57197 8308
rect 58384 8265 58390 8277
rect 56002 8237 58390 8265
rect 58384 8225 58390 8237
rect 58442 8225 58448 8277
rect 59824 8191 59830 8203
rect 55906 8163 59830 8191
rect 59824 8151 59830 8163
rect 59882 8151 59888 8203
rect 58960 8117 58966 8129
rect 53122 8089 58966 8117
rect 58960 8077 58966 8089
rect 59018 8077 59024 8129
rect 1152 8018 58848 8040
rect 1152 7966 4294 8018
rect 4346 7966 4358 8018
rect 4410 7966 4422 8018
rect 4474 7966 4486 8018
rect 4538 7966 35014 8018
rect 35066 7966 35078 8018
rect 35130 7966 35142 8018
rect 35194 7966 35206 8018
rect 35258 7966 58848 8018
rect 1152 7944 58848 7966
rect 12115 7898 12173 7904
rect 12115 7864 12127 7898
rect 12161 7895 12173 7898
rect 12400 7895 12406 7907
rect 12161 7867 12406 7895
rect 12161 7864 12173 7867
rect 12115 7858 12173 7864
rect 12400 7855 12406 7867
rect 12458 7855 12464 7907
rect 12784 7895 12790 7907
rect 12745 7867 12790 7895
rect 12784 7855 12790 7867
rect 12842 7855 12848 7907
rect 13552 7895 13558 7907
rect 13513 7867 13558 7895
rect 13552 7855 13558 7867
rect 13610 7855 13616 7907
rect 14992 7855 14998 7907
rect 15050 7895 15056 7907
rect 15091 7898 15149 7904
rect 15091 7895 15103 7898
rect 15050 7867 15103 7895
rect 15050 7855 15056 7867
rect 15091 7864 15103 7867
rect 15137 7864 15149 7898
rect 15091 7858 15149 7864
rect 17683 7898 17741 7904
rect 17683 7864 17695 7898
rect 17729 7895 17741 7898
rect 17968 7895 17974 7907
rect 17729 7867 17974 7895
rect 17729 7864 17741 7867
rect 17683 7858 17741 7864
rect 17968 7855 17974 7867
rect 18026 7855 18032 7907
rect 27952 7895 27958 7907
rect 27913 7867 27958 7895
rect 27952 7855 27958 7867
rect 28010 7895 28016 7907
rect 30832 7895 30838 7907
rect 28010 7867 28382 7895
rect 30793 7867 30838 7895
rect 28010 7855 28016 7867
rect 4531 7824 4589 7830
rect 4531 7790 4543 7824
rect 4577 7821 4589 7824
rect 23056 7821 23062 7833
rect 4577 7793 23062 7821
rect 4577 7790 4589 7793
rect 4531 7784 4589 7790
rect 3280 7707 3286 7759
rect 3338 7747 3344 7759
rect 3955 7750 4013 7756
rect 3955 7747 3967 7750
rect 3338 7719 3967 7747
rect 3338 7707 3344 7719
rect 3955 7716 3967 7719
rect 4001 7716 4013 7750
rect 3955 7710 4013 7716
rect 4048 7707 4054 7759
rect 4106 7747 4112 7759
rect 4834 7756 4862 7793
rect 23056 7781 23062 7793
rect 23114 7781 23120 7833
rect 4723 7750 4781 7756
rect 4723 7747 4735 7750
rect 4106 7719 4735 7747
rect 4106 7707 4112 7719
rect 4723 7716 4735 7719
rect 4769 7716 4781 7750
rect 4723 7710 4781 7716
rect 4819 7750 4877 7756
rect 4819 7716 4831 7750
rect 4865 7716 4877 7750
rect 4819 7710 4877 7716
rect 10099 7750 10157 7756
rect 10099 7716 10111 7750
rect 10145 7747 10157 7750
rect 10192 7747 10198 7759
rect 10145 7719 10198 7747
rect 10145 7716 10157 7719
rect 10099 7710 10157 7716
rect 10192 7707 10198 7719
rect 10250 7707 10256 7759
rect 10579 7750 10637 7756
rect 10579 7716 10591 7750
rect 10625 7747 10637 7750
rect 10864 7747 10870 7759
rect 10625 7719 10870 7747
rect 10625 7716 10637 7719
rect 10579 7710 10637 7716
rect 10864 7707 10870 7719
rect 10922 7707 10928 7759
rect 11344 7707 11350 7759
rect 11402 7747 11408 7759
rect 12307 7750 12365 7756
rect 12307 7747 12319 7750
rect 11402 7719 12319 7747
rect 11402 7707 11408 7719
rect 12307 7716 12319 7719
rect 12353 7716 12365 7750
rect 12307 7710 12365 7716
rect 12400 7707 12406 7759
rect 12458 7747 12464 7759
rect 12458 7719 12503 7747
rect 12458 7707 12464 7719
rect 12784 7707 12790 7759
rect 12842 7747 12848 7759
rect 13363 7750 13421 7756
rect 13363 7747 13375 7750
rect 12842 7719 13375 7747
rect 12842 7707 12848 7719
rect 13363 7716 13375 7719
rect 13409 7716 13421 7750
rect 13363 7710 13421 7716
rect 13552 7707 13558 7759
rect 13610 7747 13616 7759
rect 13939 7750 13997 7756
rect 13939 7747 13951 7750
rect 13610 7719 13951 7747
rect 13610 7707 13616 7719
rect 13939 7716 13951 7719
rect 13985 7716 13997 7750
rect 13939 7710 13997 7716
rect 14992 7707 14998 7759
rect 15050 7747 15056 7759
rect 15379 7750 15437 7756
rect 15379 7747 15391 7750
rect 15050 7719 15391 7747
rect 15050 7707 15056 7719
rect 15379 7716 15391 7719
rect 15425 7716 15437 7750
rect 15379 7710 15437 7716
rect 15955 7750 16013 7756
rect 15955 7716 15967 7750
rect 16001 7747 16013 7750
rect 16240 7747 16246 7759
rect 16001 7719 16246 7747
rect 16001 7716 16013 7719
rect 15955 7710 16013 7716
rect 16240 7707 16246 7719
rect 16298 7707 16304 7759
rect 20659 7750 20717 7756
rect 20659 7716 20671 7750
rect 20705 7747 20717 7750
rect 20947 7750 21005 7756
rect 20947 7747 20959 7750
rect 20705 7719 20959 7747
rect 20705 7716 20717 7719
rect 20659 7710 20717 7716
rect 20947 7716 20959 7719
rect 20993 7747 21005 7750
rect 21040 7747 21046 7759
rect 20993 7719 21046 7747
rect 20993 7716 21005 7719
rect 20947 7710 21005 7716
rect 21040 7707 21046 7719
rect 21098 7707 21104 7759
rect 23920 7747 23926 7759
rect 23881 7719 23926 7747
rect 23920 7707 23926 7719
rect 23978 7707 23984 7759
rect 24403 7750 24461 7756
rect 24403 7716 24415 7750
rect 24449 7747 24461 7750
rect 24688 7747 24694 7759
rect 24449 7719 24694 7747
rect 24449 7716 24461 7719
rect 24403 7710 24461 7716
rect 24688 7707 24694 7719
rect 24746 7707 24752 7759
rect 25459 7750 25517 7756
rect 25459 7716 25471 7750
rect 25505 7747 25517 7750
rect 25936 7747 25942 7759
rect 25505 7719 25942 7747
rect 25505 7716 25517 7719
rect 25459 7710 25517 7716
rect 25936 7707 25942 7719
rect 25994 7707 26000 7759
rect 26224 7747 26230 7759
rect 26185 7719 26230 7747
rect 26224 7707 26230 7719
rect 26282 7707 26288 7759
rect 26992 7747 26998 7759
rect 26953 7719 26998 7747
rect 26992 7707 26998 7719
rect 27050 7707 27056 7759
rect 28354 7756 28382 7867
rect 30832 7855 30838 7867
rect 30890 7855 30896 7907
rect 32368 7895 32374 7907
rect 32329 7867 32374 7895
rect 32368 7855 32374 7867
rect 32426 7855 32432 7907
rect 35827 7898 35885 7904
rect 35827 7864 35839 7898
rect 35873 7895 35885 7898
rect 35920 7895 35926 7907
rect 35873 7867 35926 7895
rect 35873 7864 35885 7867
rect 35827 7858 35885 7864
rect 35920 7855 35926 7867
rect 35978 7895 35984 7907
rect 39952 7895 39958 7907
rect 35978 7867 36062 7895
rect 39913 7867 39958 7895
rect 35978 7855 35984 7867
rect 28339 7750 28397 7756
rect 28339 7716 28351 7750
rect 28385 7716 28397 7750
rect 28339 7710 28397 7716
rect 29107 7750 29165 7756
rect 29107 7716 29119 7750
rect 29153 7747 29165 7750
rect 29392 7747 29398 7759
rect 29153 7719 29398 7747
rect 29153 7716 29165 7719
rect 29107 7710 29165 7716
rect 29392 7707 29398 7719
rect 29450 7707 29456 7759
rect 29875 7750 29933 7756
rect 29875 7716 29887 7750
rect 29921 7747 29933 7750
rect 30160 7747 30166 7759
rect 29921 7719 30166 7747
rect 29921 7716 29933 7719
rect 29875 7710 29933 7716
rect 30160 7707 30166 7719
rect 30218 7707 30224 7759
rect 30850 7747 30878 7855
rect 31123 7750 31181 7756
rect 31123 7747 31135 7750
rect 30850 7719 31135 7747
rect 31123 7716 31135 7719
rect 31169 7716 31181 7750
rect 31123 7710 31181 7716
rect 34291 7750 34349 7756
rect 34291 7716 34303 7750
rect 34337 7747 34349 7750
rect 34576 7747 34582 7759
rect 34337 7719 34582 7747
rect 34337 7716 34349 7719
rect 34291 7710 34349 7716
rect 34576 7707 34582 7719
rect 34634 7707 34640 7759
rect 35344 7747 35350 7759
rect 35305 7719 35350 7747
rect 35344 7707 35350 7719
rect 35402 7707 35408 7759
rect 36034 7756 36062 7867
rect 39952 7855 39958 7867
rect 40010 7895 40016 7907
rect 43696 7895 43702 7907
rect 40010 7867 40286 7895
rect 43657 7867 43702 7895
rect 40010 7855 40016 7867
rect 36019 7750 36077 7756
rect 36019 7716 36031 7750
rect 36065 7716 36077 7750
rect 36019 7710 36077 7716
rect 36595 7750 36653 7756
rect 36595 7716 36607 7750
rect 36641 7747 36653 7750
rect 36784 7747 36790 7759
rect 36641 7719 36790 7747
rect 36641 7716 36653 7719
rect 36595 7710 36653 7716
rect 36784 7707 36790 7719
rect 36842 7707 36848 7759
rect 38800 7747 38806 7759
rect 38761 7719 38806 7747
rect 38800 7707 38806 7719
rect 38858 7707 38864 7759
rect 39283 7750 39341 7756
rect 39283 7716 39295 7750
rect 39329 7747 39341 7750
rect 39472 7747 39478 7759
rect 39329 7719 39478 7747
rect 39329 7716 39341 7719
rect 39283 7710 39341 7716
rect 39472 7707 39478 7719
rect 39530 7707 39536 7759
rect 40258 7756 40286 7867
rect 43696 7855 43702 7867
rect 43754 7895 43760 7907
rect 44464 7895 44470 7907
rect 43754 7867 44126 7895
rect 44425 7867 44470 7895
rect 43754 7855 43760 7867
rect 40243 7750 40301 7756
rect 40243 7716 40255 7750
rect 40289 7716 40301 7750
rect 41104 7747 41110 7759
rect 41065 7719 41110 7747
rect 40243 7710 40301 7716
rect 41104 7707 41110 7719
rect 41162 7707 41168 7759
rect 41872 7747 41878 7759
rect 41833 7719 41878 7747
rect 41872 7707 41878 7719
rect 41930 7707 41936 7759
rect 42355 7750 42413 7756
rect 42355 7716 42367 7750
rect 42401 7747 42413 7750
rect 42640 7747 42646 7759
rect 42401 7719 42646 7747
rect 42401 7716 42413 7719
rect 42355 7710 42413 7716
rect 42640 7707 42646 7719
rect 42698 7707 42704 7759
rect 44098 7756 44126 7867
rect 44464 7855 44470 7867
rect 44522 7895 44528 7907
rect 45232 7895 45238 7907
rect 44522 7867 44798 7895
rect 45193 7867 45238 7895
rect 44522 7855 44528 7867
rect 44770 7756 44798 7867
rect 45232 7855 45238 7867
rect 45290 7895 45296 7907
rect 46864 7895 46870 7907
rect 45290 7867 45566 7895
rect 46825 7867 46870 7895
rect 45290 7855 45296 7867
rect 45538 7756 45566 7867
rect 46864 7855 46870 7867
rect 46922 7895 46928 7907
rect 48976 7895 48982 7907
rect 46922 7867 47102 7895
rect 48937 7867 48982 7895
rect 46922 7855 46928 7867
rect 44083 7750 44141 7756
rect 44083 7716 44095 7750
rect 44129 7716 44141 7750
rect 44083 7710 44141 7716
rect 44755 7750 44813 7756
rect 44755 7716 44767 7750
rect 44801 7716 44813 7750
rect 44755 7710 44813 7716
rect 45523 7750 45581 7756
rect 45523 7716 45535 7750
rect 45569 7716 45581 7750
rect 46384 7747 46390 7759
rect 46345 7719 46390 7747
rect 45523 7710 45581 7716
rect 46384 7707 46390 7719
rect 46442 7707 46448 7759
rect 47074 7756 47102 7867
rect 48976 7855 48982 7867
rect 49034 7855 49040 7907
rect 49744 7895 49750 7907
rect 49705 7867 49750 7895
rect 49744 7855 49750 7867
rect 49802 7855 49808 7907
rect 47059 7750 47117 7756
rect 47059 7716 47071 7750
rect 47105 7716 47117 7750
rect 47059 7710 47117 7716
rect 47824 7707 47830 7759
rect 47882 7747 47888 7759
rect 47923 7750 47981 7756
rect 47923 7747 47935 7750
rect 47882 7719 47935 7747
rect 47882 7707 47888 7719
rect 47923 7716 47935 7719
rect 47969 7716 47981 7750
rect 48994 7747 49022 7855
rect 49267 7750 49325 7756
rect 49267 7747 49279 7750
rect 48994 7719 49279 7747
rect 47923 7710 47981 7716
rect 49267 7716 49279 7719
rect 49313 7716 49325 7750
rect 49762 7747 49790 7855
rect 50035 7750 50093 7756
rect 50035 7747 50047 7750
rect 49762 7719 50047 7747
rect 49267 7710 49325 7716
rect 50035 7716 50047 7719
rect 50081 7716 50093 7750
rect 51088 7747 51094 7759
rect 51049 7719 51094 7747
rect 50035 7710 50093 7716
rect 51088 7707 51094 7719
rect 51146 7707 51152 7759
rect 52624 7747 52630 7759
rect 52585 7719 52630 7747
rect 52624 7707 52630 7719
rect 52682 7707 52688 7759
rect 52720 7707 52726 7759
rect 52778 7747 52784 7759
rect 53395 7750 53453 7756
rect 53395 7747 53407 7750
rect 52778 7719 53407 7747
rect 52778 7707 52784 7719
rect 53395 7716 53407 7719
rect 53441 7716 53453 7750
rect 53395 7710 53453 7716
rect 1456 7633 1462 7685
rect 1514 7673 1520 7685
rect 1555 7676 1613 7682
rect 1555 7673 1567 7676
rect 1514 7645 1567 7673
rect 1514 7633 1520 7645
rect 1555 7642 1567 7645
rect 1601 7642 1613 7676
rect 1555 7636 1613 7642
rect 2227 7676 2285 7682
rect 2227 7642 2239 7676
rect 2273 7673 2285 7676
rect 2515 7676 2573 7682
rect 2515 7673 2527 7676
rect 2273 7645 2527 7673
rect 2273 7642 2285 7645
rect 2227 7636 2285 7642
rect 2515 7642 2527 7645
rect 2561 7673 2573 7676
rect 3568 7673 3574 7685
rect 2561 7645 3574 7673
rect 2561 7642 2573 7645
rect 2515 7636 2573 7642
rect 3568 7633 3574 7645
rect 3626 7633 3632 7685
rect 5587 7676 5645 7682
rect 5587 7642 5599 7676
rect 5633 7673 5645 7676
rect 23152 7673 23158 7685
rect 5633 7645 23158 7673
rect 5633 7642 5645 7645
rect 5587 7636 5645 7642
rect 23152 7633 23158 7645
rect 23210 7633 23216 7685
rect 53107 7676 53165 7682
rect 53107 7642 53119 7676
rect 53153 7673 53165 7676
rect 53200 7673 53206 7685
rect 53153 7645 53206 7673
rect 53153 7642 53165 7645
rect 53107 7636 53165 7642
rect 53200 7633 53206 7645
rect 53258 7673 53264 7685
rect 53299 7676 53357 7682
rect 53299 7673 53311 7676
rect 53258 7645 53311 7673
rect 53258 7633 53264 7645
rect 53299 7642 53311 7645
rect 53345 7642 53357 7676
rect 53299 7636 53357 7642
rect 55123 7676 55181 7682
rect 55123 7642 55135 7676
rect 55169 7642 55181 7676
rect 55792 7673 55798 7685
rect 55753 7645 55798 7673
rect 55123 7636 55181 7642
rect 2995 7602 3053 7608
rect 2995 7568 3007 7602
rect 3041 7599 3053 7602
rect 3283 7602 3341 7608
rect 3283 7599 3295 7602
rect 3041 7571 3295 7599
rect 3041 7568 3053 7571
rect 2995 7562 3053 7568
rect 3283 7568 3295 7571
rect 3329 7568 3341 7602
rect 3283 7562 3341 7568
rect 4051 7602 4109 7608
rect 4051 7568 4063 7602
rect 4097 7599 4109 7602
rect 4144 7599 4150 7611
rect 4097 7571 4150 7599
rect 4097 7568 4109 7571
rect 4051 7562 4109 7568
rect 3298 7525 3326 7562
rect 4144 7559 4150 7571
rect 4202 7559 4208 7611
rect 9331 7602 9389 7608
rect 9331 7568 9343 7602
rect 9377 7568 9389 7602
rect 9331 7562 9389 7568
rect 6832 7525 6838 7537
rect 3298 7497 6838 7525
rect 6832 7485 6838 7497
rect 6890 7485 6896 7537
rect 9346 7525 9374 7562
rect 12880 7559 12886 7611
rect 12938 7599 12944 7611
rect 13075 7602 13133 7608
rect 13075 7599 13087 7602
rect 12938 7571 13087 7599
rect 12938 7559 12944 7571
rect 13075 7568 13087 7571
rect 13121 7568 13133 7602
rect 13075 7562 13133 7568
rect 13282 7571 15518 7599
rect 13282 7525 13310 7571
rect 9346 7497 13310 7525
rect 13363 7528 13421 7534
rect 13363 7494 13375 7528
rect 13409 7525 13421 7528
rect 15490 7525 15518 7571
rect 18352 7559 18358 7611
rect 18410 7599 18416 7611
rect 18643 7602 18701 7608
rect 18643 7599 18655 7602
rect 18410 7571 18655 7599
rect 18410 7559 18416 7571
rect 18643 7568 18655 7571
rect 18689 7568 18701 7602
rect 18643 7562 18701 7568
rect 21715 7602 21773 7608
rect 21715 7568 21727 7602
rect 21761 7568 21773 7602
rect 21715 7562 21773 7568
rect 33811 7602 33869 7608
rect 33811 7568 33823 7602
rect 33857 7599 33869 7602
rect 34096 7599 34102 7611
rect 33857 7571 34102 7599
rect 33857 7568 33869 7571
rect 33811 7562 33869 7568
rect 21730 7525 21758 7562
rect 34096 7559 34102 7571
rect 34154 7559 34160 7611
rect 51859 7602 51917 7608
rect 51859 7568 51871 7602
rect 51905 7599 51917 7602
rect 52912 7599 52918 7611
rect 51905 7571 52918 7599
rect 51905 7568 51917 7571
rect 51859 7562 51917 7568
rect 52912 7559 52918 7571
rect 52970 7559 52976 7611
rect 55138 7599 55166 7636
rect 55792 7633 55798 7645
rect 55850 7633 55856 7685
rect 56176 7633 56182 7685
rect 56234 7673 56240 7685
rect 56563 7676 56621 7682
rect 56563 7673 56575 7676
rect 56234 7645 56575 7673
rect 56234 7633 56240 7645
rect 56563 7642 56575 7645
rect 56609 7642 56621 7676
rect 57328 7673 57334 7685
rect 57289 7645 57334 7673
rect 56563 7636 56621 7642
rect 57328 7633 57334 7645
rect 57386 7633 57392 7685
rect 58768 7599 58774 7611
rect 55138 7571 58774 7599
rect 58768 7559 58774 7571
rect 58826 7559 58832 7611
rect 13409 7497 13886 7525
rect 15490 7497 21758 7525
rect 13409 7494 13421 7497
rect 13363 7488 13421 7494
rect 2416 7451 2422 7463
rect 2377 7423 2422 7451
rect 2416 7411 2422 7423
rect 2474 7411 2480 7463
rect 3187 7454 3245 7460
rect 3187 7420 3199 7454
rect 3233 7451 3245 7454
rect 3376 7451 3382 7463
rect 3233 7423 3382 7451
rect 3233 7420 3245 7423
rect 3187 7414 3245 7420
rect 3376 7411 3382 7423
rect 3434 7411 3440 7463
rect 5296 7411 5302 7463
rect 5354 7451 5360 7463
rect 5491 7454 5549 7460
rect 5491 7451 5503 7454
rect 5354 7423 5503 7451
rect 5354 7411 5360 7423
rect 5491 7420 5503 7423
rect 5537 7420 5549 7454
rect 5491 7414 5549 7420
rect 9136 7411 9142 7463
rect 9194 7451 9200 7463
rect 9235 7454 9293 7460
rect 9235 7451 9247 7454
rect 9194 7423 9247 7451
rect 9194 7411 9200 7423
rect 9235 7420 9247 7423
rect 9281 7420 9293 7454
rect 9235 7414 9293 7420
rect 9904 7411 9910 7463
rect 9962 7451 9968 7463
rect 10003 7454 10061 7460
rect 10003 7451 10015 7454
rect 9962 7423 10015 7451
rect 9962 7411 9968 7423
rect 10003 7420 10015 7423
rect 10049 7420 10061 7454
rect 10003 7414 10061 7420
rect 10771 7454 10829 7460
rect 10771 7420 10783 7454
rect 10817 7451 10829 7454
rect 11056 7451 11062 7463
rect 10817 7423 11062 7451
rect 10817 7420 10829 7423
rect 10771 7414 10829 7420
rect 11056 7411 11062 7423
rect 11114 7411 11120 7463
rect 12208 7411 12214 7463
rect 12266 7451 12272 7463
rect 13858 7460 13886 7497
rect 39952 7485 39958 7537
rect 40010 7525 40016 7537
rect 40010 7497 41054 7525
rect 40010 7485 40016 7497
rect 13171 7454 13229 7460
rect 13171 7451 13183 7454
rect 12266 7423 13183 7451
rect 12266 7411 12272 7423
rect 13171 7420 13183 7423
rect 13217 7420 13229 7454
rect 13171 7414 13229 7420
rect 13843 7454 13901 7460
rect 13843 7420 13855 7454
rect 13889 7420 13901 7454
rect 13843 7414 13901 7420
rect 15280 7411 15286 7463
rect 15338 7451 15344 7463
rect 15475 7454 15533 7460
rect 15475 7451 15487 7454
rect 15338 7423 15487 7451
rect 15338 7411 15344 7423
rect 15475 7420 15487 7423
rect 15521 7420 15533 7454
rect 15475 7414 15533 7420
rect 15664 7411 15670 7463
rect 15722 7451 15728 7463
rect 16147 7454 16205 7460
rect 16147 7451 16159 7454
rect 15722 7423 16159 7451
rect 15722 7411 15728 7423
rect 16147 7420 16159 7423
rect 16193 7420 16205 7454
rect 16147 7414 16205 7420
rect 20752 7411 20758 7463
rect 20810 7451 20816 7463
rect 20851 7454 20909 7460
rect 20851 7451 20863 7454
rect 20810 7423 20863 7451
rect 20810 7411 20816 7423
rect 20851 7420 20863 7423
rect 20897 7420 20909 7454
rect 20851 7414 20909 7420
rect 23728 7411 23734 7463
rect 23786 7451 23792 7463
rect 23827 7454 23885 7460
rect 23827 7451 23839 7454
rect 23786 7423 23839 7451
rect 23786 7411 23792 7423
rect 23827 7420 23839 7423
rect 23873 7420 23885 7454
rect 24592 7451 24598 7463
rect 24553 7423 24598 7451
rect 23827 7414 23885 7420
rect 24592 7411 24598 7423
rect 24650 7411 24656 7463
rect 24784 7411 24790 7463
rect 24842 7451 24848 7463
rect 25363 7454 25421 7460
rect 25363 7451 25375 7454
rect 24842 7423 25375 7451
rect 24842 7411 24848 7423
rect 25363 7420 25375 7423
rect 25409 7420 25421 7454
rect 25363 7414 25421 7420
rect 25936 7411 25942 7463
rect 25994 7451 26000 7463
rect 26131 7454 26189 7460
rect 26131 7451 26143 7454
rect 25994 7423 26143 7451
rect 25994 7411 26000 7423
rect 26131 7420 26143 7423
rect 26177 7420 26189 7454
rect 26131 7414 26189 7420
rect 26704 7411 26710 7463
rect 26762 7451 26768 7463
rect 26899 7454 26957 7460
rect 26899 7451 26911 7454
rect 26762 7423 26911 7451
rect 26762 7411 26768 7423
rect 26899 7420 26911 7423
rect 26945 7420 26957 7454
rect 26899 7414 26957 7420
rect 28144 7411 28150 7463
rect 28202 7451 28208 7463
rect 28243 7454 28301 7460
rect 28243 7451 28255 7454
rect 28202 7423 28255 7451
rect 28202 7411 28208 7423
rect 28243 7420 28255 7423
rect 28289 7420 28301 7454
rect 28243 7414 28301 7420
rect 29200 7411 29206 7463
rect 29258 7451 29264 7463
rect 29299 7454 29357 7460
rect 29299 7451 29311 7454
rect 29258 7423 29311 7451
rect 29258 7411 29264 7423
rect 29299 7420 29311 7423
rect 29345 7420 29357 7454
rect 29299 7414 29357 7420
rect 29584 7411 29590 7463
rect 29642 7451 29648 7463
rect 30067 7454 30125 7460
rect 30067 7451 30079 7454
rect 29642 7423 30079 7451
rect 29642 7411 29648 7423
rect 30067 7420 30079 7423
rect 30113 7420 30125 7454
rect 30067 7414 30125 7420
rect 31024 7411 31030 7463
rect 31082 7451 31088 7463
rect 31219 7454 31277 7460
rect 31219 7451 31231 7454
rect 31082 7423 31231 7451
rect 31082 7411 31088 7423
rect 31219 7420 31231 7423
rect 31265 7420 31277 7454
rect 31219 7414 31277 7420
rect 33616 7411 33622 7463
rect 33674 7451 33680 7463
rect 33715 7454 33773 7460
rect 33715 7451 33727 7454
rect 33674 7423 33727 7451
rect 33674 7411 33680 7423
rect 33715 7420 33727 7423
rect 33761 7420 33773 7454
rect 33715 7414 33773 7420
rect 34384 7411 34390 7463
rect 34442 7451 34448 7463
rect 34483 7454 34541 7460
rect 34483 7451 34495 7454
rect 34442 7423 34495 7451
rect 34442 7411 34448 7423
rect 34483 7420 34495 7423
rect 34529 7420 34541 7454
rect 34483 7414 34541 7420
rect 34768 7411 34774 7463
rect 34826 7451 34832 7463
rect 35251 7454 35309 7460
rect 35251 7451 35263 7454
rect 34826 7423 35263 7451
rect 34826 7411 34832 7423
rect 35251 7420 35263 7423
rect 35297 7420 35309 7454
rect 35251 7414 35309 7420
rect 36016 7411 36022 7463
rect 36074 7451 36080 7463
rect 36115 7454 36173 7460
rect 36115 7451 36127 7454
rect 36074 7423 36127 7451
rect 36074 7411 36080 7423
rect 36115 7420 36127 7423
rect 36161 7420 36173 7454
rect 36115 7414 36173 7420
rect 36592 7411 36598 7463
rect 36650 7451 36656 7463
rect 36883 7454 36941 7460
rect 36883 7451 36895 7454
rect 36650 7423 36895 7451
rect 36650 7411 36656 7423
rect 36883 7420 36895 7423
rect 36929 7420 36941 7454
rect 36883 7414 36941 7420
rect 38032 7411 38038 7463
rect 38090 7451 38096 7463
rect 38707 7454 38765 7460
rect 38707 7451 38719 7454
rect 38090 7423 38719 7451
rect 38090 7411 38096 7423
rect 38707 7420 38719 7423
rect 38753 7420 38765 7454
rect 38707 7414 38765 7420
rect 38800 7411 38806 7463
rect 38858 7451 38864 7463
rect 39571 7454 39629 7460
rect 39571 7451 39583 7454
rect 38858 7423 39583 7451
rect 38858 7411 38864 7423
rect 39571 7420 39583 7423
rect 39617 7420 39629 7454
rect 39571 7414 39629 7420
rect 39664 7411 39670 7463
rect 39722 7451 39728 7463
rect 41026 7460 41054 7497
rect 41680 7485 41686 7537
rect 41738 7525 41744 7537
rect 41738 7497 42590 7525
rect 41738 7485 41744 7497
rect 40339 7454 40397 7460
rect 40339 7451 40351 7454
rect 39722 7423 40351 7451
rect 39722 7411 39728 7423
rect 40339 7420 40351 7423
rect 40385 7420 40397 7454
rect 40339 7414 40397 7420
rect 41011 7454 41069 7460
rect 41011 7420 41023 7454
rect 41057 7420 41069 7454
rect 41011 7414 41069 7420
rect 41104 7411 41110 7463
rect 41162 7451 41168 7463
rect 42562 7460 42590 7497
rect 45424 7485 45430 7537
rect 45482 7525 45488 7537
rect 45482 7497 46334 7525
rect 45482 7485 45488 7497
rect 41779 7454 41837 7460
rect 41779 7451 41791 7454
rect 41162 7423 41791 7451
rect 41162 7411 41168 7423
rect 41779 7420 41791 7423
rect 41825 7420 41837 7454
rect 41779 7414 41837 7420
rect 42547 7454 42605 7460
rect 42547 7420 42559 7454
rect 42593 7420 42605 7454
rect 42547 7414 42605 7420
rect 43216 7411 43222 7463
rect 43274 7451 43280 7463
rect 43987 7454 44045 7460
rect 43987 7451 43999 7454
rect 43274 7423 43999 7451
rect 43274 7411 43280 7423
rect 43987 7420 43999 7423
rect 44033 7420 44045 7454
rect 43987 7414 44045 7420
rect 44368 7411 44374 7463
rect 44426 7451 44432 7463
rect 44851 7454 44909 7460
rect 44851 7451 44863 7454
rect 44426 7423 44863 7451
rect 44426 7411 44432 7423
rect 44851 7420 44863 7423
rect 44897 7420 44909 7454
rect 44851 7414 44909 7420
rect 45040 7411 45046 7463
rect 45098 7451 45104 7463
rect 46306 7460 46334 7497
rect 46864 7485 46870 7537
rect 46922 7525 46928 7537
rect 59344 7525 59350 7537
rect 46922 7497 47870 7525
rect 46922 7485 46928 7497
rect 45619 7454 45677 7460
rect 45619 7451 45631 7454
rect 45098 7423 45631 7451
rect 45098 7411 45104 7423
rect 45619 7420 45631 7423
rect 45665 7420 45677 7454
rect 45619 7414 45677 7420
rect 46291 7454 46349 7460
rect 46291 7420 46303 7454
rect 46337 7420 46349 7454
rect 46291 7414 46349 7420
rect 46384 7411 46390 7463
rect 46442 7451 46448 7463
rect 47842 7460 47870 7497
rect 51010 7497 59350 7525
rect 47155 7454 47213 7460
rect 47155 7451 47167 7454
rect 46442 7423 47167 7451
rect 46442 7411 46448 7423
rect 47155 7420 47167 7423
rect 47201 7420 47213 7454
rect 47155 7414 47213 7420
rect 47827 7454 47885 7460
rect 47827 7420 47839 7454
rect 47873 7420 47885 7454
rect 47827 7414 47885 7420
rect 48304 7411 48310 7463
rect 48362 7451 48368 7463
rect 49363 7454 49421 7460
rect 49363 7451 49375 7454
rect 48362 7423 49375 7451
rect 48362 7411 48368 7423
rect 49363 7420 49375 7423
rect 49409 7420 49421 7454
rect 49363 7414 49421 7420
rect 50032 7411 50038 7463
rect 50090 7451 50096 7463
rect 51010 7460 51038 7497
rect 59344 7485 59350 7497
rect 59402 7485 59408 7537
rect 50131 7454 50189 7460
rect 50131 7451 50143 7454
rect 50090 7423 50143 7451
rect 50090 7411 50096 7423
rect 50131 7420 50143 7423
rect 50177 7420 50189 7454
rect 50131 7414 50189 7420
rect 50995 7454 51053 7460
rect 50995 7420 51007 7454
rect 51041 7420 51053 7454
rect 50995 7414 51053 7420
rect 51664 7411 51670 7463
rect 51722 7451 51728 7463
rect 51763 7454 51821 7460
rect 51763 7451 51775 7454
rect 51722 7423 51775 7451
rect 51722 7411 51728 7423
rect 51763 7420 51775 7423
rect 51809 7420 51821 7454
rect 51763 7414 51821 7420
rect 52336 7411 52342 7463
rect 52394 7451 52400 7463
rect 52531 7454 52589 7460
rect 52531 7451 52543 7454
rect 52394 7423 52543 7451
rect 52394 7411 52400 7423
rect 52531 7420 52543 7423
rect 52577 7420 52589 7454
rect 52531 7414 52589 7420
rect 1152 7352 58848 7374
rect 1152 7300 19654 7352
rect 19706 7300 19718 7352
rect 19770 7300 19782 7352
rect 19834 7300 19846 7352
rect 19898 7300 50374 7352
rect 50426 7300 50438 7352
rect 50490 7300 50502 7352
rect 50554 7300 50566 7352
rect 50618 7300 58848 7352
rect 1152 7278 58848 7300
rect 17203 7232 17261 7238
rect 17203 7198 17215 7232
rect 17249 7198 17261 7232
rect 17203 7192 17261 7198
rect 31603 7232 31661 7238
rect 31603 7198 31615 7232
rect 31649 7198 31661 7232
rect 31603 7192 31661 7198
rect 6448 7155 6454 7167
rect 6409 7127 6454 7155
rect 6448 7115 6454 7127
rect 6506 7155 6512 7167
rect 7984 7155 7990 7167
rect 6506 7127 6878 7155
rect 7945 7127 7990 7155
rect 6506 7115 6512 7127
rect 6850 7090 6878 7127
rect 7984 7115 7990 7127
rect 8042 7155 8048 7167
rect 17011 7158 17069 7164
rect 17011 7155 17023 7158
rect 8042 7127 8414 7155
rect 8042 7115 8048 7127
rect 6835 7084 6893 7090
rect 6835 7050 6847 7084
rect 6881 7050 6893 7084
rect 6835 7044 6893 7050
rect 7315 7084 7373 7090
rect 7315 7050 7327 7084
rect 7361 7081 7373 7084
rect 7600 7081 7606 7093
rect 7361 7053 7606 7081
rect 7361 7050 7373 7053
rect 7315 7044 7373 7050
rect 7600 7041 7606 7053
rect 7658 7041 7664 7093
rect 8386 7090 8414 7127
rect 9826 7127 17023 7155
rect 9826 7090 9854 7127
rect 17011 7124 17023 7127
rect 17057 7124 17069 7158
rect 17011 7118 17069 7124
rect 17104 7115 17110 7167
rect 17162 7155 17168 7167
rect 17218 7155 17246 7192
rect 22288 7155 22294 7167
rect 17162 7127 17246 7155
rect 17698 7127 21182 7155
rect 22249 7127 22294 7155
rect 17162 7115 17168 7127
rect 8371 7084 8429 7090
rect 8371 7050 8383 7084
rect 8417 7050 8429 7084
rect 8371 7044 8429 7050
rect 9811 7084 9869 7090
rect 9811 7050 9823 7084
rect 9857 7050 9869 7084
rect 9811 7044 9869 7050
rect 15091 7084 15149 7090
rect 15091 7050 15103 7084
rect 15137 7081 15149 7084
rect 15184 7081 15190 7093
rect 15137 7053 15190 7081
rect 15137 7050 15149 7053
rect 15091 7044 15149 7050
rect 15184 7041 15190 7053
rect 15242 7041 15248 7093
rect 15760 7041 15766 7093
rect 15818 7081 15824 7093
rect 15859 7084 15917 7090
rect 15859 7081 15871 7084
rect 15818 7053 15871 7081
rect 15818 7041 15824 7053
rect 15859 7050 15871 7053
rect 15905 7050 15917 7084
rect 15859 7044 15917 7050
rect 16528 7041 16534 7093
rect 16586 7081 16592 7093
rect 17698 7081 17726 7127
rect 16586 7053 17726 7081
rect 17779 7084 17837 7090
rect 16586 7041 16592 7053
rect 17779 7050 17791 7084
rect 17825 7081 17837 7084
rect 18064 7081 18070 7093
rect 17825 7053 18070 7081
rect 17825 7050 17837 7053
rect 17779 7044 17837 7050
rect 18064 7041 18070 7053
rect 18122 7041 18128 7093
rect 18832 7081 18838 7093
rect 18793 7053 18838 7081
rect 18832 7041 18838 7053
rect 18890 7041 18896 7093
rect 20083 7084 20141 7090
rect 20083 7050 20095 7084
rect 20129 7081 20141 7084
rect 20368 7081 20374 7093
rect 20129 7053 20374 7081
rect 20129 7050 20141 7053
rect 20083 7044 20141 7050
rect 20368 7041 20374 7053
rect 20426 7041 20432 7093
rect 21154 7090 21182 7127
rect 22288 7115 22294 7127
rect 22346 7155 22352 7167
rect 22346 7127 22622 7155
rect 22346 7115 22352 7127
rect 21139 7084 21197 7090
rect 21139 7050 21151 7084
rect 21185 7050 21197 7084
rect 21904 7081 21910 7093
rect 21865 7053 21910 7081
rect 21139 7044 21197 7050
rect 21904 7041 21910 7053
rect 21962 7041 21968 7093
rect 22594 7090 22622 7127
rect 23056 7115 23062 7167
rect 23114 7155 23120 7167
rect 28048 7155 28054 7167
rect 23114 7127 28054 7155
rect 23114 7115 23120 7127
rect 28048 7115 28054 7127
rect 28106 7115 28112 7167
rect 28336 7155 28342 7167
rect 28297 7127 28342 7155
rect 28336 7115 28342 7127
rect 28394 7155 28400 7167
rect 28394 7127 28670 7155
rect 28394 7115 28400 7127
rect 22579 7084 22637 7090
rect 22579 7050 22591 7084
rect 22625 7050 22637 7084
rect 23440 7081 23446 7093
rect 23401 7053 23446 7081
rect 22579 7044 22637 7050
rect 23440 7041 23446 7053
rect 23498 7041 23504 7093
rect 24208 7081 24214 7093
rect 24169 7053 24214 7081
rect 24208 7041 24214 7053
rect 24266 7041 24272 7093
rect 25648 7081 25654 7093
rect 25609 7053 25654 7081
rect 25648 7041 25654 7053
rect 25706 7041 25712 7093
rect 26416 7081 26422 7093
rect 26377 7053 26422 7081
rect 26416 7041 26422 7053
rect 26474 7041 26480 7093
rect 27184 7081 27190 7093
rect 27145 7053 27190 7081
rect 27184 7041 27190 7053
rect 27242 7041 27248 7093
rect 27955 7084 28013 7090
rect 27955 7050 27967 7084
rect 28001 7081 28013 7084
rect 28240 7081 28246 7093
rect 28001 7053 28246 7081
rect 28001 7050 28013 7053
rect 27955 7044 28013 7050
rect 28240 7041 28246 7053
rect 28298 7041 28304 7093
rect 28642 7090 28670 7127
rect 30736 7115 30742 7167
rect 30794 7155 30800 7167
rect 31618 7155 31646 7192
rect 32944 7189 32950 7241
rect 33002 7229 33008 7241
rect 33907 7232 33965 7238
rect 33907 7229 33919 7232
rect 33002 7201 33919 7229
rect 33002 7189 33008 7201
rect 33907 7198 33919 7201
rect 33953 7198 33965 7232
rect 33907 7192 33965 7198
rect 42163 7232 42221 7238
rect 42163 7198 42175 7232
rect 42209 7198 42221 7232
rect 42163 7192 42221 7198
rect 30794 7127 31646 7155
rect 30794 7115 30800 7127
rect 35440 7115 35446 7167
rect 35498 7155 35504 7167
rect 38896 7155 38902 7167
rect 35498 7127 38558 7155
rect 38857 7127 38902 7155
rect 35498 7115 35504 7127
rect 28627 7084 28685 7090
rect 28627 7050 28639 7084
rect 28673 7050 28685 7084
rect 29488 7081 29494 7093
rect 29449 7053 29494 7081
rect 28627 7044 28685 7050
rect 29488 7041 29494 7053
rect 29546 7041 29552 7093
rect 31696 7081 31702 7093
rect 31657 7053 31702 7081
rect 31696 7041 31702 7053
rect 31754 7041 31760 7093
rect 32464 7081 32470 7093
rect 32425 7053 32470 7081
rect 32464 7041 32470 7053
rect 32522 7041 32528 7093
rect 33232 7081 33238 7093
rect 33193 7053 33238 7081
rect 33232 7041 33238 7053
rect 33290 7041 33296 7093
rect 34000 7081 34006 7093
rect 33961 7053 34006 7081
rect 34000 7041 34006 7053
rect 34058 7041 34064 7093
rect 36691 7084 36749 7090
rect 36691 7050 36703 7084
rect 36737 7081 36749 7084
rect 36880 7081 36886 7093
rect 36737 7053 36886 7081
rect 36737 7050 36749 7053
rect 36691 7044 36749 7050
rect 36880 7041 36886 7053
rect 36938 7081 36944 7093
rect 37171 7084 37229 7090
rect 37171 7081 37183 7084
rect 36938 7053 37183 7081
rect 36938 7041 36944 7053
rect 37171 7050 37183 7053
rect 37217 7050 37229 7084
rect 37171 7044 37229 7050
rect 37459 7084 37517 7090
rect 37459 7050 37471 7084
rect 37505 7081 37517 7084
rect 37648 7081 37654 7093
rect 37505 7053 37654 7081
rect 37505 7050 37517 7053
rect 37459 7044 37517 7050
rect 37648 7041 37654 7053
rect 37706 7041 37712 7093
rect 38530 7090 38558 7127
rect 38896 7115 38902 7127
rect 38954 7155 38960 7167
rect 38954 7127 39326 7155
rect 38954 7115 38960 7127
rect 39298 7090 39326 7127
rect 40624 7115 40630 7167
rect 40682 7155 40688 7167
rect 42178 7155 42206 7192
rect 40682 7127 42206 7155
rect 42274 7127 53294 7155
rect 40682 7115 40688 7127
rect 38515 7084 38573 7090
rect 38515 7050 38527 7084
rect 38561 7050 38573 7084
rect 38515 7044 38573 7050
rect 39283 7084 39341 7090
rect 39283 7050 39295 7084
rect 39329 7050 39341 7084
rect 40048 7081 40054 7093
rect 40009 7053 40054 7081
rect 39283 7044 39341 7050
rect 40048 7041 40054 7053
rect 40106 7041 40112 7093
rect 41488 7081 41494 7093
rect 41449 7053 41494 7081
rect 41488 7041 41494 7053
rect 41546 7041 41552 7093
rect 42274 7090 42302 7127
rect 42259 7084 42317 7090
rect 42259 7050 42271 7084
rect 42305 7050 42317 7084
rect 42259 7044 42317 7050
rect 42739 7084 42797 7090
rect 42739 7050 42751 7084
rect 42785 7081 42797 7084
rect 42928 7081 42934 7093
rect 42785 7053 42934 7081
rect 42785 7050 42797 7053
rect 42739 7044 42797 7050
rect 42928 7041 42934 7053
rect 42986 7041 42992 7093
rect 43120 7041 43126 7093
rect 43178 7081 43184 7093
rect 43715 7084 43773 7090
rect 43715 7081 43727 7084
rect 43178 7053 43727 7081
rect 43178 7041 43184 7053
rect 43715 7050 43727 7053
rect 43761 7050 43773 7084
rect 43715 7044 43773 7050
rect 44275 7084 44333 7090
rect 44275 7050 44287 7084
rect 44321 7081 44333 7084
rect 44560 7081 44566 7093
rect 44321 7053 44566 7081
rect 44321 7050 44333 7053
rect 44275 7044 44333 7050
rect 44560 7041 44566 7053
rect 44618 7041 44624 7093
rect 46576 7041 46582 7093
rect 46634 7081 46640 7093
rect 46771 7084 46829 7090
rect 46771 7081 46783 7084
rect 46634 7053 46783 7081
rect 46634 7041 46640 7053
rect 46771 7050 46783 7053
rect 46817 7050 46829 7084
rect 47152 7081 47158 7093
rect 47113 7053 47158 7081
rect 46771 7044 46829 7050
rect 47152 7041 47158 7053
rect 47210 7081 47216 7093
rect 47443 7084 47501 7090
rect 47443 7081 47455 7084
rect 47210 7053 47455 7081
rect 47210 7041 47216 7053
rect 47443 7050 47455 7053
rect 47489 7050 47501 7084
rect 47443 7044 47501 7050
rect 48112 7041 48118 7093
rect 48170 7081 48176 7093
rect 48307 7084 48365 7090
rect 48307 7081 48319 7084
rect 48170 7053 48319 7081
rect 48170 7041 48176 7053
rect 48307 7050 48319 7053
rect 48353 7050 48365 7084
rect 49072 7081 49078 7093
rect 49033 7053 49078 7081
rect 48307 7044 48365 7050
rect 49072 7041 49078 7053
rect 49130 7041 49136 7093
rect 49936 7041 49942 7093
rect 49994 7081 50000 7093
rect 50323 7084 50381 7090
rect 50323 7081 50335 7084
rect 49994 7053 50335 7081
rect 49994 7041 50000 7053
rect 50323 7050 50335 7053
rect 50369 7050 50381 7084
rect 52048 7081 52054 7093
rect 52009 7053 52054 7081
rect 50323 7044 50381 7050
rect 52048 7041 52054 7053
rect 52106 7041 52112 7093
rect 52432 7081 52438 7093
rect 52393 7053 52438 7081
rect 52432 7041 52438 7053
rect 52490 7081 52496 7093
rect 52723 7084 52781 7090
rect 52723 7081 52735 7084
rect 52490 7053 52735 7081
rect 52490 7041 52496 7053
rect 52723 7050 52735 7053
rect 52769 7050 52781 7084
rect 53266 7081 53294 7127
rect 56368 7115 56374 7167
rect 56426 7155 56432 7167
rect 56752 7155 56758 7167
rect 56426 7127 56758 7155
rect 56426 7115 56432 7127
rect 56752 7115 56758 7127
rect 56810 7115 56816 7167
rect 54352 7081 54358 7093
rect 53266 7053 54358 7081
rect 52723 7044 52781 7050
rect 54352 7041 54358 7053
rect 54410 7041 54416 7093
rect 1648 7007 1654 7019
rect 1609 6979 1654 7007
rect 1648 6967 1654 6979
rect 1706 6967 1712 7019
rect 2512 7007 2518 7019
rect 2473 6979 2518 7007
rect 2512 6967 2518 6979
rect 2570 6967 2576 7019
rect 4243 7010 4301 7016
rect 4243 6976 4255 7010
rect 4289 7007 4301 7010
rect 4531 7010 4589 7016
rect 4531 7007 4543 7010
rect 4289 6979 4543 7007
rect 4289 6976 4301 6979
rect 4243 6970 4301 6976
rect 4531 6976 4543 6979
rect 4577 7007 4589 7010
rect 11248 7007 11254 7019
rect 4577 6979 7214 7007
rect 11209 6979 11254 7007
rect 4577 6976 4589 6979
rect 4531 6970 4589 6976
rect 4435 6936 4493 6942
rect 4435 6902 4447 6936
rect 4481 6933 4493 6936
rect 5104 6933 5110 6945
rect 4481 6905 5110 6933
rect 4481 6902 4493 6905
rect 4435 6896 4493 6902
rect 5104 6893 5110 6905
rect 5162 6893 5168 6945
rect 5203 6936 5261 6942
rect 5203 6902 5215 6936
rect 5249 6902 5261 6936
rect 5203 6896 5261 6902
rect 5299 6936 5357 6942
rect 5299 6902 5311 6936
rect 5345 6933 5357 6936
rect 5680 6933 5686 6945
rect 5345 6905 5686 6933
rect 5345 6902 5357 6905
rect 5299 6896 5357 6902
rect 3664 6819 3670 6871
rect 3722 6859 3728 6871
rect 5218 6859 5246 6896
rect 5680 6893 5686 6905
rect 5738 6893 5744 6945
rect 5872 6893 5878 6945
rect 5930 6933 5936 6945
rect 5971 6936 6029 6942
rect 5971 6933 5983 6936
rect 5930 6905 5983 6933
rect 5930 6893 5936 6905
rect 5971 6902 5983 6905
rect 6017 6902 6029 6936
rect 5971 6896 6029 6902
rect 6067 6936 6125 6942
rect 6067 6902 6079 6936
rect 6113 6933 6125 6936
rect 6160 6933 6166 6945
rect 6113 6905 6166 6933
rect 6113 6902 6125 6905
rect 6067 6896 6125 6902
rect 3722 6831 5246 6859
rect 5779 6862 5837 6868
rect 3722 6819 3728 6831
rect 5779 6828 5791 6862
rect 5825 6859 5837 6862
rect 6082 6859 6110 6896
rect 6160 6893 6166 6905
rect 6218 6893 6224 6945
rect 6544 6893 6550 6945
rect 6602 6933 6608 6945
rect 6739 6936 6797 6942
rect 6739 6933 6751 6936
rect 6602 6905 6751 6933
rect 6602 6893 6608 6905
rect 6739 6902 6751 6905
rect 6785 6902 6797 6936
rect 6739 6896 6797 6902
rect 5825 6831 6110 6859
rect 5825 6828 5837 6831
rect 5779 6822 5837 6828
rect 7186 6785 7214 6979
rect 11248 6967 11254 6979
rect 11306 6967 11312 7019
rect 12688 7007 12694 7019
rect 12649 6979 12694 7007
rect 12688 6967 12694 6979
rect 12746 6967 12752 7019
rect 23363 7010 23421 7016
rect 12802 6979 23294 7007
rect 7312 6893 7318 6945
rect 7370 6933 7376 6945
rect 7507 6936 7565 6942
rect 7507 6933 7519 6936
rect 7370 6905 7519 6933
rect 7370 6893 7376 6905
rect 7507 6902 7519 6905
rect 7553 6902 7565 6936
rect 7507 6896 7565 6902
rect 8080 6893 8086 6945
rect 8138 6933 8144 6945
rect 8275 6936 8333 6942
rect 8275 6933 8287 6936
rect 8138 6905 8287 6933
rect 8138 6893 8144 6905
rect 8275 6902 8287 6905
rect 8321 6902 8333 6936
rect 8275 6896 8333 6902
rect 8848 6893 8854 6945
rect 8906 6933 8912 6945
rect 9715 6936 9773 6942
rect 9715 6933 9727 6936
rect 8906 6905 9727 6933
rect 8906 6893 8912 6905
rect 9715 6902 9727 6905
rect 9761 6902 9773 6936
rect 10483 6936 10541 6942
rect 10483 6933 10495 6936
rect 9715 6896 9773 6902
rect 9826 6905 10495 6933
rect 9520 6819 9526 6871
rect 9578 6859 9584 6871
rect 9826 6859 9854 6905
rect 10483 6902 10495 6905
rect 10529 6902 10541 6936
rect 10483 6896 10541 6902
rect 10579 6936 10637 6942
rect 10579 6902 10591 6936
rect 10625 6933 10637 6936
rect 12802 6933 12830 6979
rect 10625 6905 12830 6933
rect 10625 6902 10637 6905
rect 10579 6896 10637 6902
rect 9578 6831 9854 6859
rect 10291 6862 10349 6868
rect 9578 6819 9584 6831
rect 10291 6828 10303 6862
rect 10337 6859 10349 6862
rect 10594 6859 10622 6896
rect 13456 6893 13462 6945
rect 13514 6933 13520 6945
rect 13555 6936 13613 6942
rect 13555 6933 13567 6936
rect 13514 6905 13567 6933
rect 13514 6893 13520 6905
rect 13555 6902 13567 6905
rect 13601 6902 13613 6936
rect 13555 6896 13613 6902
rect 13648 6893 13654 6945
rect 13706 6933 13712 6945
rect 13706 6905 13751 6933
rect 13706 6893 13712 6905
rect 14512 6893 14518 6945
rect 14570 6933 14576 6945
rect 14995 6936 15053 6942
rect 14995 6933 15007 6936
rect 14570 6905 15007 6933
rect 14570 6893 14576 6905
rect 14995 6902 15007 6905
rect 15041 6902 15053 6936
rect 14995 6896 15053 6902
rect 15088 6893 15094 6945
rect 15146 6933 15152 6945
rect 15763 6936 15821 6942
rect 15763 6933 15775 6936
rect 15146 6905 15775 6933
rect 15146 6893 15152 6905
rect 15763 6902 15775 6905
rect 15809 6902 15821 6936
rect 17296 6933 17302 6945
rect 17257 6905 17302 6933
rect 15763 6896 15821 6902
rect 17296 6893 17302 6905
rect 17354 6893 17360 6945
rect 17872 6893 17878 6945
rect 17930 6933 17936 6945
rect 17971 6936 18029 6942
rect 17971 6933 17983 6936
rect 17930 6905 17983 6933
rect 17930 6893 17936 6905
rect 17971 6902 17983 6905
rect 18017 6902 18029 6936
rect 17971 6896 18029 6902
rect 18640 6893 18646 6945
rect 18698 6933 18704 6945
rect 18739 6936 18797 6942
rect 18739 6933 18751 6936
rect 18698 6905 18751 6933
rect 18698 6893 18704 6905
rect 18739 6902 18751 6905
rect 18785 6902 18797 6936
rect 18739 6896 18797 6902
rect 20275 6936 20333 6942
rect 20275 6902 20287 6936
rect 20321 6933 20333 6936
rect 20368 6933 20374 6945
rect 20321 6905 20374 6933
rect 20321 6902 20333 6905
rect 20275 6896 20333 6902
rect 20368 6893 20374 6905
rect 20426 6893 20432 6945
rect 20848 6893 20854 6945
rect 20906 6933 20912 6945
rect 21043 6936 21101 6942
rect 21043 6933 21055 6936
rect 20906 6905 21055 6933
rect 20906 6893 20912 6905
rect 21043 6902 21055 6905
rect 21089 6902 21101 6936
rect 21043 6896 21101 6902
rect 21232 6893 21238 6945
rect 21290 6933 21296 6945
rect 21811 6936 21869 6942
rect 21811 6933 21823 6936
rect 21290 6905 21823 6933
rect 21290 6893 21296 6905
rect 21811 6902 21823 6905
rect 21857 6902 21869 6936
rect 21811 6896 21869 6902
rect 21904 6893 21910 6945
rect 21962 6933 21968 6945
rect 22675 6936 22733 6942
rect 22675 6933 22687 6936
rect 21962 6905 22687 6933
rect 21962 6893 21968 6905
rect 22675 6902 22687 6905
rect 22721 6902 22733 6936
rect 23266 6933 23294 6979
rect 23363 6976 23375 7010
rect 23409 7007 23421 7010
rect 23632 7007 23638 7019
rect 23409 6979 23638 7007
rect 23409 6976 23421 6979
rect 23363 6970 23421 6976
rect 23632 6967 23638 6979
rect 23690 6967 23696 7019
rect 25168 6967 25174 7019
rect 25226 7007 25232 7019
rect 25226 6979 26366 7007
rect 25226 6967 25232 6979
rect 23920 6933 23926 6945
rect 23266 6905 23926 6933
rect 22675 6896 22733 6902
rect 23920 6893 23926 6905
rect 23978 6893 23984 6945
rect 24112 6933 24118 6945
rect 24073 6905 24118 6933
rect 24112 6893 24118 6905
rect 24170 6893 24176 6945
rect 24880 6893 24886 6945
rect 24938 6933 24944 6945
rect 26338 6942 26366 6979
rect 27760 6967 27766 7019
rect 27818 7007 27824 7019
rect 30931 7010 30989 7016
rect 27818 6979 28766 7007
rect 27818 6967 27824 6979
rect 25555 6936 25613 6942
rect 25555 6933 25567 6936
rect 24938 6905 25567 6933
rect 24938 6893 24944 6905
rect 25555 6902 25567 6905
rect 25601 6902 25613 6936
rect 25555 6896 25613 6902
rect 26323 6936 26381 6942
rect 26323 6902 26335 6936
rect 26369 6902 26381 6936
rect 27088 6933 27094 6945
rect 27049 6905 27094 6933
rect 26323 6896 26381 6902
rect 27088 6893 27094 6905
rect 27146 6893 27152 6945
rect 27376 6893 27382 6945
rect 27434 6933 27440 6945
rect 28738 6942 28766 6979
rect 30931 6976 30943 7010
rect 30977 7007 30989 7010
rect 32272 7007 32278 7019
rect 30977 6979 32278 7007
rect 30977 6976 30989 6979
rect 30931 6970 30989 6976
rect 32272 6967 32278 6979
rect 32330 6967 32336 7019
rect 36211 7010 36269 7016
rect 36211 6976 36223 7010
rect 36257 7007 36269 7010
rect 45616 7007 45622 7019
rect 36257 6979 45622 7007
rect 36257 6976 36269 6979
rect 36211 6970 36269 6976
rect 45616 6967 45622 6979
rect 45674 6967 45680 7019
rect 46480 6967 46486 7019
rect 46538 7007 46544 7019
rect 54067 7010 54125 7016
rect 46538 6979 48254 7007
rect 46538 6967 46544 6979
rect 27859 6936 27917 6942
rect 27859 6933 27871 6936
rect 27434 6905 27871 6933
rect 27434 6893 27440 6905
rect 27859 6902 27871 6905
rect 27905 6902 27917 6936
rect 27859 6896 27917 6902
rect 28723 6936 28781 6942
rect 28723 6902 28735 6936
rect 28769 6902 28781 6936
rect 29392 6933 29398 6945
rect 29353 6905 29398 6933
rect 28723 6896 28781 6902
rect 29392 6893 29398 6905
rect 29450 6893 29456 6945
rect 29968 6893 29974 6945
rect 30026 6933 30032 6945
rect 30835 6936 30893 6942
rect 30835 6933 30847 6936
rect 30026 6905 30847 6933
rect 30026 6893 30032 6905
rect 30835 6902 30847 6905
rect 30881 6902 30893 6936
rect 30835 6896 30893 6902
rect 31408 6893 31414 6945
rect 31466 6933 31472 6945
rect 32371 6936 32429 6942
rect 32371 6933 32383 6936
rect 31466 6905 32383 6933
rect 31466 6893 31472 6905
rect 32371 6902 32383 6905
rect 32417 6902 32429 6936
rect 32371 6896 32429 6902
rect 32464 6893 32470 6945
rect 32522 6933 32528 6945
rect 33139 6936 33197 6942
rect 33139 6933 33151 6936
rect 32522 6905 33151 6933
rect 32522 6893 32528 6905
rect 33139 6902 33151 6905
rect 33185 6902 33197 6936
rect 33139 6896 33197 6902
rect 34000 6893 34006 6945
rect 34058 6933 34064 6945
rect 34675 6936 34733 6942
rect 34675 6933 34687 6936
rect 34058 6905 34687 6933
rect 34058 6893 34064 6905
rect 34675 6902 34687 6905
rect 34721 6902 34733 6936
rect 34675 6896 34733 6902
rect 34771 6936 34829 6942
rect 34771 6902 34783 6936
rect 34817 6933 34829 6936
rect 35344 6933 35350 6945
rect 34817 6905 35350 6933
rect 34817 6902 34829 6905
rect 34771 6896 34829 6902
rect 35344 6893 35350 6905
rect 35402 6893 35408 6945
rect 35536 6893 35542 6945
rect 35594 6933 35600 6945
rect 36115 6936 36173 6942
rect 36115 6933 36127 6936
rect 35594 6905 36127 6933
rect 35594 6893 35600 6905
rect 36115 6902 36127 6905
rect 36161 6902 36173 6936
rect 36115 6896 36173 6902
rect 36496 6893 36502 6945
rect 36554 6933 36560 6945
rect 36979 6936 37037 6942
rect 36979 6933 36991 6936
rect 36554 6905 36991 6933
rect 36554 6893 36560 6905
rect 36979 6902 36991 6905
rect 37025 6902 37037 6936
rect 36979 6896 37037 6902
rect 37072 6893 37078 6945
rect 37130 6933 37136 6945
rect 37747 6936 37805 6942
rect 37747 6933 37759 6936
rect 37130 6905 37759 6933
rect 37130 6893 37136 6905
rect 37747 6902 37759 6905
rect 37793 6902 37805 6936
rect 37747 6896 37805 6902
rect 38419 6936 38477 6942
rect 38419 6902 38431 6936
rect 38465 6902 38477 6936
rect 38419 6896 38477 6902
rect 39187 6936 39245 6942
rect 39187 6902 39199 6936
rect 39233 6902 39245 6936
rect 39187 6896 39245 6902
rect 37264 6859 37270 6871
rect 10337 6831 10622 6859
rect 12946 6831 23486 6859
rect 10337 6828 10349 6831
rect 10291 6822 10349 6828
rect 12946 6785 12974 6831
rect 7186 6757 12974 6785
rect 17011 6788 17069 6794
rect 17011 6754 17023 6788
rect 17057 6785 17069 6788
rect 23056 6785 23062 6797
rect 17057 6757 23062 6785
rect 17057 6754 17069 6757
rect 17011 6748 17069 6754
rect 23056 6745 23062 6757
rect 23114 6745 23120 6797
rect 23458 6785 23486 6831
rect 23650 6831 37270 6859
rect 23650 6785 23678 6831
rect 37264 6819 37270 6831
rect 37322 6819 37328 6871
rect 37360 6819 37366 6871
rect 37418 6859 37424 6871
rect 38434 6859 38462 6896
rect 37418 6831 38462 6859
rect 37418 6819 37424 6831
rect 23458 6757 23678 6785
rect 23920 6745 23926 6797
rect 23978 6785 23984 6797
rect 34672 6785 34678 6797
rect 23978 6757 34678 6785
rect 23978 6745 23984 6757
rect 34672 6745 34678 6757
rect 34730 6745 34736 6797
rect 37648 6745 37654 6797
rect 37706 6785 37712 6797
rect 39202 6785 39230 6896
rect 39280 6893 39286 6945
rect 39338 6933 39344 6945
rect 39955 6936 40013 6942
rect 39955 6933 39967 6936
rect 39338 6905 39967 6933
rect 39338 6893 39344 6905
rect 39955 6902 39967 6905
rect 40001 6902 40013 6936
rect 39955 6896 40013 6902
rect 41395 6936 41453 6942
rect 41395 6902 41407 6936
rect 41441 6902 41453 6936
rect 41395 6896 41453 6902
rect 39856 6819 39862 6871
rect 39914 6859 39920 6871
rect 41410 6859 41438 6896
rect 41584 6893 41590 6945
rect 41642 6933 41648 6945
rect 43027 6936 43085 6942
rect 43027 6933 43039 6936
rect 41642 6905 43039 6933
rect 41642 6893 41648 6905
rect 43027 6902 43039 6905
rect 43073 6902 43085 6936
rect 43792 6933 43798 6945
rect 43753 6905 43798 6933
rect 43027 6896 43085 6902
rect 43792 6893 43798 6905
rect 43850 6893 43856 6945
rect 44467 6936 44525 6942
rect 44467 6902 44479 6936
rect 44513 6902 44525 6936
rect 44467 6896 44525 6902
rect 45235 6936 45293 6942
rect 45235 6902 45247 6936
rect 45281 6902 45293 6936
rect 45235 6896 45293 6902
rect 45331 6936 45389 6942
rect 45331 6902 45343 6936
rect 45377 6902 45389 6936
rect 45331 6896 45389 6902
rect 39914 6831 41438 6859
rect 39914 6819 39920 6831
rect 42736 6819 42742 6871
rect 42794 6859 42800 6871
rect 44482 6859 44510 6896
rect 42794 6831 44510 6859
rect 42794 6819 42800 6831
rect 37706 6757 39230 6785
rect 37706 6745 37712 6757
rect 43600 6745 43606 6797
rect 43658 6785 43664 6797
rect 45250 6785 45278 6896
rect 43658 6757 45278 6785
rect 45346 6785 45374 6896
rect 45808 6893 45814 6945
rect 45866 6933 45872 6945
rect 48226 6942 48254 6979
rect 54067 6976 54079 7010
rect 54113 6976 54125 7010
rect 54736 7007 54742 7019
rect 54697 6979 54742 7007
rect 54067 6970 54125 6976
rect 46675 6936 46733 6942
rect 46675 6933 46687 6936
rect 45866 6905 46687 6933
rect 45866 6893 45872 6905
rect 46675 6902 46687 6905
rect 46721 6902 46733 6936
rect 47539 6936 47597 6942
rect 47539 6933 47551 6936
rect 46675 6896 46733 6902
rect 46786 6905 47551 6933
rect 45712 6819 45718 6871
rect 45770 6859 45776 6871
rect 46786 6859 46814 6905
rect 47539 6902 47551 6905
rect 47585 6902 47597 6936
rect 47539 6896 47597 6902
rect 48211 6936 48269 6942
rect 48211 6902 48223 6936
rect 48257 6902 48269 6936
rect 48211 6896 48269 6902
rect 48979 6936 49037 6942
rect 48979 6902 48991 6936
rect 49025 6902 49037 6936
rect 48979 6896 49037 6902
rect 45770 6831 46814 6859
rect 45770 6819 45776 6831
rect 47248 6819 47254 6871
rect 47306 6859 47312 6871
rect 48994 6859 49022 6896
rect 50128 6893 50134 6945
rect 50186 6933 50192 6945
rect 50227 6936 50285 6942
rect 50227 6933 50239 6936
rect 50186 6905 50239 6933
rect 50186 6893 50192 6905
rect 50227 6902 50239 6905
rect 50273 6902 50285 6936
rect 50227 6896 50285 6902
rect 51280 6893 51286 6945
rect 51338 6933 51344 6945
rect 51955 6936 52013 6942
rect 51955 6933 51967 6936
rect 51338 6905 51967 6933
rect 51338 6893 51344 6905
rect 51955 6902 51967 6905
rect 52001 6902 52013 6936
rect 52816 6933 52822 6945
rect 52777 6905 52822 6933
rect 51955 6896 52013 6902
rect 52816 6893 52822 6905
rect 52874 6893 52880 6945
rect 54082 6933 54110 6970
rect 54736 6967 54742 6979
rect 54794 6967 54800 7019
rect 55408 6967 55414 7019
rect 55466 7007 55472 7019
rect 55507 7010 55565 7016
rect 55507 7007 55519 7010
rect 55466 6979 55519 7007
rect 55466 6967 55472 6979
rect 55507 6976 55519 6979
rect 55553 6976 55565 7010
rect 55507 6970 55565 6976
rect 57811 7010 57869 7016
rect 57811 6976 57823 7010
rect 57857 7007 57869 7010
rect 58480 7007 58486 7019
rect 57857 6979 58486 7007
rect 57857 6976 57869 6979
rect 57811 6970 57869 6976
rect 58480 6967 58486 6979
rect 58538 6967 58544 7019
rect 56272 6933 56278 6945
rect 54082 6905 56278 6933
rect 56272 6893 56278 6905
rect 56330 6893 56336 6945
rect 47306 6831 49022 6859
rect 47306 6819 47312 6831
rect 49168 6785 49174 6797
rect 45346 6757 49174 6785
rect 43658 6745 43664 6757
rect 49168 6745 49174 6757
rect 49226 6745 49232 6797
rect 1152 6686 58848 6708
rect 1152 6634 4294 6686
rect 4346 6634 4358 6686
rect 4410 6634 4422 6686
rect 4474 6634 4486 6686
rect 4538 6634 35014 6686
rect 35066 6634 35078 6686
rect 35130 6634 35142 6686
rect 35194 6634 35206 6686
rect 35258 6634 58848 6686
rect 1152 6612 58848 6634
rect 6160 6523 6166 6575
rect 6218 6563 6224 6575
rect 12112 6563 12118 6575
rect 6218 6535 12118 6563
rect 6218 6523 6224 6535
rect 12112 6523 12118 6535
rect 12170 6523 12176 6575
rect 18931 6566 18989 6572
rect 18931 6532 18943 6566
rect 18977 6563 18989 6566
rect 19024 6563 19030 6575
rect 18977 6535 19030 6563
rect 18977 6532 18989 6535
rect 18931 6526 18989 6532
rect 19024 6523 19030 6535
rect 19082 6523 19088 6575
rect 33136 6523 33142 6575
rect 33194 6563 33200 6575
rect 33194 6535 33239 6563
rect 33194 6523 33200 6535
rect 36688 6523 36694 6575
rect 36746 6563 36752 6575
rect 36883 6566 36941 6572
rect 36883 6563 36895 6566
rect 36746 6535 36895 6563
rect 36746 6523 36752 6535
rect 36883 6532 36895 6535
rect 36929 6532 36941 6566
rect 36883 6526 36941 6532
rect 38416 6523 38422 6575
rect 38474 6563 38480 6575
rect 39280 6563 39286 6575
rect 38474 6535 39286 6563
rect 38474 6523 38480 6535
rect 39280 6523 39286 6535
rect 39338 6523 39344 6575
rect 50611 6566 50669 6572
rect 50611 6532 50623 6566
rect 50657 6563 50669 6566
rect 50704 6563 50710 6575
rect 50657 6535 50710 6563
rect 50657 6532 50669 6535
rect 50611 6526 50669 6532
rect 50704 6523 50710 6535
rect 50762 6563 50768 6575
rect 50762 6535 50846 6563
rect 50762 6523 50768 6535
rect 8371 6492 8429 6498
rect 8371 6458 8383 6492
rect 8417 6489 8429 6492
rect 8851 6492 8909 6498
rect 8851 6489 8863 6492
rect 8417 6461 8863 6489
rect 8417 6458 8429 6461
rect 8371 6452 8429 6458
rect 8851 6458 8863 6461
rect 8897 6458 8909 6492
rect 8851 6452 8909 6458
rect 9139 6492 9197 6498
rect 9139 6458 9151 6492
rect 9185 6489 9197 6492
rect 9185 6461 33134 6489
rect 9185 6458 9197 6461
rect 9139 6452 9197 6458
rect 7120 6415 7126 6427
rect 7081 6387 7126 6415
rect 7120 6375 7126 6387
rect 7178 6375 7184 6427
rect 8464 6375 8470 6427
rect 8522 6415 8528 6427
rect 9442 6424 9470 6461
rect 9331 6418 9389 6424
rect 9331 6415 9343 6418
rect 8522 6387 9343 6415
rect 8522 6375 8528 6387
rect 9331 6384 9343 6387
rect 9377 6384 9389 6418
rect 9331 6378 9389 6384
rect 9427 6418 9485 6424
rect 9427 6384 9439 6418
rect 9473 6384 9485 6418
rect 13936 6415 13942 6427
rect 13897 6387 13942 6415
rect 9427 6378 9485 6384
rect 13936 6375 13942 6387
rect 13994 6375 14000 6427
rect 14704 6415 14710 6427
rect 14665 6387 14710 6415
rect 14704 6375 14710 6387
rect 14762 6375 14768 6427
rect 15187 6418 15245 6424
rect 15187 6384 15199 6418
rect 15233 6415 15245 6418
rect 15472 6415 15478 6427
rect 15233 6387 15478 6415
rect 15233 6384 15245 6387
rect 15187 6378 15245 6384
rect 15472 6375 15478 6387
rect 15530 6375 15536 6427
rect 16432 6415 16438 6427
rect 15586 6387 16438 6415
rect 1552 6341 1558 6353
rect 1513 6313 1558 6341
rect 1552 6301 1558 6313
rect 1610 6301 1616 6353
rect 2032 6301 2038 6353
rect 2090 6341 2096 6353
rect 2323 6344 2381 6350
rect 2323 6341 2335 6344
rect 2090 6313 2335 6341
rect 2090 6301 2096 6313
rect 2323 6310 2335 6313
rect 2369 6310 2381 6344
rect 3184 6341 3190 6353
rect 3145 6313 3190 6341
rect 2323 6304 2381 6310
rect 3184 6301 3190 6313
rect 3242 6301 3248 6353
rect 3856 6301 3862 6353
rect 3914 6341 3920 6353
rect 3955 6344 4013 6350
rect 3955 6341 3967 6344
rect 3914 6313 3967 6341
rect 3914 6301 3920 6313
rect 3955 6310 3967 6313
rect 4001 6310 4013 6344
rect 3955 6304 4013 6310
rect 4624 6301 4630 6353
rect 4682 6341 4688 6353
rect 4723 6344 4781 6350
rect 4723 6341 4735 6344
rect 4682 6313 4735 6341
rect 4682 6301 4688 6313
rect 4723 6310 4735 6313
rect 4769 6310 4781 6344
rect 4723 6304 4781 6310
rect 5683 6344 5741 6350
rect 5683 6310 5695 6344
rect 5729 6341 5741 6344
rect 8752 6341 8758 6353
rect 5729 6313 8758 6341
rect 5729 6310 5741 6313
rect 5683 6304 5741 6310
rect 8752 6301 8758 6313
rect 8810 6301 8816 6353
rect 10096 6341 10102 6353
rect 10057 6313 10102 6341
rect 10096 6301 10102 6313
rect 10154 6301 10160 6353
rect 10864 6341 10870 6353
rect 10825 6313 10870 6341
rect 10864 6301 10870 6313
rect 10922 6301 10928 6353
rect 11632 6301 11638 6353
rect 11690 6341 11696 6353
rect 12211 6344 12269 6350
rect 12211 6341 12223 6344
rect 11690 6313 12223 6341
rect 11690 6301 11696 6313
rect 12211 6310 12223 6313
rect 12257 6310 12269 6344
rect 12211 6304 12269 6310
rect 12304 6301 12310 6353
rect 12362 6341 12368 6353
rect 12979 6344 13037 6350
rect 12979 6341 12991 6344
rect 12362 6313 12991 6341
rect 12362 6301 12368 6313
rect 12979 6310 12991 6313
rect 13025 6310 13037 6344
rect 15586 6341 15614 6387
rect 16432 6375 16438 6387
rect 16490 6375 16496 6427
rect 18448 6415 18454 6427
rect 18409 6387 18454 6415
rect 18448 6375 18454 6387
rect 18506 6375 18512 6427
rect 19024 6375 19030 6427
rect 19082 6415 19088 6427
rect 19219 6418 19277 6424
rect 19219 6415 19231 6418
rect 19082 6387 19231 6415
rect 19082 6375 19088 6387
rect 19219 6384 19231 6387
rect 19265 6384 19277 6418
rect 19219 6378 19277 6384
rect 19699 6418 19757 6424
rect 19699 6384 19711 6418
rect 19745 6415 19757 6418
rect 19984 6415 19990 6427
rect 19745 6387 19990 6415
rect 19745 6384 19757 6387
rect 19699 6378 19757 6384
rect 19984 6375 19990 6387
rect 20042 6375 20048 6427
rect 20467 6418 20525 6424
rect 20467 6384 20479 6418
rect 20513 6415 20525 6418
rect 20755 6418 20813 6424
rect 20755 6415 20767 6418
rect 20513 6387 20767 6415
rect 20513 6384 20525 6387
rect 20467 6378 20525 6384
rect 20755 6384 20767 6387
rect 20801 6415 20813 6418
rect 20944 6415 20950 6427
rect 20801 6387 20950 6415
rect 20801 6384 20813 6387
rect 20755 6378 20813 6384
rect 20944 6375 20950 6387
rect 21002 6375 21008 6427
rect 21235 6418 21293 6424
rect 21235 6384 21247 6418
rect 21281 6415 21293 6418
rect 21520 6415 21526 6427
rect 21281 6387 21526 6415
rect 21281 6384 21293 6387
rect 21235 6378 21293 6384
rect 21520 6375 21526 6387
rect 21578 6375 21584 6427
rect 22675 6418 22733 6424
rect 22675 6384 22687 6418
rect 22721 6415 22733 6418
rect 22960 6415 22966 6427
rect 22721 6387 22966 6415
rect 22721 6384 22733 6387
rect 22675 6378 22733 6384
rect 22960 6375 22966 6387
rect 23018 6375 23024 6427
rect 23248 6375 23254 6427
rect 23306 6415 23312 6427
rect 23731 6418 23789 6424
rect 23731 6415 23743 6418
rect 23306 6387 23743 6415
rect 23306 6375 23312 6387
rect 23731 6384 23743 6387
rect 23777 6384 23789 6418
rect 23731 6378 23789 6384
rect 24211 6418 24269 6424
rect 24211 6384 24223 6418
rect 24257 6415 24269 6418
rect 24496 6415 24502 6427
rect 24257 6387 24502 6415
rect 24257 6384 24269 6387
rect 24211 6378 24269 6384
rect 24496 6375 24502 6387
rect 24554 6375 24560 6427
rect 27955 6418 28013 6424
rect 27955 6384 27967 6418
rect 28001 6415 28013 6418
rect 28147 6418 28205 6424
rect 28147 6415 28159 6418
rect 28001 6387 28159 6415
rect 28001 6384 28013 6387
rect 27955 6378 28013 6384
rect 28147 6384 28159 6387
rect 28193 6415 28205 6418
rect 28528 6415 28534 6427
rect 28193 6387 28534 6415
rect 28193 6384 28205 6387
rect 28147 6378 28205 6384
rect 28528 6375 28534 6387
rect 28586 6375 28592 6427
rect 28723 6418 28781 6424
rect 28723 6384 28735 6418
rect 28769 6415 28781 6418
rect 29008 6415 29014 6427
rect 28769 6387 29014 6415
rect 28769 6384 28781 6387
rect 28723 6378 28781 6384
rect 29008 6375 29014 6387
rect 29066 6375 29072 6427
rect 30640 6415 30646 6427
rect 30601 6387 30646 6415
rect 30640 6375 30646 6387
rect 30698 6375 30704 6427
rect 32080 6375 32086 6427
rect 32138 6415 32144 6427
rect 32179 6418 32237 6424
rect 32179 6415 32191 6418
rect 32138 6387 32191 6415
rect 32138 6375 32144 6387
rect 32179 6384 32191 6387
rect 32225 6384 32237 6418
rect 33106 6415 33134 6461
rect 37264 6449 37270 6501
rect 37322 6489 37328 6501
rect 42064 6489 42070 6501
rect 37322 6461 42070 6489
rect 37322 6449 37328 6461
rect 42064 6449 42070 6461
rect 42122 6449 42128 6501
rect 46960 6449 46966 6501
rect 47018 6489 47024 6501
rect 47152 6489 47158 6501
rect 47018 6461 47158 6489
rect 47018 6449 47024 6461
rect 47152 6449 47158 6461
rect 47210 6449 47216 6501
rect 47344 6415 47350 6427
rect 33106 6387 47350 6415
rect 32179 6378 32237 6384
rect 47344 6375 47350 6387
rect 47402 6375 47408 6427
rect 50818 6424 50846 6535
rect 50803 6418 50861 6424
rect 50803 6384 50815 6418
rect 50849 6384 50861 6418
rect 50803 6378 50861 6384
rect 51472 6375 51478 6427
rect 51530 6415 51536 6427
rect 51667 6418 51725 6424
rect 51667 6415 51679 6418
rect 51530 6387 51679 6415
rect 51530 6375 51536 6387
rect 51667 6384 51679 6387
rect 51713 6384 51725 6418
rect 51667 6378 51725 6384
rect 52339 6418 52397 6424
rect 52339 6384 52351 6418
rect 52385 6384 52397 6418
rect 56848 6415 56854 6427
rect 52339 6378 52397 6384
rect 53314 6387 56854 6415
rect 12979 6304 13037 6310
rect 13858 6313 15614 6341
rect 16339 6344 16397 6350
rect 7891 6270 7949 6276
rect 7891 6236 7903 6270
rect 7937 6267 7949 6270
rect 8560 6267 8566 6279
rect 7937 6239 8566 6267
rect 7937 6236 7949 6239
rect 7891 6230 7949 6236
rect 8560 6227 8566 6239
rect 8618 6227 8624 6279
rect 8659 6270 8717 6276
rect 8659 6236 8671 6270
rect 8705 6267 8717 6270
rect 8851 6270 8909 6276
rect 8851 6267 8863 6270
rect 8705 6239 8863 6267
rect 8705 6236 8717 6239
rect 8659 6230 8717 6236
rect 8851 6236 8863 6239
rect 8897 6267 8909 6270
rect 13858 6267 13886 6313
rect 16339 6310 16351 6344
rect 16385 6341 16397 6344
rect 16528 6341 16534 6353
rect 16385 6313 16534 6341
rect 16385 6310 16397 6313
rect 16339 6304 16397 6310
rect 16528 6301 16534 6313
rect 16586 6301 16592 6353
rect 25648 6341 25654 6353
rect 25609 6313 25654 6341
rect 25648 6301 25654 6313
rect 25706 6301 25712 6353
rect 26800 6341 26806 6353
rect 26761 6313 26806 6341
rect 26800 6301 26806 6313
rect 26858 6301 26864 6353
rect 29680 6341 29686 6353
rect 29641 6313 29686 6341
rect 29680 6301 29686 6313
rect 29738 6301 29744 6353
rect 31216 6341 31222 6353
rect 31177 6313 31222 6341
rect 31216 6301 31222 6313
rect 31274 6301 31280 6353
rect 32560 6301 32566 6353
rect 32618 6341 32624 6353
rect 34211 6344 34269 6350
rect 34211 6341 34223 6344
rect 32618 6313 34223 6341
rect 32618 6301 32624 6313
rect 34211 6310 34223 6313
rect 34257 6310 34269 6344
rect 36304 6341 36310 6353
rect 36265 6313 36310 6341
rect 34211 6304 34269 6310
rect 36304 6301 36310 6313
rect 36362 6301 36368 6353
rect 37251 6344 37309 6350
rect 37251 6341 37263 6344
rect 36418 6313 37263 6341
rect 17680 6267 17686 6279
rect 8897 6239 13886 6267
rect 17641 6239 17686 6267
rect 8897 6236 8909 6239
rect 8851 6230 8909 6236
rect 17680 6227 17686 6239
rect 17738 6227 17744 6279
rect 18064 6227 18070 6279
rect 18122 6267 18128 6279
rect 18122 6239 19166 6267
rect 18122 6227 18128 6239
rect 6928 6153 6934 6205
rect 6986 6193 6992 6205
rect 6986 6165 7214 6193
rect 6986 6153 6992 6165
rect 5488 6079 5494 6131
rect 5546 6119 5552 6131
rect 5587 6122 5645 6128
rect 5587 6119 5599 6122
rect 5546 6091 5599 6119
rect 5546 6079 5552 6091
rect 5587 6088 5599 6091
rect 5633 6088 5645 6122
rect 5587 6082 5645 6088
rect 6256 6079 6262 6131
rect 6314 6119 6320 6131
rect 7027 6122 7085 6128
rect 7027 6119 7039 6122
rect 6314 6091 7039 6119
rect 6314 6079 6320 6091
rect 7027 6088 7039 6091
rect 7073 6088 7085 6122
rect 7186 6119 7214 6165
rect 7984 6153 7990 6205
rect 8042 6193 8048 6205
rect 8042 6165 8606 6193
rect 8042 6153 8048 6165
rect 8578 6128 8606 6165
rect 14128 6153 14134 6205
rect 14186 6193 14192 6205
rect 14186 6165 15422 6193
rect 14186 6153 14192 6165
rect 7795 6122 7853 6128
rect 7795 6119 7807 6122
rect 7186 6091 7807 6119
rect 7027 6082 7085 6088
rect 7795 6088 7807 6091
rect 7841 6088 7853 6122
rect 7795 6082 7853 6088
rect 8563 6122 8621 6128
rect 8563 6088 8575 6122
rect 8609 6088 8621 6122
rect 8563 6082 8621 6088
rect 13264 6079 13270 6131
rect 13322 6119 13328 6131
rect 13843 6122 13901 6128
rect 13843 6119 13855 6122
rect 13322 6091 13855 6119
rect 13322 6079 13328 6091
rect 13843 6088 13855 6091
rect 13889 6088 13901 6122
rect 13843 6082 13901 6088
rect 13936 6079 13942 6131
rect 13994 6119 14000 6131
rect 15394 6128 15422 6165
rect 17488 6153 17494 6205
rect 17546 6193 17552 6205
rect 17546 6165 18398 6193
rect 17546 6153 17552 6165
rect 14611 6122 14669 6128
rect 14611 6119 14623 6122
rect 13994 6091 14623 6119
rect 13994 6079 14000 6091
rect 14611 6088 14623 6091
rect 14657 6088 14669 6122
rect 14611 6082 14669 6088
rect 15379 6122 15437 6128
rect 15379 6088 15391 6122
rect 15425 6088 15437 6122
rect 15379 6082 15437 6088
rect 16720 6079 16726 6131
rect 16778 6119 16784 6131
rect 18370 6128 18398 6165
rect 19138 6128 19166 6239
rect 33136 6227 33142 6279
rect 33194 6267 33200 6279
rect 33523 6270 33581 6276
rect 33523 6267 33535 6270
rect 33194 6239 33535 6267
rect 33194 6227 33200 6239
rect 33523 6236 33535 6239
rect 33569 6236 33581 6270
rect 34288 6267 34294 6279
rect 34249 6239 34294 6267
rect 33523 6230 33581 6236
rect 34288 6227 34294 6239
rect 34346 6227 34352 6279
rect 35059 6270 35117 6276
rect 35059 6236 35071 6270
rect 35105 6236 35117 6270
rect 35059 6230 35117 6236
rect 22288 6153 22294 6205
rect 22346 6193 22352 6205
rect 22346 6165 23054 6193
rect 22346 6153 22352 6165
rect 17587 6122 17645 6128
rect 17587 6119 17599 6122
rect 16778 6091 17599 6119
rect 16778 6079 16784 6091
rect 17587 6088 17599 6091
rect 17633 6088 17645 6122
rect 17587 6082 17645 6088
rect 18355 6122 18413 6128
rect 18355 6088 18367 6122
rect 18401 6088 18413 6122
rect 18355 6082 18413 6088
rect 19123 6122 19181 6128
rect 19123 6088 19135 6122
rect 19169 6088 19181 6122
rect 19123 6082 19181 6088
rect 19312 6079 19318 6131
rect 19370 6119 19376 6131
rect 19891 6122 19949 6128
rect 19891 6119 19903 6122
rect 19370 6091 19903 6119
rect 19370 6079 19376 6091
rect 19891 6088 19903 6091
rect 19937 6088 19949 6122
rect 19891 6082 19949 6088
rect 19984 6079 19990 6131
rect 20042 6119 20048 6131
rect 20659 6122 20717 6128
rect 20659 6119 20671 6122
rect 20042 6091 20671 6119
rect 20042 6079 20048 6091
rect 20659 6088 20671 6091
rect 20705 6088 20717 6122
rect 21424 6119 21430 6131
rect 21385 6091 21430 6119
rect 20659 6082 20717 6088
rect 21424 6079 21430 6091
rect 21482 6079 21488 6131
rect 22864 6119 22870 6131
rect 22825 6091 22870 6119
rect 22864 6079 22870 6091
rect 22922 6079 22928 6131
rect 23026 6119 23054 6165
rect 31792 6153 31798 6205
rect 31850 6193 31856 6205
rect 35074 6193 35102 6230
rect 35728 6227 35734 6279
rect 35786 6267 35792 6279
rect 36418 6267 36446 6313
rect 37251 6310 37263 6313
rect 37297 6310 37309 6344
rect 38896 6341 38902 6353
rect 38857 6313 38902 6341
rect 37251 6304 37309 6310
rect 38896 6301 38902 6313
rect 38954 6301 38960 6353
rect 40336 6341 40342 6353
rect 40297 6313 40342 6341
rect 40336 6301 40342 6313
rect 40394 6301 40400 6353
rect 41488 6341 41494 6353
rect 41449 6313 41494 6341
rect 41488 6301 41494 6313
rect 41546 6301 41552 6353
rect 41872 6301 41878 6353
rect 41930 6341 41936 6353
rect 42259 6344 42317 6350
rect 42259 6341 42271 6344
rect 41930 6313 42271 6341
rect 41930 6301 41936 6313
rect 42259 6310 42271 6313
rect 42305 6310 42317 6344
rect 42259 6304 42317 6310
rect 43312 6301 43318 6353
rect 43370 6341 43376 6353
rect 43891 6344 43949 6350
rect 43891 6341 43903 6344
rect 43370 6313 43903 6341
rect 43370 6301 43376 6313
rect 43891 6310 43903 6313
rect 43937 6310 43949 6344
rect 44752 6341 44758 6353
rect 44713 6313 44758 6341
rect 43891 6304 43949 6310
rect 44752 6301 44758 6313
rect 44810 6301 44816 6353
rect 45520 6341 45526 6353
rect 45481 6313 45526 6341
rect 45520 6301 45526 6313
rect 45578 6301 45584 6353
rect 46960 6341 46966 6353
rect 46921 6313 46966 6341
rect 46960 6301 46966 6313
rect 47018 6301 47024 6353
rect 47728 6341 47734 6353
rect 47689 6313 47734 6341
rect 47728 6301 47734 6313
rect 47786 6301 47792 6353
rect 48784 6301 48790 6353
rect 48842 6341 48848 6353
rect 49171 6344 49229 6350
rect 49171 6341 49183 6344
rect 48842 6313 49183 6341
rect 48842 6301 48848 6313
rect 49171 6310 49183 6313
rect 49217 6310 49229 6344
rect 49171 6304 49229 6310
rect 49552 6301 49558 6353
rect 49610 6341 49616 6353
rect 49939 6344 49997 6350
rect 49939 6341 49951 6344
rect 49610 6313 49951 6341
rect 49610 6301 49616 6313
rect 49939 6310 49951 6313
rect 49985 6310 49997 6344
rect 49939 6304 49997 6310
rect 51568 6301 51574 6353
rect 51626 6341 51632 6353
rect 52354 6341 52382 6378
rect 53314 6350 53342 6387
rect 56848 6375 56854 6387
rect 56906 6375 56912 6427
rect 51626 6313 52382 6341
rect 53299 6344 53357 6350
rect 51626 6301 51632 6313
rect 53299 6310 53311 6344
rect 53345 6310 53357 6344
rect 53299 6304 53357 6310
rect 53968 6301 53974 6353
rect 54026 6341 54032 6353
rect 54451 6344 54509 6350
rect 54451 6341 54463 6344
rect 54026 6313 54463 6341
rect 54026 6301 54032 6313
rect 54451 6310 54463 6313
rect 54497 6310 54509 6344
rect 54451 6304 54509 6310
rect 54640 6301 54646 6353
rect 54698 6341 54704 6353
rect 55219 6344 55277 6350
rect 55219 6341 55231 6344
rect 54698 6313 55231 6341
rect 54698 6301 54704 6313
rect 55219 6310 55231 6313
rect 55265 6310 55277 6344
rect 55219 6304 55277 6310
rect 55987 6344 56045 6350
rect 55987 6310 55999 6344
rect 56033 6310 56045 6344
rect 55987 6304 56045 6310
rect 57043 6344 57101 6350
rect 57043 6310 57055 6344
rect 57089 6310 57101 6344
rect 57043 6304 57101 6310
rect 57811 6344 57869 6350
rect 57811 6310 57823 6344
rect 57857 6341 57869 6344
rect 58096 6341 58102 6353
rect 57857 6313 58102 6341
rect 57857 6310 57869 6313
rect 57811 6304 57869 6310
rect 35786 6239 36446 6267
rect 35786 6227 35792 6239
rect 36688 6227 36694 6279
rect 36746 6267 36752 6279
rect 37171 6270 37229 6276
rect 37171 6267 37183 6270
rect 36746 6239 37183 6267
rect 36746 6227 36752 6239
rect 37171 6236 37183 6239
rect 37217 6236 37229 6270
rect 37171 6230 37229 6236
rect 51184 6227 51190 6279
rect 51242 6267 51248 6279
rect 52435 6270 52493 6276
rect 52435 6267 52447 6270
rect 51242 6239 52447 6267
rect 51242 6227 51248 6239
rect 52435 6236 52447 6239
rect 52481 6236 52493 6270
rect 52435 6230 52493 6236
rect 55120 6227 55126 6279
rect 55178 6267 55184 6279
rect 56002 6267 56030 6304
rect 55178 6239 56030 6267
rect 57058 6267 57086 6304
rect 58096 6301 58102 6313
rect 58154 6301 58160 6353
rect 58864 6267 58870 6279
rect 57058 6239 58870 6267
rect 55178 6227 55184 6239
rect 58864 6227 58870 6239
rect 58922 6227 58928 6279
rect 45328 6193 45334 6205
rect 31850 6165 33470 6193
rect 35074 6165 45334 6193
rect 31850 6153 31856 6165
rect 23635 6122 23693 6128
rect 23635 6119 23647 6122
rect 23026 6091 23647 6119
rect 23635 6088 23647 6091
rect 23681 6088 23693 6122
rect 23635 6082 23693 6088
rect 24304 6079 24310 6131
rect 24362 6119 24368 6131
rect 24403 6122 24461 6128
rect 24403 6119 24415 6122
rect 24362 6091 24415 6119
rect 24362 6079 24368 6091
rect 24403 6088 24415 6091
rect 24449 6088 24461 6122
rect 24403 6082 24461 6088
rect 27568 6079 27574 6131
rect 27626 6119 27632 6131
rect 28243 6122 28301 6128
rect 28243 6119 28255 6122
rect 27626 6091 28255 6119
rect 27626 6079 27632 6091
rect 28243 6088 28255 6091
rect 28289 6088 28301 6122
rect 28243 6082 28301 6088
rect 28915 6122 28973 6128
rect 28915 6088 28927 6122
rect 28961 6119 28973 6122
rect 29296 6119 29302 6131
rect 28961 6091 29302 6119
rect 28961 6088 28973 6091
rect 28915 6082 28973 6088
rect 29296 6079 29302 6091
rect 29354 6079 29360 6131
rect 29776 6079 29782 6131
rect 29834 6119 29840 6131
rect 30547 6122 30605 6128
rect 30547 6119 30559 6122
rect 29834 6091 30559 6119
rect 29834 6079 29840 6091
rect 30547 6088 30559 6091
rect 30593 6088 30605 6122
rect 30547 6082 30605 6088
rect 30640 6079 30646 6131
rect 30698 6119 30704 6131
rect 33442 6128 33470 6165
rect 45328 6153 45334 6165
rect 45386 6153 45392 6205
rect 32083 6122 32141 6128
rect 32083 6119 32095 6122
rect 30698 6091 32095 6119
rect 30698 6079 30704 6091
rect 32083 6088 32095 6091
rect 32129 6088 32141 6122
rect 32083 6082 32141 6088
rect 33427 6122 33485 6128
rect 33427 6088 33439 6122
rect 33473 6088 33485 6122
rect 33427 6082 33485 6088
rect 33520 6079 33526 6131
rect 33578 6119 33584 6131
rect 34963 6122 35021 6128
rect 34963 6119 34975 6122
rect 33578 6091 34975 6119
rect 33578 6079 33584 6091
rect 34963 6088 34975 6091
rect 35009 6088 35021 6122
rect 34963 6082 35021 6088
rect 49744 6079 49750 6131
rect 49802 6119 49808 6131
rect 50899 6122 50957 6128
rect 50899 6119 50911 6122
rect 49802 6091 50911 6119
rect 49802 6079 49808 6091
rect 50899 6088 50911 6091
rect 50945 6088 50957 6122
rect 50899 6082 50957 6088
rect 51088 6079 51094 6131
rect 51146 6119 51152 6131
rect 51571 6122 51629 6128
rect 51571 6119 51583 6122
rect 51146 6091 51583 6119
rect 51146 6079 51152 6091
rect 51571 6088 51583 6091
rect 51617 6088 51629 6122
rect 51571 6082 51629 6088
rect 1152 6020 58848 6042
rect 1152 5968 19654 6020
rect 19706 5968 19718 6020
rect 19770 5968 19782 6020
rect 19834 5968 19846 6020
rect 19898 5968 50374 6020
rect 50426 5968 50438 6020
rect 50490 5968 50502 6020
rect 50554 5968 50566 6020
rect 50618 5968 58848 6020
rect 1152 5946 58848 5968
rect 36208 5897 36214 5909
rect 23026 5869 36214 5897
rect 5680 5783 5686 5835
rect 5738 5823 5744 5835
rect 23026 5823 23054 5869
rect 36208 5857 36214 5869
rect 36266 5857 36272 5909
rect 54928 5857 54934 5909
rect 54986 5897 54992 5909
rect 55027 5900 55085 5906
rect 55027 5897 55039 5900
rect 54986 5869 55039 5897
rect 54986 5857 54992 5869
rect 55027 5866 55039 5869
rect 55073 5897 55085 5900
rect 55219 5900 55277 5906
rect 55219 5897 55231 5900
rect 55073 5869 55231 5897
rect 55073 5866 55085 5869
rect 55027 5860 55085 5866
rect 55219 5866 55231 5869
rect 55265 5866 55277 5900
rect 55219 5860 55277 5866
rect 5738 5795 23054 5823
rect 5738 5783 5744 5795
rect 23344 5783 23350 5835
rect 23402 5823 23408 5835
rect 24112 5823 24118 5835
rect 23402 5795 24118 5823
rect 23402 5783 23408 5795
rect 24112 5783 24118 5795
rect 24170 5783 24176 5835
rect 43024 5783 43030 5835
rect 43082 5823 43088 5835
rect 43082 5795 43200 5823
rect 43082 5783 43088 5795
rect 56272 5783 56278 5835
rect 56330 5823 56336 5835
rect 57712 5823 57718 5835
rect 56330 5795 57718 5823
rect 56330 5783 56336 5795
rect 57712 5783 57718 5795
rect 57770 5783 57776 5835
rect 6064 5749 6070 5761
rect 6025 5721 6070 5749
rect 6064 5709 6070 5721
rect 6122 5709 6128 5761
rect 7504 5709 7510 5761
rect 7562 5749 7568 5761
rect 34288 5749 34294 5761
rect 7562 5721 34294 5749
rect 7562 5709 7568 5721
rect 34288 5709 34294 5721
rect 34346 5709 34352 5761
rect 1072 5635 1078 5687
rect 1130 5675 1136 5687
rect 1555 5678 1613 5684
rect 1555 5675 1567 5678
rect 1130 5647 1567 5675
rect 1130 5635 1136 5647
rect 1555 5644 1567 5647
rect 1601 5644 1613 5678
rect 2896 5675 2902 5687
rect 2857 5647 2902 5675
rect 1555 5638 1613 5644
rect 2896 5635 2902 5647
rect 2954 5635 2960 5687
rect 4435 5678 4493 5684
rect 4435 5644 4447 5678
rect 4481 5675 4493 5678
rect 4912 5675 4918 5687
rect 4481 5647 4918 5675
rect 4481 5644 4493 5647
rect 4435 5638 4493 5644
rect 4912 5635 4918 5647
rect 4970 5635 4976 5687
rect 5104 5675 5110 5687
rect 5065 5647 5110 5675
rect 5104 5635 5110 5647
rect 5162 5635 5168 5687
rect 7216 5635 7222 5687
rect 7274 5675 7280 5687
rect 7274 5647 7319 5675
rect 7274 5635 7280 5647
rect 7888 5635 7894 5687
rect 7946 5675 7952 5687
rect 7987 5678 8045 5684
rect 7987 5675 7999 5678
rect 7946 5647 7999 5675
rect 7946 5635 7952 5647
rect 7987 5644 7999 5647
rect 8033 5644 8045 5678
rect 7987 5638 8045 5644
rect 9040 5635 9046 5687
rect 9098 5675 9104 5687
rect 9619 5678 9677 5684
rect 9619 5675 9631 5678
rect 9098 5647 9631 5675
rect 9098 5635 9104 5647
rect 9619 5644 9631 5647
rect 9665 5644 9677 5678
rect 9619 5638 9677 5644
rect 10192 5635 10198 5687
rect 10250 5675 10256 5687
rect 10387 5678 10445 5684
rect 10387 5675 10399 5678
rect 10250 5647 10399 5675
rect 10250 5635 10256 5647
rect 10387 5644 10399 5647
rect 10433 5644 10445 5678
rect 10387 5638 10445 5644
rect 10480 5635 10486 5687
rect 10538 5675 10544 5687
rect 11155 5678 11213 5684
rect 11155 5675 11167 5678
rect 10538 5647 11167 5675
rect 10538 5635 10544 5647
rect 11155 5644 11167 5647
rect 11201 5644 11213 5678
rect 12592 5675 12598 5687
rect 12553 5647 12598 5675
rect 11155 5638 11213 5644
rect 12592 5635 12598 5647
rect 12650 5635 12656 5687
rect 13360 5675 13366 5687
rect 13321 5647 13366 5675
rect 13360 5635 13366 5647
rect 13418 5635 13424 5687
rect 14992 5675 14998 5687
rect 14953 5647 14998 5675
rect 14992 5635 14998 5647
rect 15050 5635 15056 5687
rect 15856 5675 15862 5687
rect 15817 5647 15862 5675
rect 15856 5635 15862 5647
rect 15914 5635 15920 5687
rect 16144 5635 16150 5687
rect 16202 5675 16208 5687
rect 16531 5678 16589 5684
rect 16531 5675 16543 5678
rect 16202 5647 16543 5675
rect 16202 5635 16208 5647
rect 16531 5644 16543 5647
rect 16577 5644 16589 5678
rect 17968 5675 17974 5687
rect 17929 5647 17974 5675
rect 16531 5638 16589 5644
rect 17968 5635 17974 5647
rect 18026 5635 18032 5687
rect 18736 5675 18742 5687
rect 18697 5647 18742 5675
rect 18736 5635 18742 5647
rect 18794 5635 18800 5687
rect 20176 5675 20182 5687
rect 20137 5647 20182 5675
rect 20176 5635 20182 5647
rect 20234 5635 20240 5687
rect 20464 5635 20470 5687
rect 20522 5675 20528 5687
rect 20947 5678 21005 5684
rect 20947 5675 20959 5678
rect 20522 5647 20959 5675
rect 20522 5635 20528 5647
rect 20947 5644 20959 5647
rect 20993 5644 21005 5678
rect 21712 5675 21718 5687
rect 21673 5647 21718 5675
rect 20947 5638 21005 5644
rect 21712 5635 21718 5647
rect 21770 5635 21776 5687
rect 22480 5675 22486 5687
rect 22441 5647 22486 5675
rect 22480 5635 22486 5647
rect 22538 5635 22544 5687
rect 23056 5635 23062 5687
rect 23114 5675 23120 5687
rect 23251 5678 23309 5684
rect 23251 5675 23263 5678
rect 23114 5647 23263 5675
rect 23114 5635 23120 5647
rect 23251 5644 23263 5647
rect 23297 5644 23309 5678
rect 23251 5638 23309 5644
rect 23440 5635 23446 5687
rect 23498 5675 23504 5687
rect 24019 5678 24077 5684
rect 24019 5675 24031 5678
rect 23498 5647 24031 5675
rect 23498 5635 23504 5647
rect 24019 5644 24031 5647
rect 24065 5644 24077 5678
rect 24019 5638 24077 5644
rect 24592 5635 24598 5687
rect 24650 5675 24656 5687
rect 25459 5678 25517 5684
rect 25459 5675 25471 5678
rect 24650 5647 25471 5675
rect 24650 5635 24656 5647
rect 25459 5644 25471 5647
rect 25505 5644 25517 5678
rect 26224 5675 26230 5687
rect 26185 5647 26230 5675
rect 25459 5638 25517 5644
rect 26224 5635 26230 5647
rect 26282 5635 26288 5687
rect 26995 5678 27053 5684
rect 26995 5644 27007 5678
rect 27041 5644 27053 5678
rect 26995 5638 27053 5644
rect 5968 5601 5974 5613
rect 5929 5573 5974 5601
rect 5968 5561 5974 5573
rect 6026 5561 6032 5613
rect 26032 5561 26038 5613
rect 26090 5601 26096 5613
rect 27010 5601 27038 5638
rect 27184 5635 27190 5687
rect 27242 5675 27248 5687
rect 27763 5678 27821 5684
rect 27763 5675 27775 5678
rect 27242 5647 27775 5675
rect 27242 5635 27248 5647
rect 27763 5644 27775 5647
rect 27809 5644 27821 5678
rect 27763 5638 27821 5644
rect 27856 5635 27862 5687
rect 27914 5675 27920 5687
rect 28531 5678 28589 5684
rect 28531 5675 28543 5678
rect 27914 5647 28543 5675
rect 27914 5635 27920 5647
rect 28531 5644 28543 5647
rect 28577 5644 28589 5678
rect 28531 5638 28589 5644
rect 28816 5635 28822 5687
rect 28874 5675 28880 5687
rect 29299 5678 29357 5684
rect 29299 5675 29311 5678
rect 28874 5647 29311 5675
rect 28874 5635 28880 5647
rect 29299 5644 29311 5647
rect 29345 5644 29357 5678
rect 29299 5638 29357 5644
rect 30256 5635 30262 5687
rect 30314 5675 30320 5687
rect 30739 5678 30797 5684
rect 30739 5675 30751 5678
rect 30314 5647 30751 5675
rect 30314 5635 30320 5647
rect 30739 5644 30751 5647
rect 30785 5644 30797 5678
rect 30739 5638 30797 5644
rect 30832 5635 30838 5687
rect 30890 5675 30896 5687
rect 31507 5678 31565 5684
rect 31507 5675 31519 5678
rect 30890 5647 31519 5675
rect 30890 5635 30896 5647
rect 31507 5644 31519 5647
rect 31553 5644 31565 5678
rect 31507 5638 31565 5644
rect 31696 5635 31702 5687
rect 31754 5675 31760 5687
rect 32275 5678 32333 5684
rect 32275 5675 32287 5678
rect 31754 5647 32287 5675
rect 31754 5635 31760 5647
rect 32275 5644 32287 5647
rect 32321 5644 32333 5678
rect 32275 5638 32333 5644
rect 33136 5635 33142 5687
rect 33194 5675 33200 5687
rect 33811 5678 33869 5684
rect 33194 5647 33239 5675
rect 33194 5635 33200 5647
rect 33811 5644 33823 5678
rect 33857 5644 33869 5678
rect 34672 5675 34678 5687
rect 34633 5647 34678 5675
rect 33811 5638 33869 5644
rect 26090 5573 27038 5601
rect 26090 5561 26096 5573
rect 33232 5561 33238 5613
rect 33290 5601 33296 5613
rect 33826 5601 33854 5638
rect 34672 5635 34678 5647
rect 34730 5635 34736 5687
rect 36115 5678 36173 5684
rect 36115 5644 36127 5678
rect 36161 5675 36173 5678
rect 36208 5675 36214 5687
rect 36161 5647 36214 5675
rect 36161 5644 36173 5647
rect 36115 5638 36173 5644
rect 36208 5635 36214 5647
rect 36266 5635 36272 5687
rect 36400 5635 36406 5687
rect 36458 5675 36464 5687
rect 36787 5678 36845 5684
rect 36787 5675 36799 5678
rect 36458 5647 36799 5675
rect 36458 5635 36464 5647
rect 36787 5644 36799 5647
rect 36833 5644 36845 5678
rect 37552 5675 37558 5687
rect 37513 5647 37558 5675
rect 36787 5638 36845 5644
rect 37552 5635 37558 5647
rect 37610 5635 37616 5687
rect 38323 5678 38381 5684
rect 38323 5644 38335 5678
rect 38369 5644 38381 5678
rect 39088 5675 39094 5687
rect 39049 5647 39094 5675
rect 38323 5638 38381 5644
rect 33290 5573 33854 5601
rect 33290 5561 33296 5573
rect 37456 5561 37462 5613
rect 37514 5601 37520 5613
rect 38338 5601 38366 5638
rect 39088 5635 39094 5647
rect 39146 5635 39152 5687
rect 39280 5635 39286 5687
rect 39338 5675 39344 5687
rect 39859 5678 39917 5684
rect 39859 5675 39871 5678
rect 39338 5647 39871 5675
rect 39338 5635 39344 5647
rect 39859 5644 39871 5647
rect 39905 5644 39917 5678
rect 39859 5638 39917 5644
rect 40720 5635 40726 5687
rect 40778 5675 40784 5687
rect 41299 5678 41357 5684
rect 41299 5675 41311 5678
rect 40778 5647 41311 5675
rect 40778 5635 40784 5647
rect 41299 5644 41311 5647
rect 41345 5644 41357 5678
rect 41299 5638 41357 5644
rect 42598 5650 42650 5656
rect 37514 5573 38366 5601
rect 42598 5592 42650 5598
rect 42886 5650 42938 5656
rect 43504 5635 43510 5687
rect 43562 5675 43568 5687
rect 43891 5678 43949 5684
rect 43891 5675 43903 5678
rect 43562 5647 43903 5675
rect 43562 5635 43568 5647
rect 43891 5644 43903 5647
rect 43937 5644 43949 5678
rect 44656 5675 44662 5687
rect 44617 5647 44662 5675
rect 43891 5638 43949 5644
rect 44656 5635 44662 5647
rect 44714 5635 44720 5687
rect 46096 5635 46102 5687
rect 46154 5675 46160 5687
rect 46579 5678 46637 5684
rect 46579 5675 46591 5678
rect 46154 5647 46591 5675
rect 46154 5635 46160 5647
rect 46579 5644 46591 5647
rect 46625 5644 46637 5678
rect 46579 5638 46637 5644
rect 46672 5635 46678 5687
rect 46730 5675 46736 5687
rect 47347 5678 47405 5684
rect 47347 5675 47359 5678
rect 46730 5647 47359 5675
rect 46730 5635 46736 5647
rect 47347 5644 47359 5647
rect 47393 5644 47405 5678
rect 47347 5638 47405 5644
rect 47536 5635 47542 5687
rect 47594 5675 47600 5687
rect 48115 5678 48173 5684
rect 48115 5675 48127 5678
rect 47594 5647 48127 5675
rect 47594 5635 47600 5647
rect 48115 5644 48127 5647
rect 48161 5644 48173 5678
rect 48976 5675 48982 5687
rect 48937 5647 48982 5675
rect 48115 5638 48173 5644
rect 48976 5635 48982 5647
rect 49034 5635 49040 5687
rect 49648 5675 49654 5687
rect 49609 5647 49654 5675
rect 49648 5635 49654 5647
rect 49706 5635 49712 5687
rect 50515 5678 50573 5684
rect 50515 5644 50527 5678
rect 50561 5675 50573 5678
rect 50704 5675 50710 5687
rect 50561 5647 50710 5675
rect 50561 5644 50573 5647
rect 50515 5638 50573 5644
rect 50704 5635 50710 5647
rect 50762 5635 50768 5687
rect 52144 5675 52150 5687
rect 52105 5647 52150 5675
rect 52144 5635 52150 5647
rect 52202 5635 52208 5687
rect 52528 5635 52534 5687
rect 52586 5675 52592 5687
rect 52915 5678 52973 5684
rect 52915 5675 52927 5678
rect 52586 5647 52927 5675
rect 52586 5635 52592 5647
rect 52915 5644 52927 5647
rect 52961 5644 52973 5678
rect 53680 5675 53686 5687
rect 53641 5647 53686 5675
rect 52915 5638 52973 5644
rect 53680 5635 53686 5647
rect 53738 5635 53744 5687
rect 54451 5678 54509 5684
rect 54451 5644 54463 5678
rect 54497 5644 54509 5678
rect 54451 5638 54509 5644
rect 55987 5678 56045 5684
rect 55987 5644 55999 5678
rect 56033 5644 56045 5678
rect 57424 5675 57430 5687
rect 57385 5647 57430 5675
rect 55987 5638 56045 5644
rect 42886 5592 42938 5598
rect 37514 5561 37520 5573
rect 53584 5561 53590 5613
rect 53642 5601 53648 5613
rect 54466 5601 54494 5638
rect 53642 5573 54494 5601
rect 56002 5601 56030 5638
rect 57424 5635 57430 5647
rect 57482 5635 57488 5687
rect 59632 5601 59638 5613
rect 56002 5573 59638 5601
rect 53642 5561 53648 5573
rect 59632 5561 59638 5573
rect 59690 5561 59696 5613
rect 17680 5487 17686 5539
rect 17738 5527 17744 5539
rect 17738 5499 42480 5527
rect 17738 5487 17744 5499
rect 11827 5456 11885 5462
rect 11827 5422 11839 5456
rect 11873 5453 11885 5456
rect 12112 5453 12118 5465
rect 11873 5425 12118 5453
rect 11873 5422 11885 5425
rect 11827 5416 11885 5422
rect 12112 5413 12118 5425
rect 12170 5413 12176 5465
rect 17203 5456 17261 5462
rect 17203 5422 17215 5456
rect 17249 5453 17261 5456
rect 17491 5456 17549 5462
rect 17491 5453 17503 5456
rect 17249 5425 17503 5453
rect 17249 5422 17261 5425
rect 17203 5416 17261 5422
rect 17491 5422 17503 5425
rect 17537 5453 17549 5456
rect 28432 5453 28438 5465
rect 17537 5425 28438 5453
rect 17537 5422 17549 5425
rect 17491 5416 17549 5422
rect 28432 5413 28438 5425
rect 28490 5413 28496 5465
rect 37840 5413 37846 5465
rect 37898 5453 37904 5465
rect 42592 5453 42598 5465
rect 37898 5425 42598 5453
rect 37898 5413 37904 5425
rect 42592 5413 42598 5425
rect 42650 5413 42656 5465
rect 1152 5354 58848 5376
rect 1152 5302 4294 5354
rect 4346 5302 4358 5354
rect 4410 5302 4422 5354
rect 4474 5302 4486 5354
rect 4538 5302 35014 5354
rect 35066 5302 35078 5354
rect 35130 5302 35142 5354
rect 35194 5302 35206 5354
rect 35258 5302 58848 5354
rect 1152 5280 58848 5302
rect 18352 5191 18358 5243
rect 18410 5231 18416 5243
rect 43792 5231 43798 5243
rect 18410 5203 43798 5231
rect 18410 5191 18416 5203
rect 43792 5191 43798 5203
rect 43850 5191 43856 5243
rect 59248 5157 59254 5169
rect 55618 5129 59254 5157
rect 12112 5043 12118 5095
rect 12170 5083 12176 5095
rect 47056 5083 47062 5095
rect 12170 5055 47062 5083
rect 12170 5043 12176 5055
rect 47056 5043 47062 5055
rect 47114 5043 47120 5095
rect 304 4969 310 5021
rect 362 5009 368 5021
rect 1555 5012 1613 5018
rect 1555 5009 1567 5012
rect 362 4981 1567 5009
rect 362 4969 368 4981
rect 1555 4978 1567 4981
rect 1601 4978 1613 5012
rect 1555 4972 1613 4978
rect 1840 4969 1846 5021
rect 1898 5009 1904 5021
rect 2323 5012 2381 5018
rect 2323 5009 2335 5012
rect 1898 4981 2335 5009
rect 1898 4969 1904 4981
rect 2323 4978 2335 4981
rect 2369 4978 2381 5012
rect 3088 5009 3094 5021
rect 3049 4981 3094 5009
rect 2323 4972 2381 4978
rect 3088 4969 3094 4981
rect 3146 4969 3152 5021
rect 4144 5009 4150 5021
rect 4105 4981 4150 5009
rect 4144 4969 4150 4981
rect 4202 4969 4208 5021
rect 5392 5009 5398 5021
rect 5353 4981 5398 5009
rect 5392 4969 5398 4981
rect 5450 4969 5456 5021
rect 6064 4969 6070 5021
rect 6122 5009 6128 5021
rect 6931 5012 6989 5018
rect 6931 5009 6943 5012
rect 6122 4981 6943 5009
rect 6122 4969 6128 4981
rect 6931 4978 6943 4981
rect 6977 4978 6989 5012
rect 7696 5009 7702 5021
rect 7657 4981 7702 5009
rect 6931 4972 6989 4978
rect 7696 4969 7702 4981
rect 7754 4969 7760 5021
rect 8467 5012 8525 5018
rect 8467 4978 8479 5012
rect 8513 4978 8525 5012
rect 9232 5009 9238 5021
rect 9193 4981 9238 5009
rect 8467 4972 8525 4978
rect 7600 4895 7606 4947
rect 7658 4935 7664 4947
rect 8482 4935 8510 4972
rect 9232 4969 9238 4981
rect 9290 4969 9296 5021
rect 10099 5012 10157 5018
rect 10099 4978 10111 5012
rect 10145 5009 10157 5012
rect 10288 5009 10294 5021
rect 10145 4981 10294 5009
rect 10145 4978 10157 4981
rect 10099 4972 10157 4978
rect 10288 4969 10294 4981
rect 10346 4969 10352 5021
rect 10672 4969 10678 5021
rect 10730 5009 10736 5021
rect 10771 5012 10829 5018
rect 10771 5009 10783 5012
rect 10730 4981 10783 5009
rect 10730 4969 10736 4981
rect 10771 4978 10783 4981
rect 10817 4978 10829 5012
rect 10771 4972 10829 4978
rect 11824 4969 11830 5021
rect 11882 5009 11888 5021
rect 12211 5012 12269 5018
rect 12211 5009 12223 5012
rect 11882 4981 12223 5009
rect 11882 4969 11888 4981
rect 12211 4978 12223 4981
rect 12257 4978 12269 5012
rect 12211 4972 12269 4978
rect 12976 4969 12982 5021
rect 13034 5009 13040 5021
rect 13936 5009 13942 5021
rect 13034 4981 13079 5009
rect 13897 4981 13942 5009
rect 13034 4969 13040 4981
rect 13936 4969 13942 4981
rect 13994 4969 14000 5021
rect 14416 4969 14422 5021
rect 14474 5009 14480 5021
rect 14707 5012 14765 5018
rect 14707 5009 14719 5012
rect 14474 4981 14719 5009
rect 14474 4969 14480 4981
rect 14707 4978 14719 4981
rect 14753 4978 14765 5012
rect 14707 4972 14765 4978
rect 14800 4969 14806 5021
rect 14858 5009 14864 5021
rect 15475 5012 15533 5018
rect 15475 5009 15487 5012
rect 14858 4981 15487 5009
rect 14858 4969 14864 4981
rect 15475 4978 15487 4981
rect 15521 4978 15533 5012
rect 15475 4972 15533 4978
rect 16339 5012 16397 5018
rect 16339 4978 16351 5012
rect 16385 5009 16397 5012
rect 16432 5009 16438 5021
rect 16385 4981 16438 5009
rect 16385 4978 16397 4981
rect 16339 4972 16397 4978
rect 16432 4969 16438 4981
rect 16490 4969 16496 5021
rect 17296 4969 17302 5021
rect 17354 5009 17360 5021
rect 17491 5012 17549 5018
rect 17491 5009 17503 5012
rect 17354 4981 17503 5009
rect 17354 4969 17360 4981
rect 17491 4978 17503 4981
rect 17537 4978 17549 5012
rect 17491 4972 17549 4978
rect 17584 4969 17590 5021
rect 17642 5009 17648 5021
rect 18259 5012 18317 5018
rect 18259 5009 18271 5012
rect 17642 4981 18271 5009
rect 17642 4969 17648 4981
rect 18259 4978 18271 4981
rect 18305 4978 18317 5012
rect 19024 5009 19030 5021
rect 18985 4981 19030 5009
rect 18259 4972 18317 4978
rect 19024 4969 19030 4981
rect 19082 4969 19088 5021
rect 19216 4969 19222 5021
rect 19274 5009 19280 5021
rect 19795 5012 19853 5018
rect 19795 5009 19807 5012
rect 19274 4981 19807 5009
rect 19274 4969 19280 4981
rect 19795 4978 19807 4981
rect 19841 4978 19853 5012
rect 20560 5009 20566 5021
rect 20521 4981 20566 5009
rect 19795 4972 19853 4978
rect 20560 4969 20566 4981
rect 20618 4969 20624 5021
rect 21232 4969 21238 5021
rect 21290 5009 21296 5021
rect 21331 5012 21389 5018
rect 21331 5009 21343 5012
rect 21290 4981 21343 5009
rect 21290 4969 21296 4981
rect 21331 4978 21343 4981
rect 21377 4978 21389 5012
rect 22768 5009 22774 5021
rect 22729 4981 22774 5009
rect 21331 4972 21389 4978
rect 22768 4969 22774 4981
rect 22826 4969 22832 5021
rect 23152 4969 23158 5021
rect 23210 5009 23216 5021
rect 23539 5012 23597 5018
rect 23539 5009 23551 5012
rect 23210 4981 23551 5009
rect 23210 4969 23216 4981
rect 23539 4978 23551 4981
rect 23585 4978 23597 5012
rect 23539 4972 23597 4978
rect 23824 4969 23830 5021
rect 23882 5009 23888 5021
rect 24307 5012 24365 5018
rect 24307 5009 24319 5012
rect 23882 4981 24319 5009
rect 23882 4969 23888 4981
rect 24307 4978 24319 4981
rect 24353 4978 24365 5012
rect 24307 4972 24365 4978
rect 24400 4969 24406 5021
rect 24458 5009 24464 5021
rect 25075 5012 25133 5018
rect 25075 5009 25087 5012
rect 24458 4981 25087 5009
rect 24458 4969 24464 4981
rect 25075 4978 25087 4981
rect 25121 4978 25133 5012
rect 25840 5009 25846 5021
rect 25801 4981 25846 5009
rect 25075 4972 25133 4978
rect 25840 4969 25846 4981
rect 25898 4969 25904 5021
rect 26608 5009 26614 5021
rect 26569 4981 26614 5009
rect 26608 4969 26614 4981
rect 26666 4969 26672 5021
rect 27379 5012 27437 5018
rect 27379 4978 27391 5012
rect 27425 5009 27437 5012
rect 28051 5012 28109 5018
rect 28051 5009 28063 5012
rect 27425 4981 28063 5009
rect 27425 4978 27437 4981
rect 27379 4972 27437 4978
rect 28051 4978 28063 4981
rect 28097 4978 28109 5012
rect 28912 5009 28918 5021
rect 28873 4981 28918 5009
rect 28051 4972 28109 4978
rect 28912 4969 28918 4981
rect 28970 4969 28976 5021
rect 29008 4969 29014 5021
rect 29066 5009 29072 5021
rect 29587 5012 29645 5018
rect 29587 5009 29599 5012
rect 29066 4981 29599 5009
rect 29066 4969 29072 4981
rect 29587 4978 29599 4981
rect 29633 4978 29645 5012
rect 30352 5009 30358 5021
rect 30313 4981 30358 5009
rect 29587 4972 29645 4978
rect 30352 4969 30358 4981
rect 30410 4969 30416 5021
rect 31120 5009 31126 5021
rect 31081 4981 31126 5009
rect 31120 4969 31126 4981
rect 31178 4969 31184 5021
rect 31888 5009 31894 5021
rect 31849 4981 31894 5009
rect 31888 4969 31894 4981
rect 31946 4969 31952 5021
rect 33328 5009 33334 5021
rect 33289 4981 33334 5009
rect 33328 4969 33334 4981
rect 33386 4969 33392 5021
rect 33424 4969 33430 5021
rect 33482 5009 33488 5021
rect 34099 5012 34157 5018
rect 34099 5009 34111 5012
rect 33482 4981 34111 5009
rect 33482 4969 33488 4981
rect 34099 4978 34111 4981
rect 34145 4978 34157 5012
rect 34864 5009 34870 5021
rect 34825 4981 34870 5009
rect 34099 4972 34157 4978
rect 34864 4969 34870 4981
rect 34922 4969 34928 5021
rect 35632 5009 35638 5021
rect 35593 4981 35638 5009
rect 35632 4969 35638 4981
rect 35690 4969 35696 5021
rect 36112 4969 36118 5021
rect 36170 5009 36176 5021
rect 36403 5012 36461 5018
rect 36403 5009 36415 5012
rect 36170 4981 36415 5009
rect 36170 4969 36176 4981
rect 36403 4978 36415 4981
rect 36449 4978 36461 5012
rect 36403 4972 36461 4978
rect 36880 4969 36886 5021
rect 36938 5009 36944 5021
rect 37171 5012 37229 5018
rect 37171 5009 37183 5012
rect 36938 4981 37183 5009
rect 36938 4969 36944 4981
rect 37171 4978 37183 4981
rect 37217 4978 37229 5012
rect 38608 5009 38614 5021
rect 38569 4981 38614 5009
rect 37171 4972 37229 4978
rect 38608 4969 38614 4981
rect 38666 4969 38672 5021
rect 39376 5009 39382 5021
rect 39337 4981 39382 5009
rect 39376 4969 39382 4981
rect 39434 4969 39440 5021
rect 40144 5009 40150 5021
rect 40105 4981 40150 5009
rect 40144 4969 40150 4981
rect 40202 4969 40208 5021
rect 40912 5009 40918 5021
rect 40873 4981 40918 5009
rect 40912 4969 40918 4981
rect 40970 4969 40976 5021
rect 41296 4969 41302 5021
rect 41354 5009 41360 5021
rect 41683 5012 41741 5018
rect 41683 5009 41695 5012
rect 41354 4981 41695 5009
rect 41354 4969 41360 4981
rect 41683 4978 41695 4981
rect 41729 4978 41741 5012
rect 42448 5009 42454 5021
rect 42409 4981 42454 5009
rect 41683 4972 41741 4978
rect 42448 4969 42454 4981
rect 42506 4969 42512 5021
rect 43888 5009 43894 5021
rect 43849 4981 43894 5009
rect 43888 4969 43894 4981
rect 43946 4969 43952 5021
rect 43984 4969 43990 5021
rect 44042 5009 44048 5021
rect 44659 5012 44717 5018
rect 44659 5009 44671 5012
rect 44042 4981 44671 5009
rect 44042 4969 44048 4981
rect 44659 4978 44671 4981
rect 44705 4978 44717 5012
rect 44659 4972 44717 4978
rect 44848 4969 44854 5021
rect 44906 5009 44912 5021
rect 45427 5012 45485 5018
rect 45427 5009 45439 5012
rect 44906 4981 45439 5009
rect 44906 4969 44912 4981
rect 45427 4978 45439 4981
rect 45473 4978 45485 5012
rect 45427 4972 45485 4978
rect 45616 4969 45622 5021
rect 45674 5009 45680 5021
rect 46195 5012 46253 5018
rect 46195 5009 46207 5012
rect 45674 4981 46207 5009
rect 45674 4969 45680 4981
rect 46195 4978 46207 4981
rect 46241 4978 46253 5012
rect 46195 4972 46253 4978
rect 46480 4969 46486 5021
rect 46538 5009 46544 5021
rect 46963 5012 47021 5018
rect 46963 5009 46975 5012
rect 46538 4981 46975 5009
rect 46538 4969 46544 4981
rect 46963 4978 46975 4981
rect 47009 4978 47021 5012
rect 46963 4972 47021 4978
rect 47827 5012 47885 5018
rect 47827 4978 47839 5012
rect 47873 5009 47885 5012
rect 47920 5009 47926 5021
rect 47873 4981 47926 5009
rect 47873 4978 47885 4981
rect 47827 4972 47885 4978
rect 47920 4969 47926 4981
rect 47978 4969 47984 5021
rect 49360 5009 49366 5021
rect 49321 4981 49366 5009
rect 49360 4969 49366 4981
rect 49418 4969 49424 5021
rect 50416 5009 50422 5021
rect 50377 4981 50422 5009
rect 50416 4969 50422 4981
rect 50474 4969 50480 5021
rect 50896 4969 50902 5021
rect 50954 5009 50960 5021
rect 51091 5012 51149 5018
rect 51091 5009 51103 5012
rect 50954 4981 51103 5009
rect 50954 4969 50960 4981
rect 51091 4978 51103 4981
rect 51137 4978 51149 5012
rect 51856 5009 51862 5021
rect 51817 4981 51862 5009
rect 51091 4972 51149 4978
rect 51856 4969 51862 4981
rect 51914 4969 51920 5021
rect 51952 4969 51958 5021
rect 52010 5009 52016 5021
rect 52627 5012 52685 5018
rect 52627 5009 52639 5012
rect 52010 4981 52639 5009
rect 52010 4969 52016 4981
rect 52627 4978 52639 4981
rect 52673 4978 52685 5012
rect 52627 4972 52685 4978
rect 53296 4969 53302 5021
rect 53354 5009 53360 5021
rect 55618 5018 55646 5129
rect 59248 5117 59254 5129
rect 59306 5117 59312 5169
rect 57808 5083 57814 5095
rect 56386 5055 57814 5083
rect 56386 5018 56414 5055
rect 57808 5043 57814 5055
rect 57866 5043 57872 5095
rect 54451 5012 54509 5018
rect 54451 5009 54463 5012
rect 53354 4981 54463 5009
rect 53354 4969 53360 4981
rect 54451 4978 54463 4981
rect 54497 4978 54509 5012
rect 54451 4972 54509 4978
rect 55603 5012 55661 5018
rect 55603 4978 55615 5012
rect 55649 4978 55661 5012
rect 55603 4972 55661 4978
rect 56371 5012 56429 5018
rect 56371 4978 56383 5012
rect 56417 4978 56429 5012
rect 57040 5009 57046 5021
rect 57001 4981 57046 5009
rect 56371 4972 56429 4978
rect 57040 4969 57046 4981
rect 57098 4969 57104 5021
rect 58003 4938 58061 4944
rect 58003 4935 58015 4938
rect 7658 4907 8510 4935
rect 12946 4907 58015 4935
rect 7658 4895 7664 4907
rect 8560 4821 8566 4873
rect 8618 4861 8624 4873
rect 12946 4861 12974 4907
rect 58003 4904 58015 4907
rect 58049 4904 58061 4938
rect 58003 4898 58061 4904
rect 8618 4833 12974 4861
rect 8618 4821 8624 4833
rect 26416 4821 26422 4873
rect 26474 4861 26480 4873
rect 27379 4864 27437 4870
rect 27379 4861 27391 4864
rect 26474 4833 27391 4861
rect 26474 4821 26480 4833
rect 27379 4830 27391 4833
rect 27425 4830 27437 4864
rect 27379 4824 27437 4830
rect 15760 4747 15766 4799
rect 15818 4787 15824 4799
rect 37840 4787 37846 4799
rect 15818 4759 37846 4787
rect 15818 4747 15824 4759
rect 37840 4747 37846 4759
rect 37898 4747 37904 4799
rect 1152 4688 58848 4710
rect 1152 4636 19654 4688
rect 19706 4636 19718 4688
rect 19770 4636 19782 4688
rect 19834 4636 19846 4688
rect 19898 4636 50374 4688
rect 50426 4636 50438 4688
rect 50490 4636 50502 4688
rect 50554 4636 50566 4688
rect 50618 4636 58848 4688
rect 1152 4614 58848 4636
rect 15760 4565 15766 4577
rect 15721 4537 15766 4565
rect 15760 4525 15766 4537
rect 15818 4525 15824 4577
rect 19120 4565 19126 4577
rect 19081 4537 19126 4565
rect 19120 4525 19126 4537
rect 19178 4525 19184 4577
rect 23920 4525 23926 4577
rect 23978 4565 23984 4577
rect 24400 4565 24406 4577
rect 23978 4537 24406 4565
rect 23978 4525 23984 4537
rect 24400 4525 24406 4537
rect 24458 4525 24464 4577
rect 34192 4525 34198 4577
rect 34250 4565 34256 4577
rect 38131 4568 38189 4574
rect 38131 4565 38143 4568
rect 34250 4537 38143 4565
rect 34250 4525 34256 4537
rect 38131 4534 38143 4537
rect 38177 4565 38189 4568
rect 38323 4568 38381 4574
rect 38323 4565 38335 4568
rect 38177 4537 38335 4565
rect 38177 4534 38189 4537
rect 38131 4528 38189 4534
rect 38323 4534 38335 4537
rect 38369 4534 38381 4568
rect 38323 4528 38381 4534
rect 4720 4491 4726 4503
rect 4642 4463 4726 4491
rect 784 4377 790 4429
rect 842 4417 848 4429
rect 842 4389 2366 4417
rect 842 4377 848 4389
rect 1168 4303 1174 4355
rect 1226 4343 1232 4355
rect 2338 4352 2366 4389
rect 1555 4346 1613 4352
rect 1555 4343 1567 4346
rect 1226 4315 1567 4343
rect 1226 4303 1232 4315
rect 1555 4312 1567 4315
rect 1601 4312 1613 4346
rect 1555 4306 1613 4312
rect 2323 4346 2381 4352
rect 2323 4312 2335 4346
rect 2369 4312 2381 4346
rect 2323 4306 2381 4312
rect 3091 4346 3149 4352
rect 3091 4312 3103 4346
rect 3137 4312 3149 4346
rect 3091 4306 3149 4312
rect 4339 4346 4397 4352
rect 4339 4312 4351 4346
rect 4385 4312 4397 4346
rect 4339 4306 4397 4312
rect 1360 4229 1366 4281
rect 1418 4269 1424 4281
rect 3106 4269 3134 4306
rect 1418 4241 3134 4269
rect 1418 4229 1424 4241
rect 3760 4229 3766 4281
rect 3818 4269 3824 4281
rect 4354 4269 4382 4306
rect 3818 4241 4382 4269
rect 3818 4229 3824 4241
rect 4642 4195 4670 4463
rect 4720 4451 4726 4463
rect 4778 4451 4784 4503
rect 16531 4494 16589 4500
rect 16531 4460 16543 4494
rect 16577 4460 16589 4494
rect 16531 4454 16589 4460
rect 17299 4494 17357 4500
rect 17299 4460 17311 4494
rect 17345 4491 17357 4494
rect 42928 4491 42934 4503
rect 17345 4463 42934 4491
rect 17345 4460 17357 4463
rect 17299 4454 17357 4460
rect 16546 4417 16574 4454
rect 42928 4451 42934 4463
rect 42986 4451 42992 4503
rect 43024 4417 43030 4429
rect 16546 4389 43030 4417
rect 43024 4377 43030 4389
rect 43082 4377 43088 4429
rect 4720 4303 4726 4355
rect 4778 4343 4784 4355
rect 5107 4346 5165 4352
rect 5107 4343 5119 4346
rect 4778 4315 5119 4343
rect 4778 4303 4784 4315
rect 5107 4312 5119 4315
rect 5153 4312 5165 4346
rect 5875 4346 5933 4352
rect 5875 4343 5887 4346
rect 5107 4306 5165 4312
rect 5602 4315 5887 4343
rect 5008 4229 5014 4281
rect 5066 4269 5072 4281
rect 5602 4269 5630 4315
rect 5875 4312 5887 4315
rect 5921 4312 5933 4346
rect 5875 4306 5933 4312
rect 6643 4346 6701 4352
rect 6643 4312 6655 4346
rect 6689 4312 6701 4346
rect 7408 4343 7414 4355
rect 7369 4315 7414 4343
rect 6643 4306 6701 4312
rect 5066 4241 5630 4269
rect 5066 4229 5072 4241
rect 5680 4229 5686 4281
rect 5738 4269 5744 4281
rect 6658 4269 6686 4306
rect 7408 4303 7414 4315
rect 7466 4303 7472 4355
rect 8179 4346 8237 4352
rect 8179 4312 8191 4346
rect 8225 4312 8237 4346
rect 9616 4343 9622 4355
rect 9577 4315 9622 4343
rect 8179 4306 8237 4312
rect 5738 4241 6686 4269
rect 5738 4229 5744 4241
rect 6160 4195 6166 4207
rect 4642 4167 6166 4195
rect 6160 4155 6166 4167
rect 6218 4155 6224 4207
rect 6448 4155 6454 4207
rect 6506 4195 6512 4207
rect 8194 4195 8222 4306
rect 9616 4303 9622 4315
rect 9674 4303 9680 4355
rect 10384 4343 10390 4355
rect 10345 4315 10390 4343
rect 10384 4303 10390 4315
rect 10442 4303 10448 4355
rect 10768 4303 10774 4355
rect 10826 4343 10832 4355
rect 11155 4346 11213 4352
rect 11155 4343 11167 4346
rect 10826 4315 11167 4343
rect 10826 4303 10832 4315
rect 11155 4312 11167 4315
rect 11201 4312 11213 4346
rect 11155 4306 11213 4312
rect 11923 4346 11981 4352
rect 11923 4312 11935 4346
rect 11969 4312 11981 4346
rect 11923 4306 11981 4312
rect 12691 4346 12749 4352
rect 12691 4312 12703 4346
rect 12737 4312 12749 4346
rect 13552 4343 13558 4355
rect 13513 4315 13558 4343
rect 12691 4306 12749 4312
rect 6506 4167 8222 4195
rect 6506 4155 6512 4167
rect 11152 4155 11158 4207
rect 11210 4195 11216 4207
rect 11938 4195 11966 4306
rect 11210 4167 11966 4195
rect 11210 4155 11216 4167
rect 11440 4081 11446 4133
rect 11498 4121 11504 4133
rect 12706 4121 12734 4306
rect 13552 4303 13558 4315
rect 13610 4303 13616 4355
rect 15472 4343 15478 4355
rect 15433 4315 15478 4343
rect 15472 4303 15478 4315
rect 15530 4303 15536 4355
rect 15952 4303 15958 4355
rect 16010 4343 16016 4355
rect 16243 4346 16301 4352
rect 16243 4343 16255 4346
rect 16010 4315 16255 4343
rect 16010 4303 16016 4315
rect 16243 4312 16255 4315
rect 16289 4312 16301 4346
rect 16243 4306 16301 4312
rect 17011 4346 17069 4352
rect 17011 4312 17023 4346
rect 17057 4312 17069 4346
rect 17011 4306 17069 4312
rect 17779 4346 17837 4352
rect 17779 4312 17791 4346
rect 17825 4312 17837 4346
rect 18832 4343 18838 4355
rect 18793 4315 18838 4343
rect 17779 4306 17837 4312
rect 16240 4155 16246 4207
rect 16298 4195 16304 4207
rect 17026 4195 17054 4306
rect 17794 4269 17822 4306
rect 18832 4303 18838 4315
rect 18890 4303 18896 4355
rect 20179 4346 20237 4352
rect 20179 4312 20191 4346
rect 20225 4312 20237 4346
rect 21040 4343 21046 4355
rect 21001 4315 21046 4343
rect 20179 4306 20237 4312
rect 16298 4167 17054 4195
rect 17122 4241 17822 4269
rect 16298 4155 16304 4167
rect 11498 4093 12734 4121
rect 11498 4081 11504 4093
rect 16912 4081 16918 4133
rect 16970 4121 16976 4133
rect 17122 4121 17150 4241
rect 19504 4229 19510 4281
rect 19562 4269 19568 4281
rect 20194 4269 20222 4306
rect 21040 4303 21046 4315
rect 21098 4303 21104 4355
rect 21808 4343 21814 4355
rect 21769 4315 21814 4343
rect 21808 4303 21814 4315
rect 21866 4303 21872 4355
rect 23248 4343 23254 4355
rect 23209 4315 23254 4343
rect 23248 4303 23254 4315
rect 23306 4303 23312 4355
rect 24016 4343 24022 4355
rect 23977 4315 24022 4343
rect 24016 4303 24022 4315
rect 24074 4303 24080 4355
rect 25456 4343 25462 4355
rect 25417 4315 25462 4343
rect 25456 4303 25462 4315
rect 25514 4303 25520 4355
rect 26128 4303 26134 4355
rect 26186 4343 26192 4355
rect 26227 4346 26285 4352
rect 26227 4343 26239 4346
rect 26186 4315 26239 4343
rect 26186 4303 26192 4315
rect 26227 4312 26239 4315
rect 26273 4312 26285 4346
rect 26227 4306 26285 4312
rect 26512 4303 26518 4355
rect 26570 4343 26576 4355
rect 26995 4346 27053 4352
rect 26995 4343 27007 4346
rect 26570 4315 27007 4343
rect 26570 4303 26576 4315
rect 26995 4312 27007 4315
rect 27041 4312 27053 4346
rect 28336 4343 28342 4355
rect 28297 4315 28342 4343
rect 26995 4306 27053 4312
rect 28336 4303 28342 4315
rect 28394 4303 28400 4355
rect 29104 4343 29110 4355
rect 29065 4315 29110 4343
rect 29104 4303 29110 4315
rect 29162 4303 29168 4355
rect 30928 4343 30934 4355
rect 30889 4315 30934 4343
rect 30928 4303 30934 4315
rect 30986 4303 30992 4355
rect 31696 4343 31702 4355
rect 31657 4315 31702 4343
rect 31696 4303 31702 4315
rect 31754 4303 31760 4355
rect 32752 4343 32758 4355
rect 32713 4315 32758 4343
rect 32752 4303 32758 4315
rect 32810 4303 32816 4355
rect 33904 4343 33910 4355
rect 33865 4315 33910 4343
rect 33904 4303 33910 4315
rect 33962 4303 33968 4355
rect 34576 4303 34582 4355
rect 34634 4343 34640 4355
rect 34675 4346 34733 4352
rect 34675 4343 34687 4346
rect 34634 4315 34687 4343
rect 34634 4303 34640 4315
rect 34675 4312 34687 4315
rect 34721 4312 34733 4346
rect 36019 4346 36077 4352
rect 36019 4343 36031 4346
rect 34675 4306 34733 4312
rect 34786 4315 36031 4343
rect 19562 4241 20222 4269
rect 19562 4229 19568 4241
rect 20944 4229 20950 4281
rect 21002 4269 21008 4281
rect 21712 4269 21718 4281
rect 21002 4241 21718 4269
rect 21002 4229 21008 4241
rect 21712 4229 21718 4241
rect 21770 4229 21776 4281
rect 22771 4272 22829 4278
rect 22771 4238 22783 4272
rect 22817 4269 22829 4272
rect 28048 4269 28054 4281
rect 22817 4241 28054 4269
rect 22817 4238 22829 4241
rect 22771 4232 22829 4238
rect 28048 4229 28054 4241
rect 28106 4229 28112 4281
rect 28528 4229 28534 4281
rect 28586 4269 28592 4281
rect 29392 4269 29398 4281
rect 28586 4241 29398 4269
rect 28586 4229 28592 4241
rect 29392 4229 29398 4241
rect 29450 4229 29456 4281
rect 33106 4241 33854 4269
rect 20080 4155 20086 4207
rect 20138 4195 20144 4207
rect 21424 4195 21430 4207
rect 20138 4167 21430 4195
rect 20138 4155 20144 4167
rect 21424 4155 21430 4167
rect 21482 4155 21488 4207
rect 21520 4155 21526 4207
rect 21578 4195 21584 4207
rect 22864 4195 22870 4207
rect 21578 4167 22870 4195
rect 21578 4155 21584 4167
rect 22864 4155 22870 4167
rect 22922 4155 22928 4207
rect 24112 4155 24118 4207
rect 24170 4195 24176 4207
rect 24496 4195 24502 4207
rect 24170 4167 24502 4195
rect 24170 4155 24176 4167
rect 24496 4155 24502 4167
rect 24554 4155 24560 4207
rect 25552 4155 25558 4207
rect 25610 4195 25616 4207
rect 25936 4195 25942 4207
rect 25610 4167 25942 4195
rect 25610 4155 25616 4167
rect 25936 4155 25942 4167
rect 25994 4155 26000 4207
rect 26992 4155 26998 4207
rect 27050 4195 27056 4207
rect 27376 4195 27382 4207
rect 27050 4167 27382 4195
rect 27050 4155 27056 4167
rect 27376 4155 27382 4167
rect 27434 4155 27440 4207
rect 28240 4155 28246 4207
rect 28298 4195 28304 4207
rect 29008 4195 29014 4207
rect 28298 4167 29014 4195
rect 28298 4155 28304 4167
rect 29008 4155 29014 4167
rect 29066 4155 29072 4207
rect 16970 4093 17150 4121
rect 16970 4081 16976 4093
rect 18256 4081 18262 4133
rect 18314 4121 18320 4133
rect 33106 4121 33134 4241
rect 33826 4195 33854 4241
rect 34192 4229 34198 4281
rect 34250 4269 34256 4281
rect 34786 4269 34814 4315
rect 36019 4312 36031 4315
rect 36065 4312 36077 4346
rect 36784 4343 36790 4355
rect 36745 4315 36790 4343
rect 36019 4306 36077 4312
rect 36784 4303 36790 4315
rect 36842 4303 36848 4355
rect 37555 4346 37613 4352
rect 37555 4312 37567 4346
rect 37601 4312 37613 4346
rect 38992 4343 38998 4355
rect 38953 4315 38998 4343
rect 37555 4306 37613 4312
rect 34250 4241 34814 4269
rect 34250 4229 34256 4241
rect 37168 4229 37174 4281
rect 37226 4269 37232 4281
rect 37570 4269 37598 4306
rect 38992 4303 38998 4315
rect 39050 4303 39056 4355
rect 39760 4343 39766 4355
rect 39721 4315 39766 4343
rect 39760 4303 39766 4315
rect 39818 4303 39824 4355
rect 41968 4343 41974 4355
rect 41929 4315 41974 4343
rect 41968 4303 41974 4315
rect 42026 4303 42032 4355
rect 42256 4303 42262 4355
rect 42314 4343 42320 4355
rect 42739 4346 42797 4352
rect 42739 4343 42751 4346
rect 42314 4315 42751 4343
rect 42314 4303 42320 4315
rect 42739 4312 42751 4315
rect 42785 4312 42797 4346
rect 42739 4306 42797 4312
rect 43408 4303 43414 4355
rect 43466 4343 43472 4355
rect 43507 4346 43565 4352
rect 43507 4343 43519 4346
rect 43466 4315 43519 4343
rect 43466 4303 43472 4315
rect 43507 4312 43519 4315
rect 43553 4312 43565 4346
rect 44944 4343 44950 4355
rect 44905 4315 44950 4343
rect 43507 4306 43565 4312
rect 44944 4303 44950 4315
rect 45002 4303 45008 4355
rect 46768 4343 46774 4355
rect 46729 4315 46774 4343
rect 46768 4303 46774 4315
rect 46826 4303 46832 4355
rect 47539 4346 47597 4352
rect 47539 4312 47551 4346
rect 47585 4312 47597 4346
rect 47539 4306 47597 4312
rect 37226 4241 37598 4269
rect 37226 4229 37232 4241
rect 41392 4229 41398 4281
rect 41450 4269 41456 4281
rect 41584 4269 41590 4281
rect 41450 4241 41590 4269
rect 41450 4229 41456 4241
rect 41584 4229 41590 4241
rect 41642 4229 41648 4281
rect 42064 4229 42070 4281
rect 42122 4269 42128 4281
rect 43120 4269 43126 4281
rect 42122 4241 43126 4269
rect 42122 4229 42128 4241
rect 43120 4229 43126 4241
rect 43178 4229 43184 4281
rect 44080 4229 44086 4281
rect 44138 4269 44144 4281
rect 44656 4269 44662 4281
rect 44138 4241 44662 4269
rect 44138 4229 44144 4241
rect 44656 4229 44662 4241
rect 44714 4229 44720 4281
rect 47440 4229 47446 4281
rect 47498 4269 47504 4281
rect 47554 4269 47582 4306
rect 47824 4303 47830 4355
rect 47882 4343 47888 4355
rect 48307 4346 48365 4352
rect 48307 4343 48319 4346
rect 47882 4315 48319 4343
rect 47882 4303 47888 4315
rect 48307 4312 48319 4315
rect 48353 4312 48365 4346
rect 48307 4306 48365 4312
rect 49075 4346 49133 4352
rect 49075 4312 49087 4346
rect 49121 4312 49133 4346
rect 49075 4306 49133 4312
rect 47498 4241 47582 4269
rect 47498 4229 47504 4241
rect 48592 4229 48598 4281
rect 48650 4269 48656 4281
rect 49090 4269 49118 4306
rect 49168 4303 49174 4355
rect 49226 4343 49232 4355
rect 49843 4346 49901 4352
rect 49843 4343 49855 4346
rect 49226 4315 49855 4343
rect 49226 4303 49232 4315
rect 49843 4312 49855 4315
rect 49889 4312 49901 4346
rect 49843 4306 49901 4312
rect 50611 4346 50669 4352
rect 50611 4312 50623 4346
rect 50657 4312 50669 4346
rect 50611 4306 50669 4312
rect 51859 4346 51917 4352
rect 51859 4312 51871 4346
rect 51905 4312 51917 4346
rect 52624 4343 52630 4355
rect 52585 4315 52630 4343
rect 51859 4306 51917 4312
rect 48650 4241 49118 4269
rect 48650 4229 48656 4241
rect 41491 4198 41549 4204
rect 41491 4195 41503 4198
rect 33826 4167 41503 4195
rect 41491 4164 41503 4167
rect 41537 4164 41549 4198
rect 41491 4158 41549 4164
rect 48112 4155 48118 4207
rect 48170 4195 48176 4207
rect 48976 4195 48982 4207
rect 48170 4167 48982 4195
rect 48170 4155 48176 4167
rect 48976 4155 48982 4167
rect 49034 4155 49040 4207
rect 49840 4155 49846 4207
rect 49898 4195 49904 4207
rect 50626 4195 50654 4306
rect 50992 4229 50998 4281
rect 51050 4269 51056 4281
rect 51874 4269 51902 4306
rect 52624 4303 52630 4315
rect 52682 4303 52688 4355
rect 53395 4346 53453 4352
rect 53395 4312 53407 4346
rect 53441 4312 53453 4346
rect 53395 4306 53453 4312
rect 51050 4241 51902 4269
rect 51050 4229 51056 4241
rect 53008 4229 53014 4281
rect 53066 4269 53072 4281
rect 53410 4269 53438 4306
rect 54064 4303 54070 4355
rect 54122 4343 54128 4355
rect 54163 4346 54221 4352
rect 54163 4343 54175 4346
rect 54122 4315 54175 4343
rect 54122 4303 54128 4315
rect 54163 4312 54175 4315
rect 54209 4312 54221 4346
rect 55600 4343 55606 4355
rect 55561 4315 55606 4343
rect 54163 4306 54221 4312
rect 55600 4303 55606 4315
rect 55658 4303 55664 4355
rect 56656 4303 56662 4355
rect 56714 4343 56720 4355
rect 57139 4346 57197 4352
rect 57139 4343 57151 4346
rect 56714 4315 57151 4343
rect 56714 4303 56720 4315
rect 57139 4312 57151 4315
rect 57185 4312 57197 4346
rect 57139 4306 57197 4312
rect 53066 4241 53438 4269
rect 53066 4229 53072 4241
rect 54832 4229 54838 4281
rect 54890 4269 54896 4281
rect 55123 4272 55181 4278
rect 55123 4269 55135 4272
rect 54890 4241 55135 4269
rect 54890 4229 54896 4241
rect 55123 4238 55135 4241
rect 55169 4238 55181 4272
rect 58288 4269 58294 4281
rect 55123 4232 55181 4238
rect 57586 4241 58294 4269
rect 49898 4167 50654 4195
rect 49898 4155 49904 4167
rect 57136 4155 57142 4207
rect 57194 4195 57200 4207
rect 57586 4195 57614 4241
rect 58288 4229 58294 4241
rect 58346 4229 58352 4281
rect 57194 4167 57614 4195
rect 57194 4155 57200 4167
rect 18314 4093 33134 4121
rect 18314 4081 18320 4093
rect 33808 4081 33814 4133
rect 33866 4121 33872 4133
rect 34672 4121 34678 4133
rect 33866 4093 34678 4121
rect 33866 4081 33872 4093
rect 34672 4081 34678 4093
rect 34730 4081 34736 4133
rect 36688 4081 36694 4133
rect 36746 4121 36752 4133
rect 37552 4121 37558 4133
rect 36746 4093 37558 4121
rect 36746 4081 36752 4093
rect 37552 4081 37558 4093
rect 37610 4081 37616 4133
rect 38512 4081 38518 4133
rect 38570 4121 38576 4133
rect 40144 4121 40150 4133
rect 38570 4093 40150 4121
rect 38570 4081 38576 4093
rect 40144 4081 40150 4093
rect 40202 4081 40208 4133
rect 43792 4081 43798 4133
rect 43850 4121 43856 4133
rect 47152 4121 47158 4133
rect 43850 4093 47158 4121
rect 43850 4081 43856 4093
rect 47152 4081 47158 4093
rect 47210 4081 47216 4133
rect 48496 4081 48502 4133
rect 48554 4121 48560 4133
rect 49648 4121 49654 4133
rect 48554 4093 49654 4121
rect 48554 4081 48560 4093
rect 49648 4081 49654 4093
rect 49706 4081 49712 4133
rect 56560 4081 56566 4133
rect 56618 4121 56624 4133
rect 59152 4121 59158 4133
rect 56618 4093 59158 4121
rect 56618 4081 56624 4093
rect 59152 4081 59158 4093
rect 59210 4081 59216 4133
rect 1152 4022 58848 4044
rect 1152 3970 4294 4022
rect 4346 3970 4358 4022
rect 4410 3970 4422 4022
rect 4474 3970 4486 4022
rect 4538 3970 35014 4022
rect 35066 3970 35078 4022
rect 35130 3970 35142 4022
rect 35194 3970 35206 4022
rect 35258 3970 58848 4022
rect 1152 3948 58848 3970
rect 1936 3859 1942 3911
rect 1994 3899 2000 3911
rect 3376 3899 3382 3911
rect 1994 3871 3382 3899
rect 1994 3859 2000 3871
rect 3376 3859 3382 3871
rect 3434 3859 3440 3911
rect 8752 3859 8758 3911
rect 8810 3899 8816 3911
rect 10288 3899 10294 3911
rect 8810 3871 10294 3899
rect 8810 3859 8816 3871
rect 10288 3859 10294 3871
rect 10346 3859 10352 3911
rect 15376 3859 15382 3911
rect 15434 3899 15440 3911
rect 16432 3899 16438 3911
rect 15434 3871 16438 3899
rect 15434 3859 15440 3871
rect 16432 3859 16438 3871
rect 16490 3859 16496 3911
rect 18352 3859 18358 3911
rect 18410 3899 18416 3911
rect 19024 3899 19030 3911
rect 18410 3871 19030 3899
rect 18410 3859 18416 3871
rect 19024 3859 19030 3871
rect 19082 3859 19088 3911
rect 21328 3859 21334 3911
rect 21386 3899 21392 3911
rect 22768 3899 22774 3911
rect 21386 3871 22774 3899
rect 21386 3859 21392 3871
rect 22768 3859 22774 3871
rect 22826 3859 22832 3911
rect 24496 3859 24502 3911
rect 24554 3899 24560 3911
rect 24880 3899 24886 3911
rect 24554 3871 24886 3899
rect 24554 3859 24560 3871
rect 24880 3859 24886 3871
rect 24938 3859 24944 3911
rect 25360 3859 25366 3911
rect 25418 3899 25424 3911
rect 26224 3899 26230 3911
rect 25418 3871 26230 3899
rect 25418 3859 25424 3871
rect 26224 3859 26230 3871
rect 26282 3859 26288 3911
rect 27472 3859 27478 3911
rect 27530 3899 27536 3911
rect 28912 3899 28918 3911
rect 27530 3871 28918 3899
rect 27530 3859 27536 3871
rect 28912 3859 28918 3871
rect 28970 3859 28976 3911
rect 29008 3859 29014 3911
rect 29066 3899 29072 3911
rect 30352 3899 30358 3911
rect 29066 3871 30358 3899
rect 29066 3859 29072 3871
rect 30352 3859 30358 3871
rect 30410 3859 30416 3911
rect 34480 3859 34486 3911
rect 34538 3899 34544 3911
rect 35632 3899 35638 3911
rect 34538 3871 35638 3899
rect 34538 3859 34544 3871
rect 35632 3859 35638 3871
rect 35690 3859 35696 3911
rect 38128 3859 38134 3911
rect 38186 3899 38192 3911
rect 39088 3899 39094 3911
rect 38186 3871 39094 3899
rect 38186 3859 38192 3871
rect 39088 3859 39094 3871
rect 39146 3859 39152 3911
rect 39664 3859 39670 3911
rect 39722 3899 39728 3911
rect 40912 3899 40918 3911
rect 39722 3871 40918 3899
rect 39722 3859 39728 3871
rect 40912 3859 40918 3871
rect 40970 3859 40976 3911
rect 41200 3859 41206 3911
rect 41258 3899 41264 3911
rect 41258 3871 43646 3899
rect 41258 3859 41264 3871
rect 496 3785 502 3837
rect 554 3825 560 3837
rect 1648 3825 1654 3837
rect 554 3797 1654 3825
rect 554 3785 560 3797
rect 1648 3785 1654 3797
rect 1706 3785 1712 3837
rect 2320 3785 2326 3837
rect 2378 3825 2384 3837
rect 3088 3825 3094 3837
rect 2378 3797 3094 3825
rect 2378 3785 2384 3797
rect 3088 3785 3094 3797
rect 3146 3785 3152 3837
rect 8272 3785 8278 3837
rect 8330 3825 8336 3837
rect 9232 3825 9238 3837
rect 8330 3797 9238 3825
rect 8330 3785 8336 3797
rect 9232 3785 9238 3797
rect 9290 3785 9296 3837
rect 12016 3785 12022 3837
rect 12074 3825 12080 3837
rect 13360 3825 13366 3837
rect 12074 3797 13366 3825
rect 12074 3785 12080 3797
rect 13360 3785 13366 3797
rect 13418 3785 13424 3837
rect 13648 3785 13654 3837
rect 13706 3825 13712 3837
rect 18256 3825 18262 3837
rect 13706 3797 18262 3825
rect 13706 3785 13712 3797
rect 18256 3785 18262 3797
rect 18314 3785 18320 3837
rect 20179 3828 20237 3834
rect 20179 3794 20191 3828
rect 20225 3825 20237 3828
rect 22384 3825 22390 3837
rect 20225 3797 22390 3825
rect 20225 3794 20237 3797
rect 20179 3788 20237 3794
rect 22384 3785 22390 3797
rect 22442 3785 22448 3837
rect 24208 3785 24214 3837
rect 24266 3825 24272 3837
rect 25840 3825 25846 3837
rect 24266 3797 25846 3825
rect 24266 3785 24272 3797
rect 25840 3785 25846 3797
rect 25898 3785 25904 3837
rect 25936 3785 25942 3837
rect 25994 3825 26000 3837
rect 27088 3825 27094 3837
rect 25994 3797 27094 3825
rect 25994 3785 26000 3797
rect 27088 3785 27094 3797
rect 27146 3785 27152 3837
rect 28048 3785 28054 3837
rect 28106 3825 28112 3837
rect 35440 3825 35446 3837
rect 28106 3797 35446 3825
rect 28106 3785 28112 3797
rect 35440 3785 35446 3797
rect 35498 3785 35504 3837
rect 36016 3785 36022 3837
rect 36074 3825 36080 3837
rect 36400 3825 36406 3837
rect 36074 3797 36406 3825
rect 36074 3785 36080 3797
rect 36400 3785 36406 3797
rect 36458 3785 36464 3837
rect 37072 3785 37078 3837
rect 37130 3825 37136 3837
rect 38608 3825 38614 3837
rect 37130 3797 38614 3825
rect 37130 3785 37136 3797
rect 38608 3785 38614 3797
rect 38666 3785 38672 3837
rect 42544 3785 42550 3837
rect 42602 3825 42608 3837
rect 43504 3825 43510 3837
rect 42602 3797 43510 3825
rect 42602 3785 42608 3797
rect 43504 3785 43510 3797
rect 43562 3785 43568 3837
rect 43618 3825 43646 3871
rect 43696 3859 43702 3911
rect 43754 3899 43760 3911
rect 44848 3899 44854 3911
rect 43754 3871 44854 3899
rect 43754 3859 43760 3871
rect 44848 3859 44854 3871
rect 44906 3859 44912 3911
rect 46288 3859 46294 3911
rect 46346 3899 46352 3911
rect 47920 3899 47926 3911
rect 46346 3871 47926 3899
rect 46346 3859 46352 3871
rect 47920 3859 47926 3871
rect 47978 3859 47984 3911
rect 49264 3859 49270 3911
rect 49322 3899 49328 3911
rect 50704 3899 50710 3911
rect 49322 3871 50710 3899
rect 49322 3859 49328 3871
rect 50704 3859 50710 3871
rect 50762 3859 50768 3911
rect 51376 3859 51382 3911
rect 51434 3899 51440 3911
rect 51856 3899 51862 3911
rect 51434 3871 51862 3899
rect 51434 3859 51440 3871
rect 51856 3859 51862 3871
rect 51914 3859 51920 3911
rect 55984 3859 55990 3911
rect 56042 3899 56048 3911
rect 56042 3871 57614 3899
rect 56042 3859 56048 3871
rect 43792 3825 43798 3837
rect 43618 3797 43798 3825
rect 43792 3785 43798 3797
rect 43850 3785 43856 3837
rect 44464 3785 44470 3837
rect 44522 3825 44528 3837
rect 45616 3825 45622 3837
rect 44522 3797 45622 3825
rect 44522 3785 44528 3797
rect 45616 3785 45622 3797
rect 45674 3785 45680 3837
rect 56752 3785 56758 3837
rect 56810 3825 56816 3837
rect 57136 3825 57142 3837
rect 56810 3797 57142 3825
rect 56810 3785 56816 3797
rect 57136 3785 57142 3797
rect 57194 3785 57200 3837
rect 57586 3825 57614 3871
rect 57904 3825 57910 3837
rect 57586 3797 57910 3825
rect 57904 3785 57910 3797
rect 57962 3785 57968 3837
rect 976 3711 982 3763
rect 1034 3751 1040 3763
rect 2416 3751 2422 3763
rect 1034 3723 2422 3751
rect 1034 3711 1040 3723
rect 2416 3711 2422 3723
rect 2474 3711 2480 3763
rect 3376 3711 3382 3763
rect 3434 3751 3440 3763
rect 3434 3723 4670 3751
rect 3434 3711 3440 3723
rect 112 3637 118 3689
rect 170 3677 176 3689
rect 1555 3680 1613 3686
rect 1555 3677 1567 3680
rect 170 3649 1567 3677
rect 170 3637 176 3649
rect 1555 3646 1567 3649
rect 1601 3646 1613 3680
rect 1555 3640 1613 3646
rect 1648 3637 1654 3689
rect 1706 3677 1712 3689
rect 2323 3680 2381 3686
rect 2323 3677 2335 3680
rect 1706 3649 2335 3677
rect 1706 3637 1712 3649
rect 2323 3646 2335 3649
rect 2369 3646 2381 3680
rect 2323 3640 2381 3646
rect 2704 3637 2710 3689
rect 2762 3677 2768 3689
rect 4642 3686 4670 3723
rect 10288 3711 10294 3763
rect 10346 3751 10352 3763
rect 11056 3751 11062 3763
rect 10346 3723 11062 3751
rect 10346 3711 10352 3723
rect 11056 3711 11062 3723
rect 11114 3711 11120 3763
rect 13555 3754 13613 3760
rect 13555 3720 13567 3754
rect 13601 3751 13613 3754
rect 14224 3751 14230 3763
rect 13601 3723 14230 3751
rect 13601 3720 13613 3723
rect 13555 3714 13613 3720
rect 14224 3711 14230 3723
rect 14282 3711 14288 3763
rect 14416 3711 14422 3763
rect 14474 3751 14480 3763
rect 15283 3754 15341 3760
rect 15283 3751 15295 3754
rect 14474 3723 15295 3751
rect 14474 3711 14480 3723
rect 15283 3720 15295 3723
rect 15329 3720 15341 3754
rect 15283 3714 15341 3720
rect 17683 3754 17741 3760
rect 17683 3720 17695 3754
rect 17729 3751 17741 3754
rect 17776 3751 17782 3763
rect 17729 3723 17782 3751
rect 17729 3720 17741 3723
rect 17683 3714 17741 3720
rect 17776 3711 17782 3723
rect 17834 3711 17840 3763
rect 18544 3751 18550 3763
rect 18505 3723 18550 3751
rect 18544 3711 18550 3723
rect 18602 3711 18608 3763
rect 19408 3711 19414 3763
rect 19466 3751 19472 3763
rect 20560 3751 20566 3763
rect 19466 3723 20566 3751
rect 19466 3711 19472 3723
rect 20560 3711 20566 3723
rect 20618 3711 20624 3763
rect 22096 3711 22102 3763
rect 22154 3751 22160 3763
rect 24016 3751 24022 3763
rect 22154 3723 24022 3751
rect 22154 3711 22160 3723
rect 24016 3711 24022 3723
rect 24074 3711 24080 3763
rect 26320 3711 26326 3763
rect 26378 3751 26384 3763
rect 27568 3751 27574 3763
rect 26378 3723 27574 3751
rect 26378 3711 26384 3723
rect 27568 3711 27574 3723
rect 27626 3711 27632 3763
rect 28720 3711 28726 3763
rect 28778 3751 28784 3763
rect 28778 3723 29630 3751
rect 28778 3711 28784 3723
rect 3091 3680 3149 3686
rect 3091 3677 3103 3680
rect 2762 3649 3103 3677
rect 2762 3637 2768 3649
rect 3091 3646 3103 3649
rect 3137 3646 3149 3680
rect 3091 3640 3149 3646
rect 3859 3680 3917 3686
rect 3859 3646 3871 3680
rect 3905 3646 3917 3680
rect 3859 3640 3917 3646
rect 4627 3680 4685 3686
rect 4627 3646 4639 3680
rect 4673 3646 4685 3680
rect 5584 3677 5590 3689
rect 5545 3649 5590 3677
rect 4627 3640 4685 3646
rect 208 3563 214 3615
rect 266 3603 272 3615
rect 1744 3603 1750 3615
rect 266 3575 1750 3603
rect 266 3563 272 3575
rect 1744 3563 1750 3575
rect 1802 3563 1808 3615
rect 3088 3489 3094 3541
rect 3146 3529 3152 3541
rect 3874 3529 3902 3640
rect 5584 3637 5590 3649
rect 5642 3637 5648 3689
rect 6352 3637 6358 3689
rect 6410 3677 6416 3689
rect 6931 3680 6989 3686
rect 6931 3677 6943 3680
rect 6410 3649 6943 3677
rect 6410 3637 6416 3649
rect 6931 3646 6943 3649
rect 6977 3646 6989 3680
rect 6931 3640 6989 3646
rect 7024 3637 7030 3689
rect 7082 3677 7088 3689
rect 7699 3680 7757 3686
rect 7699 3677 7711 3680
rect 7082 3649 7711 3677
rect 7082 3637 7088 3649
rect 7699 3646 7711 3649
rect 7745 3646 7757 3680
rect 7699 3640 7757 3646
rect 7792 3637 7798 3689
rect 7850 3677 7856 3689
rect 8467 3680 8525 3686
rect 8467 3677 8479 3680
rect 7850 3649 8479 3677
rect 7850 3637 7856 3649
rect 8467 3646 8479 3649
rect 8513 3646 8525 3680
rect 8467 3640 8525 3646
rect 8560 3637 8566 3689
rect 8618 3677 8624 3689
rect 9235 3680 9293 3686
rect 9235 3677 9247 3680
rect 8618 3649 9247 3677
rect 8618 3637 8624 3649
rect 9235 3646 9247 3649
rect 9281 3646 9293 3680
rect 9235 3640 9293 3646
rect 9328 3637 9334 3689
rect 9386 3677 9392 3689
rect 10003 3680 10061 3686
rect 10003 3677 10015 3680
rect 9386 3649 10015 3677
rect 9386 3637 9392 3649
rect 10003 3646 10015 3649
rect 10049 3646 10061 3680
rect 10003 3640 10061 3646
rect 10771 3680 10829 3686
rect 10771 3646 10783 3680
rect 10817 3646 10829 3680
rect 10771 3640 10829 3646
rect 12691 3680 12749 3686
rect 12691 3646 12703 3680
rect 12737 3677 12749 3680
rect 13168 3677 13174 3689
rect 12737 3649 13174 3677
rect 12737 3646 12749 3649
rect 12691 3640 12749 3646
rect 3146 3501 3902 3529
rect 3146 3489 3152 3501
rect 10000 3489 10006 3541
rect 10058 3529 10064 3541
rect 10786 3529 10814 3640
rect 13168 3637 13174 3649
rect 13226 3637 13232 3689
rect 13360 3637 13366 3689
rect 13418 3677 13424 3689
rect 13747 3680 13805 3686
rect 13747 3677 13759 3680
rect 13418 3649 13759 3677
rect 13418 3637 13424 3649
rect 13747 3646 13759 3649
rect 13793 3646 13805 3680
rect 14611 3680 14669 3686
rect 14611 3677 14623 3680
rect 13747 3640 13805 3646
rect 13858 3649 14623 3677
rect 13648 3563 13654 3615
rect 13706 3603 13712 3615
rect 13858 3603 13886 3649
rect 14611 3646 14623 3649
rect 14657 3646 14669 3680
rect 14611 3640 14669 3646
rect 15184 3637 15190 3689
rect 15242 3677 15248 3689
rect 15859 3680 15917 3686
rect 15859 3677 15871 3680
rect 15242 3649 15871 3677
rect 15242 3637 15248 3649
rect 15859 3646 15871 3649
rect 15905 3646 15917 3680
rect 15859 3640 15917 3646
rect 17392 3637 17398 3689
rect 17450 3677 17456 3689
rect 17875 3680 17933 3686
rect 17875 3677 17887 3680
rect 17450 3649 17887 3677
rect 17450 3637 17456 3649
rect 17875 3646 17887 3649
rect 17921 3646 17933 3680
rect 17875 3640 17933 3646
rect 18256 3637 18262 3689
rect 18314 3677 18320 3689
rect 18739 3680 18797 3686
rect 18739 3677 18751 3680
rect 18314 3649 18751 3677
rect 18314 3637 18320 3649
rect 18739 3646 18751 3649
rect 18785 3646 18797 3680
rect 18739 3640 18797 3646
rect 19219 3680 19277 3686
rect 19219 3646 19231 3680
rect 19265 3646 19277 3680
rect 19219 3640 19277 3646
rect 13706 3575 13886 3603
rect 14419 3606 14477 3612
rect 13706 3563 13712 3575
rect 14419 3572 14431 3606
rect 14465 3572 14477 3606
rect 14419 3566 14477 3572
rect 10058 3501 10814 3529
rect 14434 3529 14462 3566
rect 18448 3563 18454 3615
rect 18506 3603 18512 3615
rect 19234 3603 19262 3640
rect 20272 3637 20278 3689
rect 20330 3677 20336 3689
rect 20659 3680 20717 3686
rect 20659 3677 20671 3680
rect 20330 3649 20671 3677
rect 20330 3637 20336 3649
rect 20659 3646 20671 3649
rect 20705 3646 20717 3680
rect 20659 3640 20717 3646
rect 21139 3680 21197 3686
rect 21139 3646 21151 3680
rect 21185 3646 21197 3680
rect 21139 3640 21197 3646
rect 18506 3575 19262 3603
rect 20179 3606 20237 3612
rect 18506 3563 18512 3575
rect 20179 3572 20191 3606
rect 20225 3603 20237 3606
rect 20467 3606 20525 3612
rect 20467 3603 20479 3606
rect 20225 3575 20479 3603
rect 20225 3572 20237 3575
rect 20179 3566 20237 3572
rect 20467 3572 20479 3575
rect 20513 3572 20525 3606
rect 20467 3566 20525 3572
rect 20560 3563 20566 3615
rect 20618 3603 20624 3615
rect 21154 3603 21182 3640
rect 22672 3637 22678 3689
rect 22730 3677 22736 3689
rect 22771 3680 22829 3686
rect 22771 3677 22783 3680
rect 22730 3649 22783 3677
rect 22730 3637 22736 3649
rect 22771 3646 22783 3649
rect 22817 3646 22829 3680
rect 22771 3640 22829 3646
rect 22864 3637 22870 3689
rect 22922 3677 22928 3689
rect 23539 3680 23597 3686
rect 23539 3677 23551 3680
rect 22922 3649 23551 3677
rect 22922 3637 22928 3649
rect 23539 3646 23551 3649
rect 23585 3646 23597 3680
rect 23539 3640 23597 3646
rect 23632 3637 23638 3689
rect 23690 3677 23696 3689
rect 24307 3680 24365 3686
rect 24307 3677 24319 3680
rect 23690 3649 24319 3677
rect 23690 3637 23696 3649
rect 24307 3646 24319 3649
rect 24353 3646 24365 3680
rect 24307 3640 24365 3646
rect 24400 3637 24406 3689
rect 24458 3677 24464 3689
rect 25075 3680 25133 3686
rect 25075 3677 25087 3680
rect 24458 3649 25087 3677
rect 24458 3637 24464 3649
rect 25075 3646 25087 3649
rect 25121 3646 25133 3680
rect 25075 3640 25133 3646
rect 25843 3680 25901 3686
rect 25843 3646 25855 3680
rect 25889 3646 25901 3680
rect 25843 3640 25901 3646
rect 26611 3680 26669 3686
rect 26611 3646 26623 3680
rect 26657 3646 26669 3680
rect 26611 3640 26669 3646
rect 20618 3575 21182 3603
rect 20618 3563 20624 3575
rect 22960 3563 22966 3615
rect 23018 3603 23024 3615
rect 23018 3575 24350 3603
rect 23018 3563 23024 3575
rect 24322 3541 24350 3575
rect 24688 3563 24694 3615
rect 24746 3603 24752 3615
rect 25858 3603 25886 3640
rect 24746 3575 25886 3603
rect 24746 3563 24752 3575
rect 21712 3529 21718 3541
rect 14434 3501 21718 3529
rect 10058 3489 10064 3501
rect 21712 3489 21718 3501
rect 21770 3489 21776 3541
rect 22576 3489 22582 3541
rect 22634 3529 22640 3541
rect 23536 3529 23542 3541
rect 22634 3501 23542 3529
rect 22634 3489 22640 3501
rect 23536 3489 23542 3501
rect 23594 3489 23600 3541
rect 24304 3489 24310 3541
rect 24362 3489 24368 3541
rect 25840 3489 25846 3541
rect 25898 3529 25904 3541
rect 26626 3529 26654 3640
rect 27280 3637 27286 3689
rect 27338 3677 27344 3689
rect 29602 3686 29630 3723
rect 32656 3711 32662 3763
rect 32714 3751 32720 3763
rect 33424 3751 33430 3763
rect 32714 3723 33430 3751
rect 32714 3711 32720 3723
rect 33424 3711 33430 3723
rect 33482 3711 33488 3763
rect 45232 3711 45238 3763
rect 45290 3751 45296 3763
rect 45290 3723 46238 3751
rect 45290 3711 45296 3723
rect 28051 3680 28109 3686
rect 28051 3677 28063 3680
rect 27338 3649 28063 3677
rect 27338 3637 27344 3649
rect 28051 3646 28063 3649
rect 28097 3646 28109 3680
rect 28051 3640 28109 3646
rect 28819 3680 28877 3686
rect 28819 3646 28831 3680
rect 28865 3646 28877 3680
rect 28819 3640 28877 3646
rect 29587 3680 29645 3686
rect 29587 3646 29599 3680
rect 29633 3646 29645 3680
rect 29587 3640 29645 3646
rect 30355 3680 30413 3686
rect 30355 3646 30367 3680
rect 30401 3646 30413 3680
rect 30355 3640 30413 3646
rect 25898 3501 26654 3529
rect 25898 3489 25904 3501
rect 28048 3489 28054 3541
rect 28106 3529 28112 3541
rect 28834 3529 28862 3640
rect 29488 3563 29494 3615
rect 29546 3603 29552 3615
rect 30370 3603 30398 3640
rect 30448 3637 30454 3689
rect 30506 3677 30512 3689
rect 31123 3680 31181 3686
rect 31123 3677 31135 3680
rect 30506 3649 31135 3677
rect 30506 3637 30512 3649
rect 31123 3646 31135 3649
rect 31169 3646 31181 3680
rect 31123 3640 31181 3646
rect 31312 3637 31318 3689
rect 31370 3677 31376 3689
rect 31891 3680 31949 3686
rect 31891 3677 31903 3680
rect 31370 3649 31903 3677
rect 31370 3637 31376 3649
rect 31891 3646 31903 3649
rect 31937 3646 31949 3680
rect 31891 3640 31949 3646
rect 32464 3637 32470 3689
rect 32522 3677 32528 3689
rect 33331 3680 33389 3686
rect 33331 3677 33343 3680
rect 32522 3649 33343 3677
rect 32522 3637 32528 3649
rect 33331 3646 33343 3649
rect 33377 3646 33389 3680
rect 33331 3640 33389 3646
rect 33520 3637 33526 3689
rect 33578 3677 33584 3689
rect 34099 3680 34157 3686
rect 34099 3677 34111 3680
rect 33578 3649 34111 3677
rect 33578 3637 33584 3649
rect 34099 3646 34111 3649
rect 34145 3646 34157 3680
rect 34099 3640 34157 3646
rect 34288 3637 34294 3689
rect 34346 3677 34352 3689
rect 34867 3680 34925 3686
rect 34867 3677 34879 3680
rect 34346 3649 34879 3677
rect 34346 3637 34352 3649
rect 34867 3646 34879 3649
rect 34913 3646 34925 3680
rect 34867 3640 34925 3646
rect 34960 3637 34966 3689
rect 35018 3677 35024 3689
rect 35635 3680 35693 3686
rect 35635 3677 35647 3680
rect 35018 3649 35647 3677
rect 35018 3637 35024 3649
rect 35635 3646 35647 3649
rect 35681 3646 35693 3680
rect 35635 3640 35693 3646
rect 35728 3637 35734 3689
rect 35786 3677 35792 3689
rect 36403 3680 36461 3686
rect 36403 3677 36415 3680
rect 35786 3649 36415 3677
rect 35786 3637 35792 3649
rect 36403 3646 36415 3649
rect 36449 3646 36461 3680
rect 36403 3640 36461 3646
rect 36496 3637 36502 3689
rect 36554 3677 36560 3689
rect 37171 3680 37229 3686
rect 37171 3677 37183 3680
rect 36554 3649 37183 3677
rect 36554 3637 36560 3649
rect 37171 3646 37183 3649
rect 37217 3646 37229 3680
rect 37171 3640 37229 3646
rect 37936 3637 37942 3689
rect 37994 3677 38000 3689
rect 38611 3680 38669 3686
rect 38611 3677 38623 3680
rect 37994 3649 38623 3677
rect 37994 3637 38000 3649
rect 38611 3646 38623 3649
rect 38657 3646 38669 3680
rect 38611 3640 38669 3646
rect 38704 3637 38710 3689
rect 38762 3677 38768 3689
rect 39379 3680 39437 3686
rect 39379 3677 39391 3680
rect 38762 3649 39391 3677
rect 38762 3637 38768 3649
rect 39379 3646 39391 3649
rect 39425 3646 39437 3680
rect 39379 3640 39437 3646
rect 39472 3637 39478 3689
rect 39530 3677 39536 3689
rect 40147 3680 40205 3686
rect 40147 3677 40159 3680
rect 39530 3649 40159 3677
rect 39530 3637 39536 3649
rect 40147 3646 40159 3649
rect 40193 3646 40205 3680
rect 40147 3640 40205 3646
rect 40240 3637 40246 3689
rect 40298 3677 40304 3689
rect 40915 3680 40973 3686
rect 40915 3677 40927 3680
rect 40298 3649 40927 3677
rect 40298 3637 40304 3649
rect 40915 3646 40927 3649
rect 40961 3646 40973 3680
rect 40915 3640 40973 3646
rect 41008 3637 41014 3689
rect 41066 3677 41072 3689
rect 41683 3680 41741 3686
rect 41683 3677 41695 3680
rect 41066 3649 41695 3677
rect 41066 3637 41072 3649
rect 41683 3646 41695 3649
rect 41729 3646 41741 3680
rect 41683 3640 41741 3646
rect 42451 3680 42509 3686
rect 42451 3646 42463 3680
rect 42497 3646 42509 3680
rect 42451 3640 42509 3646
rect 29546 3575 30398 3603
rect 29546 3563 29552 3575
rect 35344 3563 35350 3615
rect 35402 3603 35408 3615
rect 36208 3603 36214 3615
rect 35402 3575 36214 3603
rect 35402 3563 35408 3575
rect 36208 3563 36214 3575
rect 36266 3563 36272 3615
rect 40048 3563 40054 3615
rect 40106 3603 40112 3615
rect 41296 3603 41302 3615
rect 40106 3575 41302 3603
rect 40106 3563 40112 3575
rect 41296 3563 41302 3575
rect 41354 3563 41360 3615
rect 41584 3563 41590 3615
rect 41642 3603 41648 3615
rect 42466 3603 42494 3640
rect 42736 3637 42742 3689
rect 42794 3677 42800 3689
rect 46210 3686 46238 3723
rect 55888 3711 55894 3763
rect 55946 3751 55952 3763
rect 55946 3723 56798 3751
rect 55946 3711 55952 3723
rect 43891 3680 43949 3686
rect 43891 3677 43903 3680
rect 42794 3649 43903 3677
rect 42794 3637 42800 3649
rect 43891 3646 43903 3649
rect 43937 3646 43949 3680
rect 43891 3640 43949 3646
rect 44659 3680 44717 3686
rect 44659 3646 44671 3680
rect 44705 3646 44717 3680
rect 44659 3640 44717 3646
rect 45427 3680 45485 3686
rect 45427 3646 45439 3680
rect 45473 3646 45485 3680
rect 45427 3640 45485 3646
rect 46195 3680 46253 3686
rect 46195 3646 46207 3680
rect 46241 3646 46253 3680
rect 46195 3640 46253 3646
rect 46963 3680 47021 3686
rect 46963 3646 46975 3680
rect 47009 3646 47021 3680
rect 46963 3640 47021 3646
rect 41642 3575 42494 3603
rect 41642 3563 41648 3575
rect 43792 3563 43798 3615
rect 43850 3603 43856 3615
rect 44674 3603 44702 3640
rect 43850 3575 44702 3603
rect 43850 3563 43856 3575
rect 28106 3501 28862 3529
rect 28106 3489 28112 3501
rect 30448 3489 30454 3541
rect 30506 3529 30512 3541
rect 31888 3529 31894 3541
rect 30506 3501 31894 3529
rect 30506 3489 30512 3501
rect 31888 3489 31894 3501
rect 31946 3489 31952 3541
rect 37840 3489 37846 3541
rect 37898 3529 37904 3541
rect 39376 3529 39382 3541
rect 37898 3501 39382 3529
rect 37898 3489 37904 3501
rect 39376 3489 39382 3501
rect 39434 3489 39440 3541
rect 44560 3489 44566 3541
rect 44618 3529 44624 3541
rect 45442 3529 45470 3640
rect 46000 3563 46006 3615
rect 46058 3603 46064 3615
rect 46978 3603 47006 3640
rect 47152 3637 47158 3689
rect 47210 3677 47216 3689
rect 47731 3680 47789 3686
rect 47731 3677 47743 3680
rect 47210 3649 47743 3677
rect 47210 3637 47216 3649
rect 47731 3646 47743 3649
rect 47777 3646 47789 3680
rect 47731 3640 47789 3646
rect 48208 3637 48214 3689
rect 48266 3677 48272 3689
rect 49171 3680 49229 3686
rect 49171 3677 49183 3680
rect 48266 3649 49183 3677
rect 48266 3637 48272 3649
rect 49171 3646 49183 3649
rect 49217 3646 49229 3680
rect 49171 3640 49229 3646
rect 50515 3680 50573 3686
rect 50515 3646 50527 3680
rect 50561 3677 50573 3680
rect 50704 3677 50710 3689
rect 50561 3649 50710 3677
rect 50561 3646 50573 3649
rect 50515 3640 50573 3646
rect 50704 3637 50710 3649
rect 50762 3637 50768 3689
rect 50800 3637 50806 3689
rect 50858 3677 50864 3689
rect 51187 3680 51245 3686
rect 51187 3677 51199 3680
rect 50858 3649 51199 3677
rect 50858 3637 50864 3649
rect 51187 3646 51199 3649
rect 51233 3646 51245 3680
rect 51187 3640 51245 3646
rect 51955 3680 52013 3686
rect 51955 3646 51967 3680
rect 52001 3646 52013 3680
rect 51955 3640 52013 3646
rect 46058 3575 47006 3603
rect 46058 3563 46064 3575
rect 44618 3501 45470 3529
rect 44618 3489 44624 3501
rect 49072 3489 49078 3541
rect 49130 3529 49136 3541
rect 50032 3529 50038 3541
rect 49130 3501 50038 3529
rect 49130 3489 49136 3501
rect 50032 3489 50038 3501
rect 50090 3489 50096 3541
rect 51184 3489 51190 3541
rect 51242 3529 51248 3541
rect 51970 3529 51998 3640
rect 52048 3637 52054 3689
rect 52106 3677 52112 3689
rect 52723 3680 52781 3686
rect 52723 3677 52735 3680
rect 52106 3649 52735 3677
rect 52106 3637 52112 3649
rect 52723 3646 52735 3649
rect 52769 3646 52781 3680
rect 52723 3640 52781 3646
rect 53392 3637 53398 3689
rect 53450 3677 53456 3689
rect 56770 3686 56798 3723
rect 54451 3680 54509 3686
rect 54451 3677 54463 3680
rect 53450 3649 54463 3677
rect 53450 3637 53456 3649
rect 54451 3646 54463 3649
rect 54497 3646 54509 3680
rect 54451 3640 54509 3646
rect 55219 3680 55277 3686
rect 55219 3646 55231 3680
rect 55265 3646 55277 3680
rect 55219 3640 55277 3646
rect 55987 3680 56045 3686
rect 55987 3646 55999 3680
rect 56033 3646 56045 3680
rect 55987 3640 56045 3646
rect 56755 3680 56813 3686
rect 56755 3646 56767 3680
rect 56801 3646 56813 3680
rect 56755 3640 56813 3646
rect 57523 3680 57581 3686
rect 57523 3646 57535 3680
rect 57569 3646 57581 3680
rect 57523 3640 57581 3646
rect 54352 3563 54358 3615
rect 54410 3603 54416 3615
rect 55234 3603 55262 3640
rect 54410 3575 55262 3603
rect 54410 3563 54416 3575
rect 51242 3501 51998 3529
rect 51242 3489 51248 3501
rect 52048 3489 52054 3541
rect 52106 3529 52112 3541
rect 52816 3529 52822 3541
rect 52106 3501 52822 3529
rect 52106 3489 52112 3501
rect 52816 3489 52822 3501
rect 52874 3489 52880 3541
rect 55216 3489 55222 3541
rect 55274 3529 55280 3541
rect 56002 3529 56030 3640
rect 56272 3563 56278 3615
rect 56330 3603 56336 3615
rect 57538 3603 57566 3640
rect 58192 3637 58198 3689
rect 58250 3677 58256 3689
rect 59728 3677 59734 3689
rect 58250 3649 59734 3677
rect 58250 3637 58256 3649
rect 59728 3637 59734 3649
rect 59786 3637 59792 3689
rect 56330 3575 57566 3603
rect 56330 3563 56336 3575
rect 55274 3501 56030 3529
rect 55274 3489 55280 3501
rect 56368 3489 56374 3541
rect 56426 3529 56432 3541
rect 56752 3529 56758 3541
rect 56426 3501 56758 3529
rect 56426 3489 56432 3501
rect 56752 3489 56758 3501
rect 56810 3489 56816 3541
rect 3952 3415 3958 3467
rect 4010 3455 4016 3467
rect 5104 3455 5110 3467
rect 4010 3427 5110 3455
rect 4010 3415 4016 3427
rect 5104 3415 5110 3427
rect 5162 3415 5168 3467
rect 14032 3415 14038 3467
rect 14090 3455 14096 3467
rect 15187 3458 15245 3464
rect 15187 3455 15199 3458
rect 14090 3427 15199 3455
rect 14090 3415 14096 3427
rect 15187 3424 15199 3427
rect 15233 3424 15245 3458
rect 15187 3418 15245 3424
rect 19888 3415 19894 3467
rect 19946 3455 19952 3467
rect 20176 3455 20182 3467
rect 19946 3427 20182 3455
rect 19946 3415 19952 3427
rect 20176 3415 20182 3427
rect 20234 3415 20240 3467
rect 23056 3415 23062 3467
rect 23114 3455 23120 3467
rect 23824 3455 23830 3467
rect 23114 3427 23830 3455
rect 23114 3415 23120 3427
rect 23824 3415 23830 3427
rect 23882 3415 23888 3467
rect 24976 3415 24982 3467
rect 25034 3455 25040 3467
rect 26608 3455 26614 3467
rect 25034 3427 26614 3455
rect 25034 3415 25040 3427
rect 26608 3415 26614 3427
rect 26666 3415 26672 3467
rect 27376 3415 27382 3467
rect 27434 3455 27440 3467
rect 29296 3455 29302 3467
rect 27434 3427 29302 3455
rect 27434 3415 27440 3427
rect 29296 3415 29302 3427
rect 29354 3415 29360 3467
rect 29392 3415 29398 3467
rect 29450 3455 29456 3467
rect 31120 3455 31126 3467
rect 29450 3427 31126 3455
rect 29450 3415 29456 3427
rect 31120 3415 31126 3427
rect 31178 3415 31184 3467
rect 33424 3415 33430 3467
rect 33482 3455 33488 3467
rect 34864 3455 34870 3467
rect 33482 3427 34870 3455
rect 33482 3415 33488 3427
rect 34864 3415 34870 3427
rect 34922 3415 34928 3467
rect 56560 3415 56566 3467
rect 56618 3455 56624 3467
rect 57328 3455 57334 3467
rect 56618 3427 57334 3455
rect 56618 3415 56624 3427
rect 57328 3415 57334 3427
rect 57386 3415 57392 3467
rect 1152 3356 58848 3378
rect 1152 3304 19654 3356
rect 19706 3304 19718 3356
rect 19770 3304 19782 3356
rect 19834 3304 19846 3356
rect 19898 3304 50374 3356
rect 50426 3304 50438 3356
rect 50490 3304 50502 3356
rect 50554 3304 50566 3356
rect 50618 3304 58848 3356
rect 1152 3282 58848 3304
rect 592 3193 598 3245
rect 650 3233 656 3245
rect 1456 3233 1462 3245
rect 650 3205 1462 3233
rect 650 3193 656 3205
rect 1456 3193 1462 3205
rect 1514 3193 1520 3245
rect 2416 3193 2422 3245
rect 2474 3233 2480 3245
rect 5200 3233 5206 3245
rect 2474 3205 5206 3233
rect 2474 3193 2480 3205
rect 5200 3193 5206 3205
rect 5258 3193 5264 3245
rect 9424 3193 9430 3245
rect 9482 3233 9488 3245
rect 10672 3233 10678 3245
rect 9482 3205 10678 3233
rect 9482 3193 9488 3205
rect 10672 3193 10678 3205
rect 10730 3193 10736 3245
rect 12208 3193 12214 3245
rect 12266 3233 12272 3245
rect 12976 3233 12982 3245
rect 12266 3205 12982 3233
rect 12266 3193 12272 3205
rect 12976 3193 12982 3205
rect 13034 3193 13040 3245
rect 19696 3193 19702 3245
rect 19754 3233 19760 3245
rect 20368 3233 20374 3245
rect 19754 3205 20374 3233
rect 19754 3193 19760 3205
rect 20368 3193 20374 3205
rect 20426 3193 20432 3245
rect 21616 3233 21622 3245
rect 21577 3205 21622 3233
rect 21616 3193 21622 3205
rect 21674 3193 21680 3245
rect 21712 3193 21718 3245
rect 21770 3233 21776 3245
rect 41200 3233 41206 3245
rect 21770 3205 41206 3233
rect 21770 3193 21776 3205
rect 41200 3193 41206 3205
rect 41258 3193 41264 3245
rect 42160 3193 42166 3245
rect 42218 3233 42224 3245
rect 43888 3233 43894 3245
rect 42218 3205 43894 3233
rect 42218 3193 42224 3205
rect 43888 3193 43894 3205
rect 43946 3193 43952 3245
rect 45136 3193 45142 3245
rect 45194 3233 45200 3245
rect 46480 3233 46486 3245
rect 45194 3205 46486 3233
rect 45194 3193 45200 3205
rect 46480 3193 46486 3205
rect 46538 3193 46544 3245
rect 56848 3193 56854 3245
rect 56906 3233 56912 3245
rect 58000 3233 58006 3245
rect 56906 3205 58006 3233
rect 56906 3193 56912 3205
rect 58000 3193 58006 3205
rect 58058 3193 58064 3245
rect 3472 3119 3478 3171
rect 3530 3159 3536 3171
rect 4912 3159 4918 3171
rect 3530 3131 4918 3159
rect 3530 3119 3536 3131
rect 4912 3119 4918 3131
rect 4970 3119 4976 3171
rect 5104 3119 5110 3171
rect 5162 3159 5168 3171
rect 5968 3159 5974 3171
rect 5162 3131 5974 3159
rect 5162 3119 5168 3131
rect 5968 3119 5974 3131
rect 6026 3119 6032 3171
rect 6160 3119 6166 3171
rect 6218 3159 6224 3171
rect 19891 3162 19949 3168
rect 19891 3159 19903 3162
rect 6218 3131 17918 3159
rect 6218 3119 6224 3131
rect 1456 3045 1462 3097
rect 1514 3085 1520 3097
rect 2128 3085 2134 3097
rect 1514 3057 2134 3085
rect 1514 3045 1520 3057
rect 2128 3045 2134 3057
rect 2186 3045 2192 3097
rect 6832 3045 6838 3097
rect 6890 3085 6896 3097
rect 7696 3085 7702 3097
rect 6890 3057 7702 3085
rect 6890 3045 6896 3057
rect 7696 3045 7702 3057
rect 7754 3045 7760 3097
rect 8944 3045 8950 3097
rect 9002 3085 9008 3097
rect 15283 3088 15341 3094
rect 15283 3085 15295 3088
rect 9002 3057 10526 3085
rect 9002 3045 9008 3057
rect 16 2971 22 3023
rect 74 3011 80 3023
rect 1555 3014 1613 3020
rect 1555 3011 1567 3014
rect 74 2983 1567 3011
rect 74 2971 80 2983
rect 1555 2980 1567 2983
rect 1601 2980 1613 3014
rect 2323 3014 2381 3020
rect 2323 3011 2335 3014
rect 1555 2974 1613 2980
rect 1666 2983 2335 3011
rect 688 2897 694 2949
rect 746 2937 752 2949
rect 1666 2937 1694 2983
rect 2323 2980 2335 2983
rect 2369 2980 2381 3014
rect 2323 2974 2381 2980
rect 3091 3014 3149 3020
rect 3091 2980 3103 3014
rect 3137 2980 3149 3014
rect 4912 3011 4918 3023
rect 4873 2983 4918 3011
rect 3091 2974 3149 2980
rect 746 2909 1694 2937
rect 746 2897 752 2909
rect 2128 2897 2134 2949
rect 2186 2937 2192 2949
rect 3106 2937 3134 2974
rect 4912 2971 4918 2983
rect 4970 2971 4976 3023
rect 5200 2971 5206 3023
rect 5258 3011 5264 3023
rect 5683 3014 5741 3020
rect 5683 3011 5695 3014
rect 5258 2983 5695 3011
rect 5258 2971 5264 2983
rect 5683 2980 5695 2983
rect 5729 2980 5741 3014
rect 5683 2974 5741 2980
rect 5968 2971 5974 3023
rect 6026 3011 6032 3023
rect 7027 3014 7085 3020
rect 7027 3011 7039 3014
rect 6026 2983 7039 3011
rect 6026 2971 6032 2983
rect 7027 2980 7039 2983
rect 7073 2980 7085 3014
rect 7795 3014 7853 3020
rect 7795 3011 7807 3014
rect 7027 2974 7085 2980
rect 7186 2983 7807 3011
rect 2186 2909 3134 2937
rect 2186 2897 2192 2909
rect 6736 2897 6742 2949
rect 6794 2937 6800 2949
rect 7186 2937 7214 2983
rect 7795 2980 7807 2983
rect 7841 2980 7853 3014
rect 7795 2974 7853 2980
rect 8176 2971 8182 3023
rect 8234 3011 8240 3023
rect 10498 3020 10526 3057
rect 12946 3057 15295 3085
rect 9715 3014 9773 3020
rect 9715 3011 9727 3014
rect 8234 2983 9727 3011
rect 8234 2971 8240 2983
rect 9715 2980 9727 2983
rect 9761 2980 9773 3014
rect 9715 2974 9773 2980
rect 10483 3014 10541 3020
rect 10483 2980 10495 3014
rect 10529 2980 10541 3014
rect 10483 2974 10541 2980
rect 6794 2909 7214 2937
rect 6794 2897 6800 2909
rect 7696 2897 7702 2949
rect 7754 2937 7760 2949
rect 7984 2937 7990 2949
rect 7754 2909 7990 2937
rect 7754 2897 7760 2909
rect 7984 2897 7990 2909
rect 8042 2897 8048 2949
rect 9808 2897 9814 2949
rect 9866 2937 9872 2949
rect 10192 2937 10198 2949
rect 9866 2909 10198 2937
rect 9866 2897 9872 2909
rect 10192 2897 10198 2909
rect 10250 2897 10256 2949
rect 11536 2897 11542 2949
rect 11594 2937 11600 2949
rect 12946 2937 12974 3057
rect 15283 3054 15295 3057
rect 15329 3054 15341 3088
rect 17890 3085 17918 3131
rect 18754 3131 19903 3159
rect 18754 3085 18782 3131
rect 19891 3128 19903 3131
rect 19937 3128 19949 3162
rect 19891 3122 19949 3128
rect 22384 3119 22390 3171
rect 22442 3159 22448 3171
rect 23152 3159 23158 3171
rect 22442 3131 23158 3159
rect 22442 3119 22448 3131
rect 23152 3119 23158 3131
rect 23210 3119 23216 3171
rect 51379 3162 51437 3168
rect 51379 3159 51391 3162
rect 23266 3131 51391 3159
rect 17890 3057 18782 3085
rect 18835 3088 18893 3094
rect 15283 3048 15341 3054
rect 18835 3054 18847 3088
rect 18881 3085 18893 3088
rect 18928 3085 18934 3097
rect 18881 3057 18934 3085
rect 18881 3054 18893 3057
rect 18835 3048 18893 3054
rect 18928 3045 18934 3057
rect 18986 3045 18992 3097
rect 19426 3057 21374 3085
rect 13072 2971 13078 3023
rect 13130 3011 13136 3023
rect 13363 3014 13421 3020
rect 13363 3011 13375 3014
rect 13130 2983 13375 3011
rect 13130 2971 13136 2983
rect 13363 2980 13375 2983
rect 13409 2980 13421 3014
rect 13363 2974 13421 2980
rect 13939 3014 13997 3020
rect 13939 2980 13951 3014
rect 13985 3011 13997 3014
rect 14032 3011 14038 3023
rect 13985 2983 14038 3011
rect 13985 2980 13997 2983
rect 13939 2974 13997 2980
rect 14032 2971 14038 2983
rect 14090 2971 14096 3023
rect 14800 2971 14806 3023
rect 14858 3011 14864 3023
rect 15475 3014 15533 3020
rect 15475 3011 15487 3014
rect 14858 2983 15487 3011
rect 14858 2971 14864 2983
rect 15475 2980 15487 2983
rect 15521 2980 15533 3014
rect 16624 3011 16630 3023
rect 16585 2983 16630 3011
rect 15475 2974 15533 2980
rect 16624 2971 16630 2983
rect 16682 2971 16688 3023
rect 17008 2971 17014 3023
rect 17066 3011 17072 3023
rect 18163 3014 18221 3020
rect 18163 3011 18175 3014
rect 17066 2983 18175 3011
rect 17066 2971 17072 2983
rect 18163 2980 18175 2983
rect 18209 2980 18221 3014
rect 18163 2974 18221 2980
rect 19027 3014 19085 3020
rect 19027 2980 19039 3014
rect 19073 2980 19085 3014
rect 19027 2974 19085 2980
rect 11594 2909 12974 2937
rect 13171 2940 13229 2946
rect 11594 2897 11600 2909
rect 13171 2906 13183 2940
rect 13217 2937 13229 2940
rect 13744 2937 13750 2949
rect 13217 2909 13750 2937
rect 13217 2906 13229 2909
rect 13171 2900 13229 2906
rect 13744 2897 13750 2909
rect 13802 2897 13808 2949
rect 17776 2897 17782 2949
rect 17834 2937 17840 2949
rect 17971 2940 18029 2946
rect 17971 2937 17983 2940
rect 17834 2909 17983 2937
rect 17834 2897 17840 2909
rect 17971 2906 17983 2909
rect 18017 2906 18029 2940
rect 19042 2937 19070 2974
rect 19312 2937 19318 2949
rect 17971 2900 18029 2906
rect 18178 2909 19070 2937
rect 19138 2909 19318 2937
rect 17680 2823 17686 2875
rect 17738 2863 17744 2875
rect 18178 2863 18206 2909
rect 17738 2835 18206 2863
rect 17738 2823 17744 2835
rect 18928 2823 18934 2875
rect 18986 2863 18992 2875
rect 19138 2863 19166 2909
rect 19312 2897 19318 2909
rect 19370 2897 19376 2949
rect 18986 2835 19166 2863
rect 18986 2823 18992 2835
rect 19312 2749 19318 2801
rect 19370 2789 19376 2801
rect 19426 2789 19454 3057
rect 21346 3020 21374 3057
rect 21616 3045 21622 3097
rect 21674 3085 21680 3097
rect 22480 3085 22486 3097
rect 21674 3057 22486 3085
rect 21674 3045 21680 3057
rect 22480 3045 22486 3057
rect 22538 3045 22544 3097
rect 23266 3085 23294 3131
rect 51379 3128 51391 3131
rect 51425 3159 51437 3162
rect 51425 3131 51614 3159
rect 51425 3128 51437 3131
rect 51379 3122 51437 3128
rect 22594 3057 23294 3085
rect 20851 3014 20909 3020
rect 20851 3011 20863 3014
rect 20002 2983 20863 3011
rect 20002 2894 20030 2983
rect 20851 2980 20863 2983
rect 20897 2980 20909 3014
rect 20851 2974 20909 2980
rect 21331 3014 21389 3020
rect 21331 2980 21343 3014
rect 21377 2980 21389 3014
rect 21331 2974 21389 2980
rect 21715 3014 21773 3020
rect 21715 2980 21727 3014
rect 21761 3011 21773 3014
rect 22594 3011 22622 3057
rect 31888 3045 31894 3097
rect 31946 3085 31952 3097
rect 33328 3085 33334 3097
rect 31946 3057 33334 3085
rect 31946 3045 31952 3057
rect 33328 3045 33334 3057
rect 33386 3045 33392 3097
rect 41107 3088 41165 3094
rect 41107 3054 41119 3088
rect 41153 3085 41165 3088
rect 42448 3085 42454 3097
rect 41153 3057 42454 3085
rect 41153 3054 41165 3057
rect 41107 3048 41165 3054
rect 42448 3045 42454 3057
rect 42506 3045 42512 3097
rect 42928 3045 42934 3097
rect 42986 3085 42992 3097
rect 43984 3085 43990 3097
rect 42986 3057 43990 3085
rect 42986 3045 42992 3057
rect 43984 3045 43990 3057
rect 44042 3045 44048 3097
rect 44083 3088 44141 3094
rect 44083 3054 44095 3088
rect 44129 3085 44141 3088
rect 44368 3085 44374 3097
rect 44129 3057 44374 3085
rect 44129 3054 44141 3057
rect 44083 3048 44141 3054
rect 44368 3045 44374 3057
rect 44426 3045 44432 3097
rect 45328 3045 45334 3097
rect 45386 3085 45392 3097
rect 51586 3094 51614 3131
rect 46387 3088 46445 3094
rect 46387 3085 46399 3088
rect 45386 3057 46399 3085
rect 45386 3045 45392 3057
rect 46387 3054 46399 3057
rect 46433 3054 46445 3088
rect 46387 3048 46445 3054
rect 51571 3088 51629 3094
rect 51571 3054 51583 3088
rect 51617 3054 51629 3088
rect 51571 3048 51629 3054
rect 21761 2983 22622 3011
rect 22675 3014 22733 3020
rect 21761 2980 21773 2983
rect 21715 2974 21773 2980
rect 22675 2980 22687 3014
rect 22721 3011 22733 3014
rect 23155 3014 23213 3020
rect 23155 3011 23167 3014
rect 22721 2983 23167 3011
rect 22721 2980 22733 2983
rect 22675 2974 22733 2980
rect 23155 2980 23167 2983
rect 23201 2980 23213 3014
rect 23155 2974 23213 2980
rect 23923 3014 23981 3020
rect 23923 2980 23935 3014
rect 23969 2980 23981 3014
rect 23923 2974 23981 2980
rect 20656 2937 20662 2949
rect 20617 2909 20662 2937
rect 20656 2897 20662 2909
rect 20714 2897 20720 2949
rect 21424 2897 21430 2949
rect 21482 2937 21488 2949
rect 22387 2940 22445 2946
rect 22387 2937 22399 2940
rect 21482 2909 22399 2937
rect 21482 2897 21488 2909
rect 22387 2906 22399 2909
rect 22433 2906 22445 2940
rect 22387 2900 22445 2906
rect 22480 2897 22486 2949
rect 22538 2937 22544 2949
rect 23938 2937 23966 2974
rect 24016 2971 24022 3023
rect 24074 3011 24080 3023
rect 25843 3014 25901 3020
rect 25843 3011 25855 3014
rect 24074 2983 25855 3011
rect 24074 2971 24080 2983
rect 25843 2980 25855 2983
rect 25889 2980 25901 3014
rect 25843 2974 25901 2980
rect 26611 3014 26669 3020
rect 26611 2980 26623 3014
rect 26657 2980 26669 3014
rect 26611 2974 26669 2980
rect 22538 2909 23966 2937
rect 22538 2897 22544 2909
rect 25072 2897 25078 2949
rect 25130 2937 25136 2949
rect 26626 2937 26654 2974
rect 26896 2971 26902 3023
rect 26954 3011 26960 3023
rect 28531 3014 28589 3020
rect 28531 3011 28543 3014
rect 26954 2983 28543 3011
rect 26954 2971 26960 2983
rect 28531 2980 28543 2983
rect 28577 2980 28589 3014
rect 28531 2974 28589 2980
rect 29299 3014 29357 3020
rect 29299 2980 29311 3014
rect 29345 2980 29357 3014
rect 29299 2974 29357 2980
rect 25130 2909 26654 2937
rect 25130 2897 25136 2909
rect 27664 2897 27670 2949
rect 27722 2937 27728 2949
rect 29314 2937 29342 2974
rect 29872 2971 29878 3023
rect 29930 3011 29936 3023
rect 31219 3014 31277 3020
rect 31219 3011 31231 3014
rect 29930 2983 31231 3011
rect 29930 2971 29936 2983
rect 31219 2980 31231 2983
rect 31265 2980 31277 3014
rect 31219 2974 31277 2980
rect 31987 3014 32045 3020
rect 31987 2980 31999 3014
rect 32033 2980 32045 3014
rect 31987 2974 32045 2980
rect 29776 2937 29782 2949
rect 27722 2909 29342 2937
rect 29410 2909 29782 2937
rect 27722 2897 27728 2909
rect 19906 2866 20030 2894
rect 20083 2866 20141 2872
rect 19906 2801 19934 2866
rect 20083 2832 20095 2866
rect 20129 2863 20141 2866
rect 21715 2866 21773 2872
rect 21715 2863 21727 2866
rect 20129 2835 21727 2863
rect 20129 2832 20141 2835
rect 20083 2826 20141 2832
rect 21715 2832 21727 2835
rect 21761 2832 21773 2866
rect 21715 2826 21773 2832
rect 28912 2823 28918 2875
rect 28970 2863 28976 2875
rect 29410 2863 29438 2909
rect 29776 2897 29782 2909
rect 29834 2897 29840 2949
rect 30544 2897 30550 2949
rect 30602 2937 30608 2949
rect 32002 2937 32030 2974
rect 32080 2971 32086 3023
rect 32138 3011 32144 3023
rect 33907 3014 33965 3020
rect 33907 3011 33919 3014
rect 32138 2983 33919 3011
rect 32138 2971 32144 2983
rect 33907 2980 33919 2983
rect 33953 2980 33965 3014
rect 33907 2974 33965 2980
rect 34675 3014 34733 3020
rect 34675 2980 34687 3014
rect 34721 2980 34733 3014
rect 34675 2974 34733 2980
rect 30602 2909 32030 2937
rect 30602 2897 30608 2909
rect 32272 2897 32278 2949
rect 32330 2937 32336 2949
rect 33136 2937 33142 2949
rect 32330 2909 33142 2937
rect 32330 2897 32336 2909
rect 33136 2897 33142 2909
rect 33194 2897 33200 2949
rect 33328 2897 33334 2949
rect 33386 2937 33392 2949
rect 34690 2937 34718 2974
rect 35440 2971 35446 3023
rect 35498 3011 35504 3023
rect 36595 3014 36653 3020
rect 36595 3011 36607 3014
rect 35498 2983 36607 3011
rect 35498 2971 35504 2983
rect 36595 2980 36607 2983
rect 36641 2980 36653 3014
rect 36595 2974 36653 2980
rect 37363 3014 37421 3020
rect 37363 2980 37375 3014
rect 37409 2980 37421 3014
rect 37363 2974 37421 2980
rect 33386 2909 34718 2937
rect 33386 2897 33392 2909
rect 36208 2897 36214 2949
rect 36266 2937 36272 2949
rect 37378 2937 37406 2974
rect 37552 2971 37558 3023
rect 37610 3011 37616 3023
rect 39283 3014 39341 3020
rect 39283 3011 39295 3014
rect 37610 2983 39295 3011
rect 37610 2971 37616 2983
rect 39283 2980 39295 2983
rect 39329 2980 39341 3014
rect 39283 2974 39341 2980
rect 40051 3014 40109 3020
rect 40051 2980 40063 3014
rect 40097 2980 40109 3014
rect 40051 2974 40109 2980
rect 36266 2909 37406 2937
rect 36266 2897 36272 2909
rect 38320 2897 38326 2949
rect 38378 2937 38384 2949
rect 40066 2937 40094 2974
rect 40528 2971 40534 3023
rect 40586 3011 40592 3023
rect 41971 3014 42029 3020
rect 41971 3011 41983 3014
rect 40586 2983 41983 3011
rect 40586 2971 40592 2983
rect 41971 2980 41983 2983
rect 42017 2980 42029 3014
rect 41971 2974 42029 2980
rect 42739 3014 42797 3020
rect 42739 2980 42751 3014
rect 42785 2980 42797 3014
rect 42739 2974 42797 2980
rect 41104 2937 41110 2949
rect 38378 2909 40094 2937
rect 41065 2909 41110 2937
rect 38378 2897 38384 2909
rect 41104 2897 41110 2909
rect 41162 2897 41168 2949
rect 41200 2897 41206 2949
rect 41258 2937 41264 2949
rect 42754 2937 42782 2974
rect 43024 2971 43030 3023
rect 43082 3011 43088 3023
rect 44659 3014 44717 3020
rect 44659 3011 44671 3014
rect 43082 2983 44671 3011
rect 43082 2971 43088 2983
rect 44659 2980 44671 2983
rect 44705 2980 44717 3014
rect 44659 2974 44717 2980
rect 45427 3014 45485 3020
rect 45427 2980 45439 3014
rect 45473 2980 45485 3014
rect 45427 2974 45485 2980
rect 41258 2909 42782 2937
rect 41258 2897 41264 2909
rect 43888 2897 43894 2949
rect 43946 2937 43952 2949
rect 44083 2940 44141 2946
rect 44083 2937 44095 2940
rect 43946 2909 44095 2937
rect 43946 2897 43952 2909
rect 44083 2906 44095 2909
rect 44129 2906 44141 2940
rect 44083 2900 44141 2906
rect 44176 2897 44182 2949
rect 44234 2937 44240 2949
rect 45442 2937 45470 2974
rect 45616 2971 45622 3023
rect 45674 3011 45680 3023
rect 47347 3014 47405 3020
rect 47347 3011 47359 3014
rect 45674 2983 47359 3011
rect 45674 2971 45680 2983
rect 47347 2980 47359 2983
rect 47393 2980 47405 3014
rect 47347 2974 47405 2980
rect 48115 3014 48173 3020
rect 48115 2980 48127 3014
rect 48161 2980 48173 3014
rect 48115 2974 48173 2980
rect 44234 2909 45470 2937
rect 44234 2897 44240 2909
rect 46384 2897 46390 2949
rect 46442 2937 46448 2949
rect 48130 2937 48158 2974
rect 49648 2971 49654 3023
rect 49706 3011 49712 3023
rect 50035 3014 50093 3020
rect 50035 3011 50047 3014
rect 49706 2983 50047 3011
rect 49706 2971 49712 2983
rect 50035 2980 50047 2983
rect 50081 2980 50093 3014
rect 50035 2974 50093 2980
rect 50803 3014 50861 3020
rect 50803 2980 50815 3014
rect 50849 2980 50861 3014
rect 50803 2974 50861 2980
rect 46442 2909 48158 2937
rect 46442 2897 46448 2909
rect 49936 2897 49942 2949
rect 49994 2937 50000 2949
rect 50818 2937 50846 2974
rect 51472 2971 51478 3023
rect 51530 3011 51536 3023
rect 52723 3014 52781 3020
rect 52723 3011 52735 3014
rect 51530 2983 52735 3011
rect 51530 2971 51536 2983
rect 52723 2980 52735 2983
rect 52769 2980 52781 3014
rect 53491 3014 53549 3020
rect 53491 3011 53503 3014
rect 52723 2974 52781 2980
rect 52834 2983 53503 3011
rect 49994 2909 50846 2937
rect 49994 2897 50000 2909
rect 52240 2897 52246 2949
rect 52298 2937 52304 2949
rect 52834 2937 52862 2983
rect 53491 2980 53503 2983
rect 53537 2980 53549 3014
rect 53491 2974 53549 2980
rect 53776 2971 53782 3023
rect 53834 3011 53840 3023
rect 55411 3014 55469 3020
rect 55411 3011 55423 3014
rect 53834 2983 55423 3011
rect 53834 2971 53840 2983
rect 55411 2980 55423 2983
rect 55457 2980 55469 3014
rect 55411 2974 55469 2980
rect 56179 3014 56237 3020
rect 56179 2980 56191 3014
rect 56225 2980 56237 3014
rect 56179 2974 56237 2980
rect 52298 2909 52862 2937
rect 52298 2897 52304 2909
rect 52912 2897 52918 2949
rect 52970 2937 52976 2949
rect 53680 2937 53686 2949
rect 52970 2909 53686 2937
rect 52970 2897 52976 2909
rect 53680 2897 53686 2909
rect 53738 2897 53744 2949
rect 54832 2897 54838 2949
rect 54890 2937 54896 2949
rect 56194 2937 56222 2974
rect 54890 2909 56222 2937
rect 54890 2897 54896 2909
rect 57712 2897 57718 2949
rect 57770 2937 57776 2949
rect 59440 2937 59446 2949
rect 57770 2909 59446 2937
rect 57770 2897 57776 2909
rect 59440 2897 59446 2909
rect 59498 2897 59504 2949
rect 28970 2835 29438 2863
rect 28970 2823 28976 2835
rect 35632 2823 35638 2875
rect 35690 2863 35696 2875
rect 36880 2863 36886 2875
rect 35690 2835 36886 2863
rect 35690 2823 35696 2835
rect 36880 2823 36886 2835
rect 36938 2823 36944 2875
rect 37264 2823 37270 2875
rect 37322 2863 37328 2875
rect 57139 2866 57197 2872
rect 57139 2863 57151 2866
rect 37322 2835 57151 2863
rect 37322 2823 37328 2835
rect 57139 2832 57151 2835
rect 57185 2832 57197 2866
rect 57139 2826 57197 2832
rect 19370 2761 19454 2789
rect 19370 2749 19376 2761
rect 19888 2749 19894 2801
rect 19946 2749 19952 2801
rect 24880 2789 24886 2801
rect 24841 2761 24886 2789
rect 24880 2749 24886 2761
rect 24938 2749 24944 2801
rect 35248 2749 35254 2801
rect 35306 2789 35312 2801
rect 42448 2789 42454 2801
rect 35306 2761 42454 2789
rect 35306 2749 35312 2761
rect 42448 2749 42454 2761
rect 42506 2749 42512 2801
rect 44656 2749 44662 2801
rect 44714 2789 44720 2801
rect 45040 2789 45046 2801
rect 44714 2761 45046 2789
rect 44714 2749 44720 2761
rect 45040 2749 45046 2761
rect 45098 2749 45104 2801
rect 54448 2789 54454 2801
rect 54409 2761 54454 2789
rect 54448 2749 54454 2761
rect 54506 2749 54512 2801
rect 1152 2690 58848 2712
rect 1152 2638 4294 2690
rect 4346 2638 4358 2690
rect 4410 2638 4422 2690
rect 4474 2638 4486 2690
rect 4538 2638 35014 2690
rect 35066 2638 35078 2690
rect 35130 2638 35142 2690
rect 35194 2638 35206 2690
rect 35258 2638 58848 2690
rect 1152 2616 58848 2638
rect 3952 2527 3958 2579
rect 4010 2567 4016 2579
rect 4240 2567 4246 2579
rect 4010 2539 4246 2567
rect 4010 2527 4016 2539
rect 4240 2527 4246 2539
rect 4298 2527 4304 2579
rect 4336 2527 4342 2579
rect 4394 2567 4400 2579
rect 4816 2567 4822 2579
rect 4394 2539 4822 2567
rect 4394 2527 4400 2539
rect 4816 2527 4822 2539
rect 4874 2527 4880 2579
rect 20176 2527 20182 2579
rect 20234 2567 20240 2579
rect 21232 2567 21238 2579
rect 20234 2539 21238 2567
rect 20234 2527 20240 2539
rect 21232 2527 21238 2539
rect 21290 2527 21296 2579
rect 35152 2527 35158 2579
rect 35210 2567 35216 2579
rect 35536 2567 35542 2579
rect 35210 2539 35542 2567
rect 35210 2527 35216 2539
rect 35536 2527 35542 2539
rect 35594 2527 35600 2579
rect 42448 2527 42454 2579
rect 42506 2567 42512 2579
rect 54448 2567 54454 2579
rect 42506 2539 54454 2567
rect 42506 2527 42512 2539
rect 54448 2527 54454 2539
rect 54506 2527 54512 2579
rect 24880 2453 24886 2505
rect 24938 2493 24944 2505
rect 52816 2493 52822 2505
rect 24938 2465 52822 2493
rect 24938 2453 24944 2465
rect 52816 2453 52822 2465
rect 52874 2453 52880 2505
rect 34096 2379 34102 2431
rect 34154 2419 34160 2431
rect 37264 2419 37270 2431
rect 34154 2391 37270 2419
rect 34154 2379 34160 2391
rect 37264 2379 37270 2391
rect 37322 2379 37328 2431
rect 45040 2379 45046 2431
rect 45098 2419 45104 2431
rect 45808 2419 45814 2431
rect 45098 2391 45814 2419
rect 45098 2379 45104 2391
rect 45808 2379 45814 2391
rect 45866 2379 45872 2431
rect 4720 2009 4726 2061
rect 4778 2049 4784 2061
rect 5296 2049 5302 2061
rect 4778 2021 5302 2049
rect 4778 2009 4784 2021
rect 5296 2009 5302 2021
rect 5354 2009 5360 2061
rect 4528 1861 4534 1913
rect 4586 1901 4592 1913
rect 4816 1901 4822 1913
rect 4586 1873 4822 1901
rect 4586 1861 4592 1873
rect 4816 1861 4822 1873
rect 4874 1861 4880 1913
rect 18064 1861 18070 1913
rect 18122 1901 18128 1913
rect 18256 1901 18262 1913
rect 18122 1873 18262 1901
rect 18122 1861 18128 1873
rect 18256 1861 18262 1873
rect 18314 1861 18320 1913
rect 13072 1713 13078 1765
rect 13130 1753 13136 1765
rect 13264 1753 13270 1765
rect 13130 1725 13270 1753
rect 13130 1713 13136 1725
rect 13264 1713 13270 1725
rect 13322 1713 13328 1765
rect 30352 1713 30358 1765
rect 30410 1753 30416 1765
rect 30640 1753 30646 1765
rect 30410 1725 30646 1753
rect 30410 1713 30416 1725
rect 30640 1713 30646 1725
rect 30698 1713 30704 1765
rect 34864 1713 34870 1765
rect 34922 1753 34928 1765
rect 35920 1753 35926 1765
rect 34922 1725 35926 1753
rect 34922 1713 34928 1725
rect 35920 1713 35926 1725
rect 35978 1713 35984 1765
rect 39952 1713 39958 1765
rect 40010 1753 40016 1765
rect 40240 1753 40246 1765
rect 40010 1725 40246 1753
rect 40010 1713 40016 1725
rect 40240 1713 40246 1725
rect 40298 1713 40304 1765
rect 50704 1713 50710 1765
rect 50762 1753 50768 1765
rect 50896 1753 50902 1765
rect 50762 1725 50902 1753
rect 50762 1713 50768 1725
rect 50896 1713 50902 1725
rect 50954 1713 50960 1765
rect 54352 1713 54358 1765
rect 54410 1753 54416 1765
rect 54640 1753 54646 1765
rect 54410 1725 54646 1753
rect 54410 1713 54416 1725
rect 54640 1713 54646 1725
rect 54698 1713 54704 1765
rect 50512 1639 50518 1691
rect 50570 1679 50576 1691
rect 51088 1679 51094 1691
rect 50570 1651 51094 1679
rect 50570 1639 50576 1651
rect 51088 1639 51094 1651
rect 51146 1639 51152 1691
rect 20464 1565 20470 1617
rect 20522 1605 20528 1617
rect 20848 1605 20854 1617
rect 20522 1577 20854 1605
rect 20522 1565 20528 1577
rect 20848 1565 20854 1577
rect 20906 1565 20912 1617
rect 22096 1565 22102 1617
rect 22154 1605 22160 1617
rect 22672 1605 22678 1617
rect 22154 1577 22678 1605
rect 22154 1565 22160 1577
rect 22672 1565 22678 1577
rect 22730 1565 22736 1617
rect 50896 1565 50902 1617
rect 50954 1605 50960 1617
rect 51568 1605 51574 1617
rect 50954 1577 51574 1605
rect 50954 1565 50960 1577
rect 51568 1565 51574 1577
rect 51626 1565 51632 1617
rect 36304 1491 36310 1543
rect 36362 1491 36368 1543
rect 19312 1417 19318 1469
rect 19370 1457 19376 1469
rect 19984 1457 19990 1469
rect 19370 1429 19990 1457
rect 19370 1417 19376 1429
rect 19984 1417 19990 1429
rect 20042 1417 20048 1469
rect 33232 1417 33238 1469
rect 33290 1457 33296 1469
rect 33712 1457 33718 1469
rect 33290 1429 33718 1457
rect 33290 1417 33296 1429
rect 33712 1417 33718 1429
rect 33770 1417 33776 1469
rect 36322 1173 36350 1491
rect 36304 1121 36310 1173
rect 36362 1121 36368 1173
<< via1 >>
rect 4294 57250 4346 57302
rect 4358 57250 4410 57302
rect 4422 57250 4474 57302
rect 4486 57250 4538 57302
rect 35014 57250 35066 57302
rect 35078 57250 35130 57302
rect 35142 57250 35194 57302
rect 35206 57250 35258 57302
rect 16438 57065 16490 57117
rect 15958 56991 16010 57043
rect 17494 56991 17546 57043
rect 19126 56991 19178 57043
rect 29110 56991 29162 57043
rect 57046 57034 57098 57043
rect 57046 57000 57055 57034
rect 57055 57000 57089 57034
rect 57089 57000 57098 57034
rect 57046 56991 57098 57000
rect 214 56917 266 56969
rect 1750 56917 1802 56969
rect 3286 56917 3338 56969
rect 4918 56960 4970 56969
rect 4918 56926 4927 56960
rect 4927 56926 4961 56960
rect 4961 56926 4970 56960
rect 4918 56917 4970 56926
rect 6454 56917 6506 56969
rect 8086 56960 8138 56969
rect 8086 56926 8095 56960
rect 8095 56926 8129 56960
rect 8129 56926 8138 56960
rect 8086 56917 8138 56926
rect 9622 56917 9674 56969
rect 11254 56960 11306 56969
rect 11254 56926 11263 56960
rect 11263 56926 11297 56960
rect 11297 56926 11306 56960
rect 11254 56917 11306 56926
rect 12790 56960 12842 56969
rect 12790 56926 12799 56960
rect 12799 56926 12833 56960
rect 12833 56926 12842 56960
rect 12790 56917 12842 56926
rect 14422 56917 14474 56969
rect 20662 56917 20714 56969
rect 22294 56917 22346 56969
rect 23830 56917 23882 56969
rect 25462 56917 25514 56969
rect 26998 56960 27050 56969
rect 26998 56926 27007 56960
rect 27007 56926 27041 56960
rect 27041 56926 27050 56960
rect 26998 56917 27050 56926
rect 28630 56960 28682 56969
rect 28630 56926 28639 56960
rect 28639 56926 28673 56960
rect 28673 56926 28682 56960
rect 28630 56917 28682 56926
rect 30166 56917 30218 56969
rect 31702 56960 31754 56969
rect 31702 56926 31711 56960
rect 31711 56926 31745 56960
rect 31745 56926 31754 56960
rect 31702 56917 31754 56926
rect 33334 56917 33386 56969
rect 34870 56960 34922 56969
rect 34870 56926 34879 56960
rect 34879 56926 34913 56960
rect 34913 56926 34922 56960
rect 34870 56917 34922 56926
rect 36502 56917 36554 56969
rect 38038 56960 38090 56969
rect 38038 56926 38047 56960
rect 38047 56926 38081 56960
rect 38081 56926 38090 56960
rect 38038 56917 38090 56926
rect 41206 56917 41258 56969
rect 42838 56917 42890 56969
rect 44374 56917 44426 56969
rect 47542 56960 47594 56969
rect 47542 56926 47551 56960
rect 47551 56926 47585 56960
rect 47585 56926 47594 56960
rect 49078 56960 49130 56969
rect 47542 56917 47594 56926
rect 49078 56926 49087 56960
rect 49087 56926 49121 56960
rect 49121 56926 49130 56960
rect 49078 56917 49130 56926
rect 50710 56917 50762 56969
rect 53878 56960 53930 56969
rect 53878 56926 53887 56960
rect 53887 56926 53921 56960
rect 53921 56926 53930 56960
rect 53878 56917 53930 56926
rect 55414 56960 55466 56969
rect 55414 56926 55423 56960
rect 55423 56926 55457 56960
rect 55457 56926 55466 56960
rect 55414 56917 55466 56926
rect 7894 56843 7946 56895
rect 6070 56769 6122 56821
rect 9046 56769 9098 56821
rect 20854 56886 20906 56895
rect 20854 56852 20863 56886
rect 20863 56852 20897 56886
rect 20897 56852 20906 56886
rect 20854 56843 20906 56852
rect 21622 56843 21674 56895
rect 32566 56843 32618 56895
rect 34102 56886 34154 56895
rect 34102 56852 34111 56886
rect 34111 56852 34145 56886
rect 34145 56852 34154 56886
rect 34102 56843 34154 56852
rect 39670 56843 39722 56895
rect 40822 56886 40874 56895
rect 40822 56852 40831 56886
rect 40831 56852 40865 56886
rect 40865 56852 40874 56886
rect 40822 56843 40874 56852
rect 43030 56886 43082 56895
rect 43030 56852 43039 56886
rect 43039 56852 43073 56886
rect 43073 56852 43082 56886
rect 43030 56843 43082 56852
rect 45910 56843 45962 56895
rect 48886 56886 48938 56895
rect 48886 56852 48895 56886
rect 48895 56852 48929 56886
rect 48929 56852 48938 56886
rect 48886 56843 48938 56852
rect 50902 56886 50954 56895
rect 50902 56852 50911 56886
rect 50911 56852 50945 56886
rect 50945 56852 50954 56886
rect 50902 56843 50954 56852
rect 52246 56843 52298 56895
rect 32470 56769 32522 56821
rect 39862 56769 39914 56821
rect 42838 56769 42890 56821
rect 54838 56769 54890 56821
rect 4822 56695 4874 56747
rect 5206 56738 5258 56747
rect 5206 56704 5215 56738
rect 5215 56704 5249 56738
rect 5249 56704 5258 56738
rect 5206 56695 5258 56704
rect 5782 56738 5834 56747
rect 5782 56704 5791 56738
rect 5791 56704 5825 56738
rect 5825 56704 5834 56738
rect 5782 56695 5834 56704
rect 7318 56738 7370 56747
rect 7318 56704 7327 56738
rect 7327 56704 7361 56738
rect 7361 56704 7370 56738
rect 7318 56695 7370 56704
rect 10006 56738 10058 56747
rect 10006 56704 10015 56738
rect 10015 56704 10049 56738
rect 10049 56704 10058 56738
rect 10006 56695 10058 56704
rect 13078 56738 13130 56747
rect 13078 56704 13087 56738
rect 13087 56704 13121 56738
rect 13121 56704 13130 56738
rect 13078 56695 13130 56704
rect 13654 56738 13706 56747
rect 13654 56704 13663 56738
rect 13663 56704 13697 56738
rect 13697 56704 13706 56738
rect 13654 56695 13706 56704
rect 16054 56738 16106 56747
rect 16054 56704 16063 56738
rect 16063 56704 16097 56738
rect 16097 56704 16106 56738
rect 16054 56695 16106 56704
rect 17878 56738 17930 56747
rect 17878 56704 17887 56738
rect 17887 56704 17921 56738
rect 17921 56704 17930 56738
rect 17878 56695 17930 56704
rect 19222 56738 19274 56747
rect 19222 56704 19231 56738
rect 19231 56704 19265 56738
rect 19265 56704 19274 56738
rect 19222 56695 19274 56704
rect 21814 56695 21866 56747
rect 22006 56695 22058 56747
rect 27286 56738 27338 56747
rect 27286 56704 27295 56738
rect 27295 56704 27329 56738
rect 27329 56704 27338 56738
rect 27286 56695 27338 56704
rect 36118 56695 36170 56747
rect 36886 56738 36938 56747
rect 36886 56704 36895 56738
rect 36895 56704 36929 56738
rect 36929 56704 36938 56738
rect 36886 56695 36938 56704
rect 39670 56695 39722 56747
rect 40342 56695 40394 56747
rect 46102 56695 46154 56747
rect 52822 56738 52874 56747
rect 52822 56704 52831 56738
rect 52831 56704 52865 56738
rect 52865 56704 52874 56738
rect 52822 56695 52874 56704
rect 55702 56738 55754 56747
rect 55702 56704 55711 56738
rect 55711 56704 55745 56738
rect 55745 56704 55754 56738
rect 55702 56695 55754 56704
rect 56950 56738 57002 56747
rect 56950 56704 56959 56738
rect 56959 56704 56993 56738
rect 56993 56704 57002 56738
rect 56950 56695 57002 56704
rect 19654 56584 19706 56636
rect 19718 56584 19770 56636
rect 19782 56584 19834 56636
rect 19846 56584 19898 56636
rect 50374 56584 50426 56636
rect 50438 56584 50490 56636
rect 50502 56584 50554 56636
rect 50566 56584 50618 56636
rect 694 56473 746 56525
rect 2806 56473 2858 56525
rect 3862 56473 3914 56525
rect 5398 56473 5450 56525
rect 5974 56473 6026 56525
rect 7030 56473 7082 56525
rect 8566 56473 8618 56525
rect 10198 56473 10250 56525
rect 10678 56473 10730 56525
rect 11734 56473 11786 56525
rect 12310 56473 12362 56525
rect 13366 56473 13418 56525
rect 14902 56473 14954 56525
rect 15382 56473 15434 56525
rect 17014 56473 17066 56525
rect 18550 56473 18602 56525
rect 19990 56473 20042 56525
rect 21238 56473 21290 56525
rect 21718 56473 21770 56525
rect 22774 56473 22826 56525
rect 24406 56473 24458 56525
rect 25942 56473 25994 56525
rect 26518 56473 26570 56525
rect 27574 56473 27626 56525
rect 28054 56473 28106 56525
rect 29686 56516 29738 56525
rect 29686 56482 29695 56516
rect 29695 56482 29729 56516
rect 29729 56482 29738 56516
rect 29686 56473 29738 56482
rect 30646 56473 30698 56525
rect 31222 56473 31274 56525
rect 32278 56473 32330 56525
rect 32758 56473 32810 56525
rect 33814 56473 33866 56525
rect 34582 56473 34634 56525
rect 35446 56473 35498 56525
rect 27286 56399 27338 56451
rect 32470 56399 32522 56451
rect 36022 56399 36074 56451
rect 37558 56473 37610 56525
rect 38614 56473 38666 56525
rect 40150 56516 40202 56525
rect 40150 56482 40159 56516
rect 40159 56482 40193 56516
rect 40193 56482 40202 56516
rect 40150 56473 40202 56482
rect 41782 56473 41834 56525
rect 43318 56473 43370 56525
rect 43894 56473 43946 56525
rect 44950 56473 45002 56525
rect 46486 56473 46538 56525
rect 48022 56473 48074 56525
rect 48598 56473 48650 56525
rect 49654 56473 49706 56525
rect 50134 56473 50186 56525
rect 52918 56516 52970 56525
rect 52918 56482 52927 56516
rect 52927 56482 52961 56516
rect 52961 56482 52970 56516
rect 52918 56473 52970 56482
rect 53302 56473 53354 56525
rect 54358 56473 54410 56525
rect 54934 56473 54986 56525
rect 55990 56516 56042 56525
rect 55990 56482 55999 56516
rect 55999 56482 56033 56516
rect 56033 56482 56042 56516
rect 55990 56473 56042 56482
rect 38902 56399 38954 56451
rect 46198 56399 46250 56451
rect 48310 56325 48362 56377
rect 54838 56325 54890 56377
rect 22870 56251 22922 56303
rect 41782 56251 41834 56303
rect 46294 56251 46346 56303
rect 50038 56251 50090 56303
rect 1750 56220 1802 56229
rect 1750 56186 1759 56220
rect 1759 56186 1793 56220
rect 1793 56186 1802 56220
rect 1750 56177 1802 56186
rect 2998 56220 3050 56229
rect 2998 56186 3007 56220
rect 3007 56186 3041 56220
rect 3041 56186 3050 56220
rect 2998 56177 3050 56186
rect 4726 56177 4778 56229
rect 5590 56220 5642 56229
rect 5590 56186 5599 56220
rect 5599 56186 5633 56220
rect 5633 56186 5642 56220
rect 5590 56177 5642 56186
rect 6358 56220 6410 56229
rect 6358 56186 6367 56220
rect 6367 56186 6401 56220
rect 6401 56186 6410 56220
rect 6358 56177 6410 56186
rect 7222 56220 7274 56229
rect 7222 56186 7231 56220
rect 7231 56186 7265 56220
rect 7265 56186 7274 56220
rect 7222 56177 7274 56186
rect 8566 56220 8618 56229
rect 8566 56186 8575 56220
rect 8575 56186 8609 56220
rect 8609 56186 8618 56220
rect 10102 56220 10154 56229
rect 8566 56177 8618 56186
rect 10102 56186 10111 56220
rect 10111 56186 10145 56220
rect 10145 56186 10154 56220
rect 10102 56177 10154 56186
rect 11158 56220 11210 56229
rect 11158 56186 11167 56220
rect 11167 56186 11201 56220
rect 11201 56186 11210 56220
rect 11158 56177 11210 56186
rect 11926 56220 11978 56229
rect 11926 56186 11935 56220
rect 11935 56186 11969 56220
rect 11969 56186 11978 56220
rect 11926 56177 11978 56186
rect 12310 56220 12362 56229
rect 12310 56186 12319 56220
rect 12319 56186 12353 56220
rect 12353 56186 12362 56220
rect 12310 56177 12362 56186
rect 13558 56220 13610 56229
rect 13558 56186 13567 56220
rect 13567 56186 13601 56220
rect 13601 56186 13610 56220
rect 13558 56177 13610 56186
rect 15190 56177 15242 56229
rect 15286 56177 15338 56229
rect 16822 56220 16874 56229
rect 16822 56186 16831 56220
rect 16831 56186 16865 56220
rect 16865 56186 16874 56220
rect 16822 56177 16874 56186
rect 18070 56177 18122 56229
rect 20374 56220 20426 56229
rect 20374 56186 20383 56220
rect 20383 56186 20417 56220
rect 20417 56186 20426 56220
rect 20374 56177 20426 56186
rect 21430 56220 21482 56229
rect 21430 56186 21439 56220
rect 21439 56186 21473 56220
rect 21473 56186 21482 56220
rect 21430 56177 21482 56186
rect 22102 56220 22154 56229
rect 22102 56186 22111 56220
rect 22111 56186 22145 56220
rect 22145 56186 22154 56220
rect 22102 56177 22154 56186
rect 22678 56177 22730 56229
rect 24406 56220 24458 56229
rect 24406 56186 24415 56220
rect 24415 56186 24449 56220
rect 24449 56186 24458 56220
rect 24406 56177 24458 56186
rect 26134 56220 26186 56229
rect 26134 56186 26143 56220
rect 26143 56186 26177 56220
rect 26177 56186 26186 56220
rect 26134 56177 26186 56186
rect 27766 56220 27818 56229
rect 27766 56186 27775 56220
rect 27775 56186 27809 56220
rect 27809 56186 27818 56220
rect 27766 56177 27818 56186
rect 28438 56220 28490 56229
rect 28438 56186 28447 56220
rect 28447 56186 28481 56220
rect 28481 56186 28490 56220
rect 28438 56177 28490 56186
rect 29590 56220 29642 56229
rect 29590 56186 29599 56220
rect 29599 56186 29633 56220
rect 29633 56186 29642 56220
rect 29590 56177 29642 56186
rect 30934 56220 30986 56229
rect 30934 56186 30943 56220
rect 30943 56186 30977 56220
rect 30977 56186 30986 56220
rect 30934 56177 30986 56186
rect 32470 56220 32522 56229
rect 32470 56186 32479 56220
rect 32479 56186 32513 56220
rect 32513 56186 32522 56220
rect 32470 56177 32522 56186
rect 34198 56177 34250 56229
rect 34390 56220 34442 56229
rect 34390 56186 34399 56220
rect 34399 56186 34433 56220
rect 34433 56186 34442 56220
rect 34390 56177 34442 56186
rect 36214 56220 36266 56229
rect 36214 56186 36223 56220
rect 36223 56186 36257 56220
rect 36257 56186 36266 56220
rect 36598 56220 36650 56229
rect 36214 56177 36266 56186
rect 36598 56186 36607 56220
rect 36607 56186 36641 56220
rect 36641 56186 36650 56220
rect 36598 56177 36650 56186
rect 37750 56220 37802 56229
rect 37750 56186 37759 56220
rect 37759 56186 37793 56220
rect 37793 56186 37802 56220
rect 37750 56177 37802 56186
rect 38710 56220 38762 56229
rect 38710 56186 38719 56220
rect 38719 56186 38753 56220
rect 38753 56186 38762 56220
rect 38710 56177 38762 56186
rect 38806 56177 38858 56229
rect 41590 56220 41642 56229
rect 41590 56186 41599 56220
rect 41599 56186 41633 56220
rect 41633 56186 41642 56220
rect 41590 56177 41642 56186
rect 43414 56220 43466 56229
rect 2230 56103 2282 56155
rect 5782 56103 5834 56155
rect 18166 56103 18218 56155
rect 21814 56103 21866 56155
rect 37078 56103 37130 56155
rect 40342 56103 40394 56155
rect 40726 56103 40778 56155
rect 43414 56186 43423 56220
rect 43423 56186 43457 56220
rect 43457 56186 43466 56220
rect 43414 56177 43466 56186
rect 43894 56220 43946 56229
rect 43894 56186 43903 56220
rect 43903 56186 43937 56220
rect 43937 56186 43946 56220
rect 43894 56177 43946 56186
rect 44758 56220 44810 56229
rect 44758 56186 44767 56220
rect 44767 56186 44801 56220
rect 44801 56186 44810 56220
rect 44758 56177 44810 56186
rect 46774 56220 46826 56229
rect 46774 56186 46783 56220
rect 46783 56186 46817 56220
rect 46817 56186 46826 56220
rect 46774 56177 46826 56186
rect 47830 56220 47882 56229
rect 47830 56186 47839 56220
rect 47839 56186 47873 56220
rect 47873 56186 47882 56220
rect 47830 56177 47882 56186
rect 48598 56220 48650 56229
rect 48598 56186 48607 56220
rect 48607 56186 48641 56220
rect 48641 56186 48650 56220
rect 48598 56177 48650 56186
rect 50230 56220 50282 56229
rect 50230 56186 50239 56220
rect 50239 56186 50273 56220
rect 50273 56186 50282 56220
rect 50230 56177 50282 56186
rect 51670 56220 51722 56229
rect 51670 56186 51679 56220
rect 51679 56186 51713 56220
rect 51713 56186 51722 56220
rect 51670 56177 51722 56186
rect 53398 56220 53450 56229
rect 51190 56103 51242 56155
rect 53398 56186 53407 56220
rect 53407 56186 53441 56220
rect 53441 56186 53450 56220
rect 53398 56177 53450 56186
rect 58582 56251 58634 56303
rect 58198 56177 58250 56229
rect 4294 55918 4346 55970
rect 4358 55918 4410 55970
rect 4422 55918 4474 55970
rect 4486 55918 4538 55970
rect 35014 55918 35066 55970
rect 35078 55918 35130 55970
rect 35142 55918 35194 55970
rect 35206 55918 35258 55970
rect 36118 55807 36170 55859
rect 38902 55733 38954 55785
rect 1174 55659 1226 55711
rect 4630 55659 4682 55711
rect 7510 55659 7562 55711
rect 9142 55659 9194 55711
rect 13846 55659 13898 55711
rect 20182 55659 20234 55711
rect 23350 55659 23402 55711
rect 24886 55659 24938 55711
rect 41782 55807 41834 55859
rect 42262 55659 42314 55711
rect 45430 55659 45482 55711
rect 46966 55659 47018 55711
rect 51766 55659 51818 55711
rect 56470 55659 56522 55711
rect 57526 55659 57578 55711
rect 5398 55511 5450 55563
rect 7702 55554 7754 55563
rect 7702 55520 7711 55554
rect 7711 55520 7745 55554
rect 7745 55520 7754 55554
rect 7702 55511 7754 55520
rect 9334 55554 9386 55563
rect 9334 55520 9343 55554
rect 9343 55520 9377 55554
rect 9377 55520 9386 55554
rect 9334 55511 9386 55520
rect 12406 55554 12458 55563
rect 12406 55520 12415 55554
rect 12415 55520 12449 55554
rect 12449 55520 12458 55554
rect 12406 55511 12458 55520
rect 20470 55511 20522 55563
rect 25078 55554 25130 55563
rect 25078 55520 25087 55554
rect 25087 55520 25121 55554
rect 25121 55520 25130 55554
rect 25078 55511 25130 55520
rect 42550 55554 42602 55563
rect 42550 55520 42559 55554
rect 42559 55520 42593 55554
rect 42593 55520 42602 55554
rect 42550 55511 42602 55520
rect 45526 55554 45578 55563
rect 45526 55520 45535 55554
rect 45535 55520 45569 55554
rect 45569 55520 45578 55554
rect 45526 55511 45578 55520
rect 52054 55511 52106 55563
rect 2038 55406 2090 55415
rect 2038 55372 2047 55406
rect 2047 55372 2081 55406
rect 2081 55372 2090 55406
rect 2038 55363 2090 55372
rect 13846 55363 13898 55415
rect 23158 55406 23210 55415
rect 23158 55372 23167 55406
rect 23167 55372 23201 55406
rect 23201 55372 23210 55406
rect 23158 55363 23210 55372
rect 39766 55363 39818 55415
rect 46966 55363 47018 55415
rect 55606 55406 55658 55415
rect 55606 55372 55615 55406
rect 55615 55372 55649 55406
rect 55649 55372 55658 55406
rect 55894 55511 55946 55563
rect 57334 55406 57386 55415
rect 55606 55363 55658 55372
rect 57334 55372 57343 55406
rect 57343 55372 57377 55406
rect 57377 55372 57386 55406
rect 57334 55363 57386 55372
rect 19654 55252 19706 55304
rect 19718 55252 19770 55304
rect 19782 55252 19834 55304
rect 19846 55252 19898 55304
rect 50374 55252 50426 55304
rect 50438 55252 50490 55304
rect 50502 55252 50554 55304
rect 50566 55252 50618 55304
rect 12406 55141 12458 55193
rect 28342 55141 28394 55193
rect 39094 55141 39146 55193
rect 59158 55141 59210 55193
rect 2038 54993 2090 55045
rect 55606 54993 55658 55045
rect 39286 54888 39338 54897
rect 39286 54854 39295 54888
rect 39295 54854 39329 54888
rect 39329 54854 39338 54888
rect 39286 54845 39338 54854
rect 57910 54888 57962 54897
rect 57910 54854 57919 54888
rect 57919 54854 57953 54888
rect 57953 54854 57962 54888
rect 57910 54845 57962 54854
rect 53974 54771 54026 54823
rect 35830 54740 35882 54749
rect 35830 54706 35839 54740
rect 35839 54706 35873 54740
rect 35873 54706 35882 54740
rect 35830 54697 35882 54706
rect 39862 54740 39914 54749
rect 39862 54706 39871 54740
rect 39871 54706 39905 54740
rect 39905 54706 39914 54740
rect 39862 54697 39914 54706
rect 53878 54740 53930 54749
rect 53878 54706 53887 54740
rect 53887 54706 53921 54740
rect 53921 54706 53930 54740
rect 53878 54697 53930 54706
rect 4294 54586 4346 54638
rect 4358 54586 4410 54638
rect 4422 54586 4474 54638
rect 4486 54586 4538 54638
rect 35014 54586 35066 54638
rect 35078 54586 35130 54638
rect 35142 54586 35194 54638
rect 35206 54586 35258 54638
rect 11158 54475 11210 54527
rect 58102 54327 58154 54379
rect 31222 54179 31274 54231
rect 31126 54031 31178 54083
rect 57814 54179 57866 54231
rect 34870 54031 34922 54083
rect 36310 54074 36362 54083
rect 36310 54040 36319 54074
rect 36319 54040 36353 54074
rect 36353 54040 36362 54074
rect 36310 54031 36362 54040
rect 19654 53920 19706 53972
rect 19718 53920 19770 53972
rect 19782 53920 19834 53972
rect 19846 53920 19898 53972
rect 50374 53920 50426 53972
rect 50438 53920 50490 53972
rect 50502 53920 50554 53972
rect 50566 53920 50618 53972
rect 59638 53809 59690 53861
rect 25558 53513 25610 53565
rect 26614 53365 26666 53417
rect 49654 53365 49706 53417
rect 4294 53254 4346 53306
rect 4358 53254 4410 53306
rect 4422 53254 4474 53306
rect 4486 53254 4538 53306
rect 35014 53254 35066 53306
rect 35078 53254 35130 53306
rect 35142 53254 35194 53306
rect 35206 53254 35258 53306
rect 17014 52773 17066 52825
rect 16342 52699 16394 52751
rect 19654 52588 19706 52640
rect 19718 52588 19770 52640
rect 19782 52588 19834 52640
rect 19846 52588 19898 52640
rect 50374 52588 50426 52640
rect 50438 52588 50490 52640
rect 50502 52588 50554 52640
rect 50566 52588 50618 52640
rect 2134 52033 2186 52085
rect 22198 52033 22250 52085
rect 32662 52076 32714 52085
rect 32662 52042 32671 52076
rect 32671 52042 32705 52076
rect 32705 52042 32714 52076
rect 32662 52033 32714 52042
rect 4294 51922 4346 51974
rect 4358 51922 4410 51974
rect 4422 51922 4474 51974
rect 4486 51922 4538 51974
rect 35014 51922 35066 51974
rect 35078 51922 35130 51974
rect 35142 51922 35194 51974
rect 35206 51922 35258 51974
rect 30934 51589 30986 51641
rect 23254 51558 23306 51567
rect 23254 51524 23263 51558
rect 23263 51524 23297 51558
rect 23297 51524 23306 51558
rect 23254 51515 23306 51524
rect 53398 51515 53450 51567
rect 53206 51367 53258 51419
rect 19654 51256 19706 51308
rect 19718 51256 19770 51308
rect 19782 51256 19834 51308
rect 19846 51256 19898 51308
rect 50374 51256 50426 51308
rect 50438 51256 50490 51308
rect 50502 51256 50554 51308
rect 50566 51256 50618 51308
rect 21430 51145 21482 51197
rect 11062 50775 11114 50827
rect 14998 50775 15050 50827
rect 14038 50701 14090 50753
rect 55030 50701 55082 50753
rect 4294 50590 4346 50642
rect 4358 50590 4410 50642
rect 4422 50590 4474 50642
rect 4486 50590 4538 50642
rect 35014 50590 35066 50642
rect 35078 50590 35130 50642
rect 35142 50590 35194 50642
rect 35206 50590 35258 50642
rect 47254 50405 47306 50457
rect 25846 50257 25898 50309
rect 55702 50257 55754 50309
rect 52438 50183 52490 50235
rect 5590 50109 5642 50161
rect 27766 50109 27818 50161
rect 38806 50109 38858 50161
rect 46198 50035 46250 50087
rect 47254 50035 47306 50087
rect 54454 50035 54506 50087
rect 19654 49924 19706 49976
rect 19718 49924 19770 49976
rect 19782 49924 19834 49976
rect 19846 49924 19898 49976
rect 50374 49924 50426 49976
rect 50438 49924 50490 49976
rect 50502 49924 50554 49976
rect 50566 49924 50618 49976
rect 25558 49813 25610 49865
rect 25846 49739 25898 49791
rect 56950 49665 57002 49717
rect 46774 49517 46826 49569
rect 22966 49443 23018 49495
rect 12214 49412 12266 49421
rect 12214 49378 12223 49412
rect 12223 49378 12257 49412
rect 12257 49378 12266 49412
rect 12214 49369 12266 49378
rect 23062 49412 23114 49421
rect 23062 49378 23071 49412
rect 23071 49378 23105 49412
rect 23105 49378 23114 49412
rect 23062 49369 23114 49378
rect 4294 49258 4346 49310
rect 4358 49258 4410 49310
rect 4422 49258 4474 49310
rect 4486 49258 4538 49310
rect 35014 49258 35066 49310
rect 35078 49258 35130 49310
rect 35142 49258 35194 49310
rect 35206 49258 35258 49310
rect 26134 49147 26186 49199
rect 55894 49147 55946 49199
rect 56278 48925 56330 48977
rect 6934 48703 6986 48755
rect 46294 48703 46346 48755
rect 19654 48592 19706 48644
rect 19718 48592 19770 48644
rect 19782 48592 19834 48644
rect 19846 48592 19898 48644
rect 50374 48592 50426 48644
rect 50438 48592 50490 48644
rect 50502 48592 50554 48644
rect 50566 48592 50618 48644
rect 5398 48481 5450 48533
rect 22870 48481 22922 48533
rect 4822 48407 4874 48459
rect 6070 48407 6122 48459
rect 21958 48407 22010 48459
rect 4294 47926 4346 47978
rect 4358 47926 4410 47978
rect 4422 47926 4474 47978
rect 4486 47926 4538 47978
rect 35014 47926 35066 47978
rect 35078 47926 35130 47978
rect 35142 47926 35194 47978
rect 35206 47926 35258 47978
rect 27958 47519 28010 47571
rect 19654 47260 19706 47312
rect 19718 47260 19770 47312
rect 19782 47260 19834 47312
rect 19846 47260 19898 47312
rect 50374 47260 50426 47312
rect 50438 47260 50490 47312
rect 50502 47260 50554 47312
rect 50566 47260 50618 47312
rect 51574 46705 51626 46757
rect 4294 46594 4346 46646
rect 4358 46594 4410 46646
rect 4422 46594 4474 46646
rect 4486 46594 4538 46646
rect 35014 46594 35066 46646
rect 35078 46594 35130 46646
rect 35142 46594 35194 46646
rect 35206 46594 35258 46646
rect 29014 46335 29066 46387
rect 35830 46335 35882 46387
rect 20470 46261 20522 46313
rect 12790 46113 12842 46165
rect 13750 46156 13802 46165
rect 13750 46122 13759 46156
rect 13759 46122 13793 46156
rect 13793 46122 13802 46156
rect 13750 46113 13802 46122
rect 30838 46187 30890 46239
rect 41014 46113 41066 46165
rect 24406 46039 24458 46091
rect 50038 46082 50090 46091
rect 50038 46048 50047 46082
rect 50047 46048 50081 46082
rect 50081 46048 50090 46082
rect 50038 46039 50090 46048
rect 19654 45928 19706 45980
rect 19718 45928 19770 45980
rect 19782 45928 19834 45980
rect 19846 45928 19898 45980
rect 50374 45928 50426 45980
rect 50438 45928 50490 45980
rect 50502 45928 50554 45980
rect 50566 45928 50618 45980
rect 48310 45669 48362 45721
rect 28246 45416 28298 45425
rect 28246 45382 28255 45416
rect 28255 45382 28289 45416
rect 28289 45382 28298 45416
rect 28246 45373 28298 45382
rect 38902 45416 38954 45425
rect 38902 45382 38911 45416
rect 38911 45382 38945 45416
rect 38945 45382 38954 45416
rect 38902 45373 38954 45382
rect 4294 45262 4346 45314
rect 4358 45262 4410 45314
rect 4422 45262 4474 45314
rect 4486 45262 4538 45314
rect 35014 45262 35066 45314
rect 35078 45262 35130 45314
rect 35142 45262 35194 45314
rect 35206 45262 35258 45314
rect 30166 45151 30218 45203
rect 38902 45151 38954 45203
rect 28246 45077 28298 45129
rect 48982 45077 49034 45129
rect 44470 44707 44522 44759
rect 19654 44596 19706 44648
rect 19718 44596 19770 44648
rect 19782 44596 19834 44648
rect 19846 44596 19898 44648
rect 50374 44596 50426 44648
rect 50438 44596 50490 44648
rect 50502 44596 50554 44648
rect 50566 44596 50618 44648
rect 6358 44041 6410 44093
rect 30742 44041 30794 44093
rect 32758 44084 32810 44093
rect 32758 44050 32767 44084
rect 32767 44050 32801 44084
rect 32801 44050 32810 44084
rect 32758 44041 32810 44050
rect 33142 44084 33194 44093
rect 33142 44050 33151 44084
rect 33151 44050 33185 44084
rect 33185 44050 33194 44084
rect 33142 44041 33194 44050
rect 34774 44084 34826 44093
rect 34774 44050 34783 44084
rect 34783 44050 34817 44084
rect 34817 44050 34826 44084
rect 34774 44041 34826 44050
rect 55318 44084 55370 44093
rect 55318 44050 55327 44084
rect 55327 44050 55361 44084
rect 55361 44050 55370 44084
rect 55318 44041 55370 44050
rect 4294 43930 4346 43982
rect 4358 43930 4410 43982
rect 4422 43930 4474 43982
rect 4486 43930 4538 43982
rect 35014 43930 35066 43982
rect 35078 43930 35130 43982
rect 35142 43930 35194 43982
rect 35206 43930 35258 43982
rect 30742 43819 30794 43871
rect 55894 43819 55946 43871
rect 7606 43745 7658 43797
rect 33142 43745 33194 43797
rect 32758 43671 32810 43723
rect 49750 43671 49802 43723
rect 26710 43375 26762 43427
rect 57142 43523 57194 43575
rect 19654 43264 19706 43316
rect 19718 43264 19770 43316
rect 19782 43264 19834 43316
rect 19846 43264 19898 43316
rect 50374 43264 50426 43316
rect 50438 43264 50490 43316
rect 50502 43264 50554 43316
rect 50566 43264 50618 43316
rect 57814 43005 57866 43057
rect 38134 42783 38186 42835
rect 34678 42752 34730 42761
rect 34678 42718 34687 42752
rect 34687 42718 34721 42752
rect 34721 42718 34730 42752
rect 34678 42709 34730 42718
rect 52534 42752 52586 42761
rect 52534 42718 52543 42752
rect 52543 42718 52577 42752
rect 52577 42718 52586 42752
rect 52534 42709 52586 42718
rect 4294 42598 4346 42650
rect 4358 42598 4410 42650
rect 4422 42598 4474 42650
rect 4486 42598 4538 42650
rect 35014 42598 35066 42650
rect 35078 42598 35130 42650
rect 35142 42598 35194 42650
rect 35206 42598 35258 42650
rect 17974 42487 18026 42539
rect 34678 42487 34730 42539
rect 41110 42487 41162 42539
rect 52534 42487 52586 42539
rect 30070 42191 30122 42243
rect 43702 42191 43754 42243
rect 30070 42086 30122 42095
rect 30070 42052 30079 42086
rect 30079 42052 30113 42086
rect 30113 42052 30122 42086
rect 30070 42043 30122 42052
rect 40822 42043 40874 42095
rect 19654 41932 19706 41984
rect 19718 41932 19770 41984
rect 19782 41932 19834 41984
rect 19846 41932 19898 41984
rect 50374 41932 50426 41984
rect 50438 41932 50490 41984
rect 50502 41932 50554 41984
rect 50566 41932 50618 41984
rect 7318 41525 7370 41577
rect 9334 41451 9386 41503
rect 5206 41377 5258 41429
rect 42070 41377 42122 41429
rect 57238 41420 57290 41429
rect 57238 41386 57247 41420
rect 57247 41386 57281 41420
rect 57281 41386 57290 41420
rect 57238 41377 57290 41386
rect 4294 41266 4346 41318
rect 4358 41266 4410 41318
rect 4422 41266 4474 41318
rect 4486 41266 4538 41318
rect 35014 41266 35066 41318
rect 35078 41266 35130 41318
rect 35142 41266 35194 41318
rect 35206 41266 35258 41318
rect 8566 40933 8618 40985
rect 26806 40859 26858 40911
rect 41206 40711 41258 40763
rect 19654 40600 19706 40652
rect 19718 40600 19770 40652
rect 19782 40600 19834 40652
rect 19846 40600 19898 40652
rect 50374 40600 50426 40652
rect 50438 40600 50490 40652
rect 50502 40600 50554 40652
rect 50566 40600 50618 40652
rect 7222 40341 7274 40393
rect 18070 40267 18122 40319
rect 52054 40310 52106 40319
rect 52054 40276 52063 40310
rect 52063 40276 52097 40310
rect 52097 40276 52106 40310
rect 52054 40267 52106 40276
rect 4294 39934 4346 39986
rect 4358 39934 4410 39986
rect 4422 39934 4474 39986
rect 4486 39934 4538 39986
rect 35014 39934 35066 39986
rect 35078 39934 35130 39986
rect 35142 39934 35194 39986
rect 35206 39934 35258 39986
rect 25174 39527 25226 39579
rect 46678 39527 46730 39579
rect 25270 39453 25322 39505
rect 47542 39453 47594 39505
rect 45334 39379 45386 39431
rect 19654 39268 19706 39320
rect 19718 39268 19770 39320
rect 19782 39268 19834 39320
rect 19846 39268 19898 39320
rect 50374 39268 50426 39320
rect 50438 39268 50490 39320
rect 50502 39268 50554 39320
rect 50566 39268 50618 39320
rect 46822 39083 46874 39135
rect 47542 39157 47594 39209
rect 36214 38787 36266 38839
rect 21334 38756 21386 38765
rect 21334 38722 21343 38756
rect 21343 38722 21377 38756
rect 21377 38722 21386 38756
rect 21334 38713 21386 38722
rect 27190 38756 27242 38765
rect 27190 38722 27199 38756
rect 27199 38722 27233 38756
rect 27233 38722 27242 38756
rect 27190 38713 27242 38722
rect 41302 38713 41354 38765
rect 46870 38713 46922 38765
rect 4294 38602 4346 38654
rect 4358 38602 4410 38654
rect 4422 38602 4474 38654
rect 4486 38602 4538 38654
rect 35014 38602 35066 38654
rect 35078 38602 35130 38654
rect 35142 38602 35194 38654
rect 35206 38602 35258 38654
rect 27190 38491 27242 38543
rect 39190 38491 39242 38543
rect 13558 38343 13610 38395
rect 24694 38195 24746 38247
rect 30262 38238 30314 38247
rect 30262 38204 30271 38238
rect 30271 38204 30305 38238
rect 30305 38204 30314 38238
rect 30262 38195 30314 38204
rect 32470 38269 32522 38321
rect 15190 38121 15242 38173
rect 32374 38121 32426 38173
rect 19654 37936 19706 37988
rect 19718 37936 19770 37988
rect 19782 37936 19834 37988
rect 19846 37936 19898 37988
rect 50374 37936 50426 37988
rect 50438 37936 50490 37988
rect 50502 37936 50554 37988
rect 50566 37936 50618 37988
rect 42934 37455 42986 37507
rect 16438 37424 16490 37433
rect 16438 37390 16447 37424
rect 16447 37390 16481 37424
rect 16481 37390 16490 37424
rect 16438 37381 16490 37390
rect 41782 37424 41834 37433
rect 41782 37390 41791 37424
rect 41791 37390 41825 37424
rect 41825 37390 41834 37424
rect 41782 37381 41834 37390
rect 53782 37381 53834 37433
rect 4294 37270 4346 37322
rect 4358 37270 4410 37322
rect 4422 37270 4474 37322
rect 4486 37270 4538 37322
rect 35014 37270 35066 37322
rect 35078 37270 35130 37322
rect 35142 37270 35194 37322
rect 35206 37270 35258 37322
rect 41782 37159 41834 37211
rect 53110 37159 53162 37211
rect 32758 37085 32810 37137
rect 53782 37085 53834 37137
rect 25366 36715 25418 36767
rect 42934 36715 42986 36767
rect 19654 36604 19706 36656
rect 19718 36604 19770 36656
rect 19782 36604 19834 36656
rect 19846 36604 19898 36656
rect 50374 36604 50426 36656
rect 50438 36604 50490 36656
rect 50502 36604 50554 36656
rect 50566 36604 50618 36656
rect 20374 36197 20426 36249
rect 1942 36092 1994 36101
rect 1942 36058 1951 36092
rect 1951 36058 1985 36092
rect 1985 36058 1994 36092
rect 1942 36049 1994 36058
rect 7990 36049 8042 36101
rect 38518 36092 38570 36101
rect 38518 36058 38527 36092
rect 38527 36058 38561 36092
rect 38561 36058 38570 36092
rect 38518 36049 38570 36058
rect 54742 36092 54794 36101
rect 54742 36058 54751 36092
rect 54751 36058 54785 36092
rect 54785 36058 54794 36092
rect 54742 36049 54794 36058
rect 4294 35938 4346 35990
rect 4358 35938 4410 35990
rect 4422 35938 4474 35990
rect 4486 35938 4538 35990
rect 35014 35938 35066 35990
rect 35078 35938 35130 35990
rect 35142 35938 35194 35990
rect 35206 35938 35258 35990
rect 4534 35605 4586 35657
rect 22678 35679 22730 35731
rect 20470 35574 20522 35583
rect 20470 35540 20479 35574
rect 20479 35540 20513 35574
rect 20513 35540 20522 35574
rect 20470 35531 20522 35540
rect 39958 35531 40010 35583
rect 35926 35457 35978 35509
rect 32566 35383 32618 35435
rect 44374 35383 44426 35435
rect 47926 35383 47978 35435
rect 51190 35426 51242 35435
rect 51190 35392 51199 35426
rect 51199 35392 51233 35426
rect 51233 35392 51242 35426
rect 51190 35383 51242 35392
rect 19654 35272 19706 35324
rect 19718 35272 19770 35324
rect 19782 35272 19834 35324
rect 19846 35272 19898 35324
rect 50374 35272 50426 35324
rect 50438 35272 50490 35324
rect 50502 35272 50554 35324
rect 50566 35272 50618 35324
rect 29398 35161 29450 35213
rect 51190 35161 51242 35213
rect 21622 35087 21674 35139
rect 4534 35056 4586 35065
rect 4534 35022 4543 35056
rect 4543 35022 4577 35056
rect 4577 35022 4586 35056
rect 4534 35013 4586 35022
rect 19126 34865 19178 34917
rect 19990 34791 20042 34843
rect 17782 34760 17834 34769
rect 17782 34726 17791 34760
rect 17791 34726 17825 34760
rect 17825 34726 17834 34760
rect 17782 34717 17834 34726
rect 20374 34717 20426 34769
rect 4294 34606 4346 34658
rect 4358 34606 4410 34658
rect 4422 34606 4474 34658
rect 4486 34606 4538 34658
rect 35014 34606 35066 34658
rect 35078 34606 35130 34658
rect 35142 34606 35194 34658
rect 35206 34606 35258 34658
rect 33814 34199 33866 34251
rect 36694 34242 36746 34251
rect 36694 34208 36703 34242
rect 36703 34208 36737 34242
rect 36737 34208 36746 34242
rect 36694 34199 36746 34208
rect 17782 34051 17834 34103
rect 32470 34051 32522 34103
rect 19654 33940 19706 33992
rect 19718 33940 19770 33992
rect 19782 33940 19834 33992
rect 19846 33940 19898 33992
rect 50374 33940 50426 33992
rect 50438 33940 50490 33992
rect 50502 33940 50554 33992
rect 50566 33940 50618 33992
rect 9334 33829 9386 33881
rect 57238 33829 57290 33881
rect 41398 33459 41450 33511
rect 45718 33385 45770 33437
rect 4294 33274 4346 33326
rect 4358 33274 4410 33326
rect 4422 33274 4474 33326
rect 4486 33274 4538 33326
rect 35014 33274 35066 33326
rect 35078 33274 35130 33326
rect 35142 33274 35194 33326
rect 35206 33274 35258 33326
rect 57910 33163 57962 33215
rect 10006 33089 10058 33141
rect 8998 33015 9050 33067
rect 13078 33015 13130 33067
rect 8854 32719 8906 32771
rect 19654 32608 19706 32660
rect 19718 32608 19770 32660
rect 19782 32608 19834 32660
rect 19846 32608 19898 32660
rect 50374 32608 50426 32660
rect 50438 32608 50490 32660
rect 50502 32608 50554 32660
rect 50566 32608 50618 32660
rect 6838 32497 6890 32549
rect 8854 32497 8906 32549
rect 15286 32497 15338 32549
rect 6550 32349 6602 32401
rect 50902 32201 50954 32253
rect 42838 32127 42890 32179
rect 13078 32096 13130 32105
rect 13078 32062 13087 32096
rect 13087 32062 13121 32096
rect 13121 32062 13130 32096
rect 13078 32053 13130 32062
rect 4294 31942 4346 31994
rect 4358 31942 4410 31994
rect 4422 31942 4474 31994
rect 4486 31942 4538 31994
rect 35014 31942 35066 31994
rect 35078 31942 35130 31994
rect 35142 31942 35194 31994
rect 35206 31942 35258 31994
rect 6550 31831 6602 31883
rect 52822 31831 52874 31883
rect 6838 31757 6890 31809
rect 48886 31757 48938 31809
rect 26518 31726 26570 31735
rect 26518 31692 26527 31726
rect 26527 31692 26561 31726
rect 26561 31692 26570 31726
rect 26518 31683 26570 31692
rect 57430 31683 57482 31735
rect 19654 31276 19706 31328
rect 19718 31276 19770 31328
rect 19782 31276 19834 31328
rect 19846 31276 19898 31328
rect 50374 31276 50426 31328
rect 50438 31276 50490 31328
rect 50502 31276 50554 31328
rect 50566 31276 50618 31328
rect 1750 30869 1802 30921
rect 18838 30795 18890 30847
rect 40918 30795 40970 30847
rect 4294 30610 4346 30662
rect 4358 30610 4410 30662
rect 4422 30610 4474 30662
rect 4486 30610 4538 30662
rect 35014 30610 35066 30662
rect 35078 30610 35130 30662
rect 35142 30610 35194 30662
rect 35206 30610 35258 30662
rect 38230 30499 38282 30551
rect 45190 30499 45242 30551
rect 39286 30425 39338 30477
rect 40918 30425 40970 30477
rect 2998 30351 3050 30403
rect 36886 30351 36938 30403
rect 38326 30277 38378 30329
rect 45190 30314 45242 30366
rect 51094 30277 51146 30329
rect 44614 30129 44666 30181
rect 44902 30129 44954 30181
rect 19654 29944 19706 29996
rect 19718 29944 19770 29996
rect 19782 29944 19834 29996
rect 19846 29944 19898 29996
rect 50374 29944 50426 29996
rect 50438 29944 50490 29996
rect 50502 29944 50554 29996
rect 50566 29944 50618 29996
rect 44374 29833 44426 29885
rect 44566 29833 44618 29885
rect 3574 29463 3626 29515
rect 54742 29463 54794 29515
rect 41590 29389 41642 29441
rect 4294 29278 4346 29330
rect 4358 29278 4410 29330
rect 4422 29278 4474 29330
rect 4486 29278 4538 29330
rect 35014 29278 35066 29330
rect 35078 29278 35130 29330
rect 35142 29278 35194 29330
rect 35206 29278 35258 29330
rect 25462 28871 25514 28923
rect 52342 28797 52394 28849
rect 19654 28612 19706 28664
rect 19718 28612 19770 28664
rect 19782 28612 19834 28664
rect 19846 28612 19898 28664
rect 50374 28612 50426 28664
rect 50438 28612 50490 28664
rect 50502 28612 50554 28664
rect 50566 28612 50618 28664
rect 37750 28501 37802 28553
rect 3670 28279 3722 28331
rect 53878 28279 53930 28331
rect 13654 28205 13706 28257
rect 6262 28100 6314 28109
rect 6262 28066 6271 28100
rect 6271 28066 6305 28100
rect 6305 28066 6314 28100
rect 6262 28057 6314 28066
rect 15190 28057 15242 28109
rect 26806 28057 26858 28109
rect 55990 28057 56042 28109
rect 58006 28100 58058 28109
rect 58006 28066 58015 28100
rect 58015 28066 58049 28100
rect 58049 28066 58058 28100
rect 58006 28057 58058 28066
rect 4294 27946 4346 27998
rect 4358 27946 4410 27998
rect 4422 27946 4474 27998
rect 4486 27946 4538 27998
rect 35014 27946 35066 27998
rect 35078 27946 35130 27998
rect 35142 27946 35194 27998
rect 35206 27946 35258 27998
rect 27190 27835 27242 27887
rect 58006 27835 58058 27887
rect 19654 27280 19706 27332
rect 19718 27280 19770 27332
rect 19782 27280 19834 27332
rect 19846 27280 19898 27332
rect 50374 27280 50426 27332
rect 50438 27280 50490 27332
rect 50502 27280 50554 27332
rect 50566 27280 50618 27332
rect 43894 27021 43946 27073
rect 26518 26873 26570 26925
rect 46390 26873 46442 26925
rect 6550 26799 6602 26851
rect 32758 26799 32810 26851
rect 48214 26799 48266 26851
rect 4294 26614 4346 26666
rect 4358 26614 4410 26666
rect 4422 26614 4474 26666
rect 4486 26614 4538 26666
rect 35014 26614 35066 26666
rect 35078 26614 35130 26666
rect 35142 26614 35194 26666
rect 35206 26614 35258 26666
rect 40150 26250 40202 26259
rect 40150 26216 40159 26250
rect 40159 26216 40193 26250
rect 40193 26216 40202 26250
rect 40150 26207 40202 26216
rect 47734 26250 47786 26259
rect 47734 26216 47743 26250
rect 47743 26216 47777 26250
rect 47777 26216 47786 26250
rect 47734 26207 47786 26216
rect 54262 26207 54314 26259
rect 19654 25948 19706 26000
rect 19718 25948 19770 26000
rect 19782 25948 19834 26000
rect 19846 25948 19898 26000
rect 50374 25948 50426 26000
rect 50438 25948 50490 26000
rect 50502 25948 50554 26000
rect 50566 25948 50618 26000
rect 13846 25732 13898 25741
rect 13846 25698 13855 25732
rect 13855 25698 13889 25732
rect 13889 25698 13898 25732
rect 13846 25689 13898 25698
rect 10870 25541 10922 25593
rect 30070 25541 30122 25593
rect 22102 25467 22154 25519
rect 5398 25436 5450 25445
rect 5398 25402 5407 25436
rect 5407 25402 5441 25436
rect 5441 25402 5450 25436
rect 5398 25393 5450 25402
rect 36982 25393 37034 25445
rect 4294 25282 4346 25334
rect 4358 25282 4410 25334
rect 4422 25282 4474 25334
rect 4486 25282 4538 25334
rect 35014 25282 35066 25334
rect 35078 25282 35130 25334
rect 35142 25282 35194 25334
rect 35206 25282 35258 25334
rect 13558 25171 13610 25223
rect 36310 25171 36362 25223
rect 40150 25171 40202 25223
rect 51478 25171 51530 25223
rect 5398 25097 5450 25149
rect 45238 25097 45290 25149
rect 30646 24949 30698 25001
rect 31702 24875 31754 24927
rect 38710 24727 38762 24779
rect 19654 24616 19706 24668
rect 19718 24616 19770 24668
rect 19782 24616 19834 24668
rect 19846 24616 19898 24668
rect 50374 24616 50426 24668
rect 50438 24616 50490 24668
rect 50502 24616 50554 24668
rect 50566 24616 50618 24668
rect 4294 23950 4346 24002
rect 4358 23950 4410 24002
rect 4422 23950 4474 24002
rect 4486 23950 4538 24002
rect 35014 23950 35066 24002
rect 35078 23950 35130 24002
rect 35142 23950 35194 24002
rect 35206 23950 35258 24002
rect 1942 23691 1994 23743
rect 36886 23691 36938 23743
rect 8566 23586 8618 23595
rect 8566 23552 8575 23586
rect 8575 23552 8609 23586
rect 8609 23552 8618 23586
rect 8566 23543 8618 23552
rect 13654 23586 13706 23595
rect 13654 23552 13663 23586
rect 13663 23552 13697 23586
rect 13697 23552 13706 23586
rect 13654 23543 13706 23552
rect 26998 23469 27050 23521
rect 7126 23395 7178 23447
rect 19654 23284 19706 23336
rect 19718 23284 19770 23336
rect 19782 23284 19834 23336
rect 19846 23284 19898 23336
rect 50374 23284 50426 23336
rect 50438 23284 50490 23336
rect 50502 23284 50554 23336
rect 50566 23284 50618 23336
rect 57334 23025 57386 23077
rect 33814 22951 33866 23003
rect 38806 22951 38858 23003
rect 8758 22729 8810 22781
rect 19414 22729 19466 22781
rect 36310 22772 36362 22781
rect 36310 22738 36319 22772
rect 36319 22738 36353 22772
rect 36353 22738 36362 22772
rect 36310 22729 36362 22738
rect 49366 22729 49418 22781
rect 4294 22618 4346 22670
rect 4358 22618 4410 22670
rect 4422 22618 4474 22670
rect 4486 22618 4538 22670
rect 35014 22618 35066 22670
rect 35078 22618 35130 22670
rect 35142 22618 35194 22670
rect 35206 22618 35258 22670
rect 8566 22433 8618 22485
rect 33238 22433 33290 22485
rect 13654 22359 13706 22411
rect 40054 22359 40106 22411
rect 7894 22285 7946 22337
rect 54934 22285 54986 22337
rect 15094 22254 15146 22263
rect 15094 22220 15103 22254
rect 15103 22220 15137 22254
rect 15137 22220 15146 22254
rect 15094 22211 15146 22220
rect 22870 22211 22922 22263
rect 25558 22211 25610 22263
rect 19654 21952 19706 22004
rect 19718 21952 19770 22004
rect 19782 21952 19834 22004
rect 19846 21952 19898 22004
rect 50374 21952 50426 22004
rect 50438 21952 50490 22004
rect 50502 21952 50554 22004
rect 50566 21952 50618 22004
rect 26614 21619 26666 21671
rect 28150 21619 28202 21671
rect 38134 21545 38186 21597
rect 39478 21545 39530 21597
rect 9430 21397 9482 21449
rect 38422 21397 38474 21449
rect 4294 21286 4346 21338
rect 4358 21286 4410 21338
rect 4422 21286 4474 21338
rect 4486 21286 4538 21338
rect 35014 21286 35066 21338
rect 35078 21286 35130 21338
rect 35142 21286 35194 21338
rect 35206 21286 35258 21338
rect 13078 20953 13130 21005
rect 25078 21027 25130 21079
rect 26230 20879 26282 20931
rect 46774 20953 46826 21005
rect 19654 20620 19706 20672
rect 19718 20620 19770 20672
rect 19782 20620 19834 20672
rect 19846 20620 19898 20672
rect 50374 20620 50426 20672
rect 50438 20620 50490 20672
rect 50502 20620 50554 20672
rect 50566 20620 50618 20672
rect 24502 20139 24554 20191
rect 26710 20139 26762 20191
rect 5974 20065 6026 20117
rect 23158 20065 23210 20117
rect 4294 19954 4346 20006
rect 4358 19954 4410 20006
rect 4422 19954 4474 20006
rect 4486 19954 4538 20006
rect 35014 19954 35066 20006
rect 35078 19954 35130 20006
rect 35142 19954 35194 20006
rect 35206 19954 35258 20006
rect 19222 19769 19274 19821
rect 6166 19695 6218 19747
rect 20854 19695 20906 19747
rect 25654 19621 25706 19673
rect 4150 19547 4202 19599
rect 13942 19590 13994 19599
rect 6454 19473 6506 19525
rect 13942 19556 13951 19590
rect 13951 19556 13985 19590
rect 13985 19556 13994 19590
rect 13942 19547 13994 19556
rect 28246 19590 28298 19599
rect 28246 19556 28255 19590
rect 28255 19556 28289 19590
rect 28289 19556 28298 19590
rect 28246 19547 28298 19556
rect 5878 19399 5930 19451
rect 36790 19473 36842 19525
rect 17878 19399 17930 19451
rect 22870 19399 22922 19451
rect 49078 19399 49130 19451
rect 19654 19288 19706 19340
rect 19718 19288 19770 19340
rect 19782 19288 19834 19340
rect 19846 19288 19898 19340
rect 50374 19288 50426 19340
rect 50438 19288 50490 19340
rect 50502 19288 50554 19340
rect 50566 19288 50618 19340
rect 5974 19177 6026 19229
rect 5830 19103 5882 19155
rect 6118 19103 6170 19155
rect 6406 19103 6458 19155
rect 16054 19103 16106 19155
rect 47734 18955 47786 19007
rect 49942 18955 49994 19007
rect 30262 18733 30314 18785
rect 37654 18733 37706 18785
rect 4294 18622 4346 18674
rect 4358 18622 4410 18674
rect 4422 18622 4474 18674
rect 4486 18622 4538 18674
rect 35014 18622 35066 18674
rect 35078 18622 35130 18674
rect 35142 18622 35194 18674
rect 35206 18622 35258 18674
rect 28822 18215 28874 18267
rect 13942 18067 13994 18119
rect 46582 18067 46634 18119
rect 19654 17956 19706 18008
rect 19718 17956 19770 18008
rect 19782 17956 19834 18008
rect 19846 17956 19898 18008
rect 50374 17956 50426 18008
rect 50438 17956 50490 18008
rect 50502 17956 50554 18008
rect 50566 17956 50618 18008
rect 20758 17771 20810 17823
rect 23254 17771 23306 17823
rect 11926 17549 11978 17601
rect 37462 17475 37514 17527
rect 23158 17444 23210 17453
rect 23158 17410 23167 17444
rect 23167 17410 23201 17444
rect 23201 17410 23210 17444
rect 23158 17401 23210 17410
rect 41494 17401 41546 17453
rect 4294 17290 4346 17342
rect 4358 17290 4410 17342
rect 4422 17290 4474 17342
rect 4486 17290 4538 17342
rect 35014 17290 35066 17342
rect 35078 17290 35130 17342
rect 35142 17290 35194 17342
rect 35206 17290 35258 17342
rect 34390 16957 34442 17009
rect 16534 16883 16586 16935
rect 31510 16883 31562 16935
rect 29494 16809 29546 16861
rect 54646 16926 54698 16935
rect 54646 16892 54655 16926
rect 54655 16892 54689 16926
rect 54689 16892 54698 16926
rect 54646 16883 54698 16892
rect 10198 16735 10250 16787
rect 28822 16735 28874 16787
rect 38902 16735 38954 16787
rect 54454 16735 54506 16787
rect 19654 16624 19706 16676
rect 19718 16624 19770 16676
rect 19782 16624 19834 16676
rect 19846 16624 19898 16676
rect 50374 16624 50426 16676
rect 50438 16624 50490 16676
rect 50502 16624 50554 16676
rect 50566 16624 50618 16676
rect 19030 16513 19082 16565
rect 39862 16513 39914 16565
rect 21718 16069 21770 16121
rect 4294 15958 4346 16010
rect 4358 15958 4410 16010
rect 4422 15958 4474 16010
rect 4486 15958 4538 16010
rect 35014 15958 35066 16010
rect 35078 15958 35130 16010
rect 35142 15958 35194 16010
rect 35206 15958 35258 16010
rect 15862 15847 15914 15899
rect 15094 15699 15146 15751
rect 26422 15699 26474 15751
rect 22486 15625 22538 15677
rect 34870 15625 34922 15677
rect 18934 15551 18986 15603
rect 44662 15551 44714 15603
rect 15478 15477 15530 15529
rect 41302 15477 41354 15529
rect 18550 15403 18602 15455
rect 44950 15403 45002 15455
rect 19654 15292 19706 15344
rect 19718 15292 19770 15344
rect 19782 15292 19834 15344
rect 19846 15292 19898 15344
rect 50374 15292 50426 15344
rect 50438 15292 50490 15344
rect 50502 15292 50554 15344
rect 50566 15292 50618 15344
rect 18070 15181 18122 15233
rect 53974 15181 54026 15233
rect 15862 15107 15914 15159
rect 52630 15107 52682 15159
rect 32278 14780 32330 14789
rect 32278 14746 32287 14780
rect 32287 14746 32321 14780
rect 32321 14746 32330 14780
rect 32278 14737 32330 14746
rect 4294 14626 4346 14678
rect 4358 14626 4410 14678
rect 4422 14626 4474 14678
rect 4486 14626 4538 14678
rect 35014 14626 35066 14678
rect 35078 14626 35130 14678
rect 35142 14626 35194 14678
rect 35206 14626 35258 14678
rect 11542 14515 11594 14567
rect 17974 14515 18026 14567
rect 41206 14515 41258 14567
rect 42262 14515 42314 14567
rect 44758 14515 44810 14567
rect 12982 14441 13034 14493
rect 12598 14219 12650 14271
rect 34102 14219 34154 14271
rect 9430 14145 9482 14197
rect 24214 14145 24266 14197
rect 34582 14145 34634 14197
rect 41110 14145 41162 14197
rect 10102 14071 10154 14123
rect 19654 13960 19706 14012
rect 19718 13960 19770 14012
rect 19782 13960 19834 14012
rect 19846 13960 19898 14012
rect 50374 13960 50426 14012
rect 50438 13960 50490 14012
rect 50502 13960 50554 14012
rect 50566 13960 50618 14012
rect 33142 13849 33194 13901
rect 41398 13849 41450 13901
rect 12598 13775 12650 13827
rect 38422 13775 38474 13827
rect 52054 13775 52106 13827
rect 34006 13701 34058 13753
rect 54646 13701 54698 13753
rect 17974 13627 18026 13679
rect 47830 13553 47882 13605
rect 36598 13479 36650 13531
rect 4150 13405 4202 13457
rect 4294 13294 4346 13346
rect 4358 13294 4410 13346
rect 4422 13294 4474 13346
rect 4486 13294 4538 13346
rect 35014 13294 35066 13346
rect 35078 13294 35130 13346
rect 35142 13294 35194 13346
rect 35206 13294 35258 13346
rect 58198 13183 58250 13235
rect 21910 13035 21962 13087
rect 25462 13109 25514 13161
rect 25942 12961 25994 13013
rect 44086 13109 44138 13161
rect 41878 13035 41930 13087
rect 45622 13035 45674 13087
rect 41014 12961 41066 13013
rect 42934 12961 42986 13013
rect 50134 12961 50186 13013
rect 23446 12887 23498 12939
rect 45526 12887 45578 12939
rect 19654 12628 19706 12680
rect 19718 12628 19770 12680
rect 19782 12628 19834 12680
rect 19846 12628 19898 12680
rect 50374 12628 50426 12680
rect 50438 12628 50490 12680
rect 50502 12628 50554 12680
rect 50566 12628 50618 12680
rect 57142 12517 57194 12569
rect 13942 12443 13994 12495
rect 6070 12369 6122 12421
rect 29302 12369 29354 12421
rect 6262 12295 6314 12347
rect 56182 12295 56234 12347
rect 29590 12073 29642 12125
rect 42646 12147 42698 12199
rect 51574 12147 51626 12199
rect 57526 12147 57578 12199
rect 50230 12073 50282 12125
rect 4294 11962 4346 12014
rect 4358 11962 4410 12014
rect 4422 11962 4474 12014
rect 4486 11962 4538 12014
rect 35014 11962 35066 12014
rect 35078 11962 35130 12014
rect 35142 11962 35194 12014
rect 35206 11962 35258 12014
rect 7702 11851 7754 11903
rect 56182 11894 56234 11903
rect 56182 11860 56191 11894
rect 56191 11860 56225 11894
rect 56225 11860 56234 11894
rect 56182 11851 56234 11860
rect 23446 11777 23498 11829
rect 29302 11820 29354 11829
rect 29302 11786 29311 11820
rect 29311 11786 29345 11820
rect 29345 11786 29354 11820
rect 29302 11777 29354 11786
rect 23542 11703 23594 11755
rect 43030 11703 43082 11755
rect 58198 11777 58250 11829
rect 48118 11629 48170 11681
rect 55318 11629 55370 11681
rect 14614 11598 14666 11607
rect 14614 11564 14623 11598
rect 14623 11564 14657 11598
rect 14657 11564 14666 11598
rect 14614 11555 14666 11564
rect 56854 11555 56906 11607
rect 23254 11481 23306 11533
rect 19654 11296 19706 11348
rect 19718 11296 19770 11348
rect 19782 11296 19834 11348
rect 19846 11296 19898 11348
rect 50374 11296 50426 11348
rect 50438 11296 50490 11348
rect 50502 11296 50554 11348
rect 50566 11296 50618 11348
rect 21526 11185 21578 11237
rect 25366 11185 25418 11237
rect 43414 11185 43466 11237
rect 13846 11111 13898 11163
rect 25174 11111 25226 11163
rect 23926 11037 23978 11089
rect 37462 11037 37514 11089
rect 17590 10963 17642 11015
rect 38326 10963 38378 11015
rect 38518 10963 38570 11015
rect 4054 10889 4106 10941
rect 23254 10889 23306 10941
rect 36694 10889 36746 10941
rect 17782 10815 17834 10867
rect 38230 10815 38282 10867
rect 56374 10889 56426 10941
rect 57142 10815 57194 10867
rect 6934 10784 6986 10793
rect 6934 10750 6943 10784
rect 6943 10750 6977 10784
rect 6977 10750 6986 10784
rect 6934 10741 6986 10750
rect 32086 10741 32138 10793
rect 41110 10741 41162 10793
rect 54358 10784 54410 10793
rect 54358 10750 54367 10784
rect 54367 10750 54401 10784
rect 54401 10750 54410 10784
rect 54358 10741 54410 10750
rect 4294 10630 4346 10682
rect 4358 10630 4410 10682
rect 4422 10630 4474 10682
rect 4486 10630 4538 10682
rect 35014 10630 35066 10682
rect 35078 10630 35130 10682
rect 35142 10630 35194 10682
rect 35206 10630 35258 10682
rect 56278 10562 56330 10571
rect 56278 10528 56287 10562
rect 56287 10528 56321 10562
rect 56321 10528 56330 10562
rect 56278 10519 56330 10528
rect 6934 10445 6986 10497
rect 16150 10445 16202 10497
rect 31510 10445 31562 10497
rect 14230 10371 14282 10423
rect 25270 10371 25322 10423
rect 35350 10371 35402 10423
rect 36982 10371 37034 10423
rect 55030 10414 55082 10423
rect 55030 10380 55039 10414
rect 55039 10380 55073 10414
rect 55073 10380 55082 10414
rect 55030 10371 55082 10380
rect 55990 10371 56042 10423
rect 57430 10414 57482 10423
rect 57430 10380 57439 10414
rect 57439 10380 57473 10414
rect 57473 10380 57482 10414
rect 57430 10371 57482 10380
rect 20662 10297 20714 10349
rect 31222 10297 31274 10349
rect 52918 10297 52970 10349
rect 47830 10223 47882 10275
rect 17302 10149 17354 10201
rect 10774 10075 10826 10127
rect 12982 10075 13034 10127
rect 18454 10075 18506 10127
rect 19414 10075 19466 10127
rect 21046 10075 21098 10127
rect 31126 10149 31178 10201
rect 23446 10075 23498 10127
rect 25558 10075 25610 10127
rect 45334 10075 45386 10127
rect 47158 10075 47210 10127
rect 49654 10075 49706 10127
rect 50710 10075 50762 10127
rect 58582 10149 58634 10201
rect 55702 10075 55754 10127
rect 56086 10075 56138 10127
rect 56758 10075 56810 10127
rect 19654 9964 19706 10016
rect 19718 9964 19770 10016
rect 19782 9964 19834 10016
rect 19846 9964 19898 10016
rect 50374 9964 50426 10016
rect 50438 9964 50490 10016
rect 50502 9964 50554 10016
rect 50566 9964 50618 10016
rect 48598 9853 48650 9905
rect 14614 9779 14666 9831
rect 54166 9779 54218 9831
rect 5494 9705 5546 9757
rect 16822 9705 16874 9757
rect 28150 9705 28202 9757
rect 28534 9705 28586 9757
rect 32662 9705 32714 9757
rect 55894 9748 55946 9757
rect 55894 9714 55903 9748
rect 55903 9714 55937 9748
rect 55937 9714 55946 9748
rect 55894 9705 55946 9714
rect 39670 9631 39722 9683
rect 57622 9674 57674 9683
rect 57622 9640 57631 9674
rect 57631 9640 57665 9674
rect 57665 9640 57674 9674
rect 57622 9631 57674 9640
rect 42550 9557 42602 9609
rect 54262 9557 54314 9609
rect 54838 9557 54890 9609
rect 12502 9409 12554 9461
rect 55030 9483 55082 9535
rect 55318 9483 55370 9535
rect 45622 9452 45674 9461
rect 45622 9418 45631 9452
rect 45631 9418 45665 9452
rect 45665 9418 45674 9452
rect 45622 9409 45674 9418
rect 46774 9452 46826 9461
rect 46774 9418 46783 9452
rect 46783 9418 46817 9452
rect 46817 9418 46826 9452
rect 46774 9409 46826 9418
rect 4294 9298 4346 9350
rect 4358 9298 4410 9350
rect 4422 9298 4474 9350
rect 4486 9298 4538 9350
rect 35014 9298 35066 9350
rect 35078 9298 35130 9350
rect 35142 9298 35194 9350
rect 35206 9298 35258 9350
rect 28246 9187 28298 9239
rect 46774 9187 46826 9239
rect 54166 9187 54218 9239
rect 5494 9113 5546 9165
rect 46102 9113 46154 9165
rect 12310 9039 12362 9091
rect 53110 9082 53162 9091
rect 53110 9048 53119 9082
rect 53119 9048 53153 9082
rect 53153 9048 53162 9082
rect 55990 9113 56042 9165
rect 53110 9039 53162 9048
rect 53878 9039 53930 9091
rect 20470 8965 20522 9017
rect 56566 9008 56618 9017
rect 56566 8974 56575 9008
rect 56575 8974 56609 9008
rect 56609 8974 56618 9008
rect 56566 8965 56618 8974
rect 57238 9008 57290 9017
rect 57238 8974 57247 9008
rect 57247 8974 57281 9008
rect 57281 8974 57290 9008
rect 57238 8965 57290 8974
rect 14710 8891 14762 8943
rect 49174 8891 49226 8943
rect 54166 8891 54218 8943
rect 56374 8891 56426 8943
rect 56854 8891 56906 8943
rect 36694 8817 36746 8869
rect 51670 8743 51722 8795
rect 54550 8743 54602 8795
rect 19654 8632 19706 8684
rect 19718 8632 19770 8684
rect 19782 8632 19834 8684
rect 19846 8632 19898 8684
rect 50374 8632 50426 8684
rect 50438 8632 50490 8684
rect 50502 8632 50554 8684
rect 50566 8632 50618 8684
rect 2134 8564 2186 8573
rect 2134 8530 2143 8564
rect 2143 8530 2177 8564
rect 2177 8530 2186 8564
rect 2134 8521 2186 8530
rect 39190 8521 39242 8573
rect 42262 8564 42314 8573
rect 42262 8530 42271 8564
rect 42271 8530 42305 8564
rect 42305 8530 42314 8564
rect 42262 8521 42314 8530
rect 44086 8564 44138 8573
rect 44086 8530 44095 8564
rect 44095 8530 44129 8564
rect 44129 8530 44138 8564
rect 44086 8521 44138 8530
rect 48214 8564 48266 8573
rect 48214 8530 48223 8564
rect 48223 8530 48257 8564
rect 48257 8530 48266 8564
rect 48214 8521 48266 8530
rect 9334 8373 9386 8425
rect 10774 8416 10826 8425
rect 10774 8382 10783 8416
rect 10783 8382 10817 8416
rect 10817 8382 10826 8416
rect 10774 8373 10826 8382
rect 11542 8416 11594 8425
rect 11542 8382 11551 8416
rect 11551 8382 11585 8416
rect 11585 8382 11594 8416
rect 11542 8373 11594 8382
rect 12310 8416 12362 8425
rect 12310 8382 12319 8416
rect 12319 8382 12353 8416
rect 12353 8382 12362 8416
rect 12310 8373 12362 8382
rect 16150 8373 16202 8425
rect 17014 8416 17066 8425
rect 17014 8382 17023 8416
rect 17023 8382 17057 8416
rect 17057 8382 17066 8416
rect 17014 8373 17066 8382
rect 47926 8373 47978 8425
rect 52342 8521 52394 8573
rect 52918 8564 52970 8573
rect 52918 8530 52927 8564
rect 52927 8530 52961 8564
rect 52961 8530 52970 8564
rect 52918 8521 52970 8530
rect 49366 8416 49418 8425
rect 49366 8382 49375 8416
rect 49375 8382 49409 8416
rect 49409 8382 49418 8416
rect 49366 8373 49418 8382
rect 50134 8416 50186 8425
rect 50134 8382 50143 8416
rect 50143 8382 50177 8416
rect 50177 8382 50186 8416
rect 50134 8373 50186 8382
rect 54358 8373 54410 8425
rect 21334 8299 21386 8351
rect 53110 8299 53162 8351
rect 1654 8268 1706 8277
rect 1654 8234 1663 8268
rect 1663 8234 1697 8268
rect 1697 8234 1706 8268
rect 1654 8225 1706 8234
rect 2134 8225 2186 8277
rect 2998 8225 3050 8277
rect 4822 8225 4874 8277
rect 10582 8225 10634 8277
rect 10966 8225 11018 8277
rect 11734 8225 11786 8277
rect 12502 8225 12554 8277
rect 3670 8151 3722 8203
rect 16054 8225 16106 8277
rect 16342 8225 16394 8277
rect 39190 8225 39242 8277
rect 42358 8225 42410 8277
rect 44278 8225 44330 8277
rect 47638 8225 47690 8277
rect 48022 8225 48074 8277
rect 48694 8225 48746 8277
rect 49462 8225 49514 8277
rect 7510 8120 7562 8129
rect 7510 8086 7519 8120
rect 7519 8086 7553 8120
rect 7553 8086 7562 8120
rect 7510 8077 7562 8086
rect 12406 8077 12458 8129
rect 13750 8077 13802 8129
rect 15766 8077 15818 8129
rect 51094 8077 51146 8129
rect 53494 8225 53546 8277
rect 56950 8299 57002 8351
rect 58390 8225 58442 8277
rect 59830 8151 59882 8203
rect 58966 8077 59018 8129
rect 4294 7966 4346 8018
rect 4358 7966 4410 8018
rect 4422 7966 4474 8018
rect 4486 7966 4538 8018
rect 35014 7966 35066 8018
rect 35078 7966 35130 8018
rect 35142 7966 35194 8018
rect 35206 7966 35258 8018
rect 12406 7855 12458 7907
rect 12790 7898 12842 7907
rect 12790 7864 12799 7898
rect 12799 7864 12833 7898
rect 12833 7864 12842 7898
rect 12790 7855 12842 7864
rect 13558 7898 13610 7907
rect 13558 7864 13567 7898
rect 13567 7864 13601 7898
rect 13601 7864 13610 7898
rect 13558 7855 13610 7864
rect 14998 7855 15050 7907
rect 17974 7898 18026 7907
rect 17974 7864 17983 7898
rect 17983 7864 18017 7898
rect 18017 7864 18026 7898
rect 17974 7855 18026 7864
rect 27958 7898 28010 7907
rect 27958 7864 27967 7898
rect 27967 7864 28001 7898
rect 28001 7864 28010 7898
rect 30838 7898 30890 7907
rect 27958 7855 28010 7864
rect 3286 7707 3338 7759
rect 4054 7707 4106 7759
rect 23062 7781 23114 7833
rect 10198 7707 10250 7759
rect 10870 7750 10922 7759
rect 10870 7716 10879 7750
rect 10879 7716 10913 7750
rect 10913 7716 10922 7750
rect 10870 7707 10922 7716
rect 11350 7707 11402 7759
rect 12406 7750 12458 7759
rect 12406 7716 12415 7750
rect 12415 7716 12449 7750
rect 12449 7716 12458 7750
rect 12406 7707 12458 7716
rect 12790 7707 12842 7759
rect 13558 7707 13610 7759
rect 14998 7707 15050 7759
rect 16246 7750 16298 7759
rect 16246 7716 16255 7750
rect 16255 7716 16289 7750
rect 16289 7716 16298 7750
rect 16246 7707 16298 7716
rect 21046 7707 21098 7759
rect 23926 7750 23978 7759
rect 23926 7716 23935 7750
rect 23935 7716 23969 7750
rect 23969 7716 23978 7750
rect 23926 7707 23978 7716
rect 24694 7750 24746 7759
rect 24694 7716 24703 7750
rect 24703 7716 24737 7750
rect 24737 7716 24746 7750
rect 24694 7707 24746 7716
rect 25942 7707 25994 7759
rect 26230 7750 26282 7759
rect 26230 7716 26239 7750
rect 26239 7716 26273 7750
rect 26273 7716 26282 7750
rect 26230 7707 26282 7716
rect 26998 7750 27050 7759
rect 26998 7716 27007 7750
rect 27007 7716 27041 7750
rect 27041 7716 27050 7750
rect 26998 7707 27050 7716
rect 30838 7864 30847 7898
rect 30847 7864 30881 7898
rect 30881 7864 30890 7898
rect 30838 7855 30890 7864
rect 32374 7898 32426 7907
rect 32374 7864 32383 7898
rect 32383 7864 32417 7898
rect 32417 7864 32426 7898
rect 32374 7855 32426 7864
rect 35926 7855 35978 7907
rect 39958 7898 40010 7907
rect 29398 7750 29450 7759
rect 29398 7716 29407 7750
rect 29407 7716 29441 7750
rect 29441 7716 29450 7750
rect 29398 7707 29450 7716
rect 30166 7750 30218 7759
rect 30166 7716 30175 7750
rect 30175 7716 30209 7750
rect 30209 7716 30218 7750
rect 30166 7707 30218 7716
rect 34582 7750 34634 7759
rect 34582 7716 34591 7750
rect 34591 7716 34625 7750
rect 34625 7716 34634 7750
rect 34582 7707 34634 7716
rect 35350 7750 35402 7759
rect 35350 7716 35359 7750
rect 35359 7716 35393 7750
rect 35393 7716 35402 7750
rect 35350 7707 35402 7716
rect 39958 7864 39967 7898
rect 39967 7864 40001 7898
rect 40001 7864 40010 7898
rect 43702 7898 43754 7907
rect 39958 7855 40010 7864
rect 36790 7750 36842 7759
rect 36790 7716 36799 7750
rect 36799 7716 36833 7750
rect 36833 7716 36842 7750
rect 36790 7707 36842 7716
rect 38806 7750 38858 7759
rect 38806 7716 38815 7750
rect 38815 7716 38849 7750
rect 38849 7716 38858 7750
rect 38806 7707 38858 7716
rect 39478 7750 39530 7759
rect 39478 7716 39487 7750
rect 39487 7716 39521 7750
rect 39521 7716 39530 7750
rect 39478 7707 39530 7716
rect 43702 7864 43711 7898
rect 43711 7864 43745 7898
rect 43745 7864 43754 7898
rect 44470 7898 44522 7907
rect 43702 7855 43754 7864
rect 41110 7750 41162 7759
rect 41110 7716 41119 7750
rect 41119 7716 41153 7750
rect 41153 7716 41162 7750
rect 41110 7707 41162 7716
rect 41878 7750 41930 7759
rect 41878 7716 41887 7750
rect 41887 7716 41921 7750
rect 41921 7716 41930 7750
rect 41878 7707 41930 7716
rect 42646 7750 42698 7759
rect 42646 7716 42655 7750
rect 42655 7716 42689 7750
rect 42689 7716 42698 7750
rect 42646 7707 42698 7716
rect 44470 7864 44479 7898
rect 44479 7864 44513 7898
rect 44513 7864 44522 7898
rect 45238 7898 45290 7907
rect 44470 7855 44522 7864
rect 45238 7864 45247 7898
rect 45247 7864 45281 7898
rect 45281 7864 45290 7898
rect 46870 7898 46922 7907
rect 45238 7855 45290 7864
rect 46870 7864 46879 7898
rect 46879 7864 46913 7898
rect 46913 7864 46922 7898
rect 48982 7898 49034 7907
rect 46870 7855 46922 7864
rect 46390 7750 46442 7759
rect 46390 7716 46399 7750
rect 46399 7716 46433 7750
rect 46433 7716 46442 7750
rect 46390 7707 46442 7716
rect 48982 7864 48991 7898
rect 48991 7864 49025 7898
rect 49025 7864 49034 7898
rect 48982 7855 49034 7864
rect 49750 7898 49802 7907
rect 49750 7864 49759 7898
rect 49759 7864 49793 7898
rect 49793 7864 49802 7898
rect 49750 7855 49802 7864
rect 47830 7707 47882 7759
rect 51094 7750 51146 7759
rect 51094 7716 51103 7750
rect 51103 7716 51137 7750
rect 51137 7716 51146 7750
rect 51094 7707 51146 7716
rect 52630 7750 52682 7759
rect 52630 7716 52639 7750
rect 52639 7716 52673 7750
rect 52673 7716 52682 7750
rect 52630 7707 52682 7716
rect 52726 7707 52778 7759
rect 1462 7633 1514 7685
rect 3574 7633 3626 7685
rect 23158 7633 23210 7685
rect 53206 7633 53258 7685
rect 55798 7676 55850 7685
rect 4150 7559 4202 7611
rect 6838 7485 6890 7537
rect 12886 7559 12938 7611
rect 18358 7559 18410 7611
rect 34102 7559 34154 7611
rect 52918 7559 52970 7611
rect 55798 7642 55807 7676
rect 55807 7642 55841 7676
rect 55841 7642 55850 7676
rect 55798 7633 55850 7642
rect 56182 7633 56234 7685
rect 57334 7676 57386 7685
rect 57334 7642 57343 7676
rect 57343 7642 57377 7676
rect 57377 7642 57386 7676
rect 57334 7633 57386 7642
rect 58774 7559 58826 7611
rect 2422 7454 2474 7463
rect 2422 7420 2431 7454
rect 2431 7420 2465 7454
rect 2465 7420 2474 7454
rect 2422 7411 2474 7420
rect 3382 7411 3434 7463
rect 5302 7411 5354 7463
rect 9142 7411 9194 7463
rect 9910 7411 9962 7463
rect 11062 7411 11114 7463
rect 12214 7411 12266 7463
rect 39958 7485 40010 7537
rect 15286 7411 15338 7463
rect 15670 7411 15722 7463
rect 20758 7411 20810 7463
rect 23734 7411 23786 7463
rect 24598 7454 24650 7463
rect 24598 7420 24607 7454
rect 24607 7420 24641 7454
rect 24641 7420 24650 7454
rect 24598 7411 24650 7420
rect 24790 7411 24842 7463
rect 25942 7411 25994 7463
rect 26710 7411 26762 7463
rect 28150 7411 28202 7463
rect 29206 7411 29258 7463
rect 29590 7411 29642 7463
rect 31030 7411 31082 7463
rect 33622 7411 33674 7463
rect 34390 7411 34442 7463
rect 34774 7411 34826 7463
rect 36022 7411 36074 7463
rect 36598 7411 36650 7463
rect 38038 7411 38090 7463
rect 38806 7411 38858 7463
rect 39670 7411 39722 7463
rect 41686 7485 41738 7537
rect 41110 7411 41162 7463
rect 45430 7485 45482 7537
rect 43222 7411 43274 7463
rect 44374 7411 44426 7463
rect 45046 7411 45098 7463
rect 46870 7485 46922 7537
rect 46390 7411 46442 7463
rect 48310 7411 48362 7463
rect 50038 7411 50090 7463
rect 59350 7485 59402 7537
rect 51670 7411 51722 7463
rect 52342 7411 52394 7463
rect 19654 7300 19706 7352
rect 19718 7300 19770 7352
rect 19782 7300 19834 7352
rect 19846 7300 19898 7352
rect 50374 7300 50426 7352
rect 50438 7300 50490 7352
rect 50502 7300 50554 7352
rect 50566 7300 50618 7352
rect 6454 7158 6506 7167
rect 6454 7124 6463 7158
rect 6463 7124 6497 7158
rect 6497 7124 6506 7158
rect 7990 7158 8042 7167
rect 6454 7115 6506 7124
rect 7990 7124 7999 7158
rect 7999 7124 8033 7158
rect 8033 7124 8042 7158
rect 7990 7115 8042 7124
rect 7606 7084 7658 7093
rect 7606 7050 7615 7084
rect 7615 7050 7649 7084
rect 7649 7050 7658 7084
rect 7606 7041 7658 7050
rect 17110 7115 17162 7167
rect 22294 7158 22346 7167
rect 15190 7041 15242 7093
rect 15766 7041 15818 7093
rect 16534 7041 16586 7093
rect 18070 7084 18122 7093
rect 18070 7050 18079 7084
rect 18079 7050 18113 7084
rect 18113 7050 18122 7084
rect 18070 7041 18122 7050
rect 18838 7084 18890 7093
rect 18838 7050 18847 7084
rect 18847 7050 18881 7084
rect 18881 7050 18890 7084
rect 18838 7041 18890 7050
rect 20374 7084 20426 7093
rect 20374 7050 20383 7084
rect 20383 7050 20417 7084
rect 20417 7050 20426 7084
rect 20374 7041 20426 7050
rect 22294 7124 22303 7158
rect 22303 7124 22337 7158
rect 22337 7124 22346 7158
rect 22294 7115 22346 7124
rect 21910 7084 21962 7093
rect 21910 7050 21919 7084
rect 21919 7050 21953 7084
rect 21953 7050 21962 7084
rect 21910 7041 21962 7050
rect 23062 7115 23114 7167
rect 28054 7115 28106 7167
rect 28342 7158 28394 7167
rect 28342 7124 28351 7158
rect 28351 7124 28385 7158
rect 28385 7124 28394 7158
rect 28342 7115 28394 7124
rect 23446 7084 23498 7093
rect 23446 7050 23455 7084
rect 23455 7050 23489 7084
rect 23489 7050 23498 7084
rect 23446 7041 23498 7050
rect 24214 7084 24266 7093
rect 24214 7050 24223 7084
rect 24223 7050 24257 7084
rect 24257 7050 24266 7084
rect 24214 7041 24266 7050
rect 25654 7084 25706 7093
rect 25654 7050 25663 7084
rect 25663 7050 25697 7084
rect 25697 7050 25706 7084
rect 25654 7041 25706 7050
rect 26422 7084 26474 7093
rect 26422 7050 26431 7084
rect 26431 7050 26465 7084
rect 26465 7050 26474 7084
rect 26422 7041 26474 7050
rect 27190 7084 27242 7093
rect 27190 7050 27199 7084
rect 27199 7050 27233 7084
rect 27233 7050 27242 7084
rect 27190 7041 27242 7050
rect 28246 7041 28298 7093
rect 30742 7115 30794 7167
rect 32950 7189 33002 7241
rect 35446 7115 35498 7167
rect 38902 7158 38954 7167
rect 29494 7084 29546 7093
rect 29494 7050 29503 7084
rect 29503 7050 29537 7084
rect 29537 7050 29546 7084
rect 29494 7041 29546 7050
rect 31702 7084 31754 7093
rect 31702 7050 31711 7084
rect 31711 7050 31745 7084
rect 31745 7050 31754 7084
rect 31702 7041 31754 7050
rect 32470 7084 32522 7093
rect 32470 7050 32479 7084
rect 32479 7050 32513 7084
rect 32513 7050 32522 7084
rect 32470 7041 32522 7050
rect 33238 7084 33290 7093
rect 33238 7050 33247 7084
rect 33247 7050 33281 7084
rect 33281 7050 33290 7084
rect 33238 7041 33290 7050
rect 34006 7084 34058 7093
rect 34006 7050 34015 7084
rect 34015 7050 34049 7084
rect 34049 7050 34058 7084
rect 34006 7041 34058 7050
rect 36886 7084 36938 7093
rect 36886 7050 36895 7084
rect 36895 7050 36929 7084
rect 36929 7050 36938 7084
rect 36886 7041 36938 7050
rect 37654 7084 37706 7093
rect 37654 7050 37663 7084
rect 37663 7050 37697 7084
rect 37697 7050 37706 7084
rect 37654 7041 37706 7050
rect 38902 7124 38911 7158
rect 38911 7124 38945 7158
rect 38945 7124 38954 7158
rect 38902 7115 38954 7124
rect 40630 7115 40682 7167
rect 40054 7084 40106 7093
rect 40054 7050 40063 7084
rect 40063 7050 40097 7084
rect 40097 7050 40106 7084
rect 40054 7041 40106 7050
rect 41494 7084 41546 7093
rect 41494 7050 41503 7084
rect 41503 7050 41537 7084
rect 41537 7050 41546 7084
rect 41494 7041 41546 7050
rect 42934 7084 42986 7093
rect 42934 7050 42943 7084
rect 42943 7050 42977 7084
rect 42977 7050 42986 7084
rect 42934 7041 42986 7050
rect 43126 7041 43178 7093
rect 44566 7084 44618 7093
rect 44566 7050 44575 7084
rect 44575 7050 44609 7084
rect 44609 7050 44618 7084
rect 44566 7041 44618 7050
rect 46582 7041 46634 7093
rect 47158 7084 47210 7093
rect 47158 7050 47167 7084
rect 47167 7050 47201 7084
rect 47201 7050 47210 7084
rect 47158 7041 47210 7050
rect 48118 7041 48170 7093
rect 49078 7084 49130 7093
rect 49078 7050 49087 7084
rect 49087 7050 49121 7084
rect 49121 7050 49130 7084
rect 49078 7041 49130 7050
rect 49942 7041 49994 7093
rect 52054 7084 52106 7093
rect 52054 7050 52063 7084
rect 52063 7050 52097 7084
rect 52097 7050 52106 7084
rect 52054 7041 52106 7050
rect 52438 7084 52490 7093
rect 52438 7050 52447 7084
rect 52447 7050 52481 7084
rect 52481 7050 52490 7084
rect 52438 7041 52490 7050
rect 56374 7115 56426 7167
rect 56758 7115 56810 7167
rect 54358 7041 54410 7093
rect 1654 7010 1706 7019
rect 1654 6976 1663 7010
rect 1663 6976 1697 7010
rect 1697 6976 1706 7010
rect 1654 6967 1706 6976
rect 2518 7010 2570 7019
rect 2518 6976 2527 7010
rect 2527 6976 2561 7010
rect 2561 6976 2570 7010
rect 2518 6967 2570 6976
rect 11254 7010 11306 7019
rect 5110 6893 5162 6945
rect 3670 6819 3722 6871
rect 5686 6893 5738 6945
rect 5878 6893 5930 6945
rect 6166 6893 6218 6945
rect 6550 6893 6602 6945
rect 11254 6976 11263 7010
rect 11263 6976 11297 7010
rect 11297 6976 11306 7010
rect 11254 6967 11306 6976
rect 12694 7010 12746 7019
rect 12694 6976 12703 7010
rect 12703 6976 12737 7010
rect 12737 6976 12746 7010
rect 12694 6967 12746 6976
rect 7318 6893 7370 6945
rect 8086 6893 8138 6945
rect 8854 6893 8906 6945
rect 9526 6819 9578 6871
rect 13462 6893 13514 6945
rect 13654 6936 13706 6945
rect 13654 6902 13663 6936
rect 13663 6902 13697 6936
rect 13697 6902 13706 6936
rect 13654 6893 13706 6902
rect 14518 6893 14570 6945
rect 15094 6893 15146 6945
rect 17302 6936 17354 6945
rect 17302 6902 17311 6936
rect 17311 6902 17345 6936
rect 17345 6902 17354 6936
rect 17302 6893 17354 6902
rect 17878 6893 17930 6945
rect 18646 6893 18698 6945
rect 20374 6893 20426 6945
rect 20854 6893 20906 6945
rect 21238 6893 21290 6945
rect 21910 6893 21962 6945
rect 23638 6967 23690 7019
rect 25174 6967 25226 7019
rect 23926 6893 23978 6945
rect 24118 6936 24170 6945
rect 24118 6902 24127 6936
rect 24127 6902 24161 6936
rect 24161 6902 24170 6936
rect 24118 6893 24170 6902
rect 24886 6893 24938 6945
rect 27766 6967 27818 7019
rect 27094 6936 27146 6945
rect 27094 6902 27103 6936
rect 27103 6902 27137 6936
rect 27137 6902 27146 6936
rect 27094 6893 27146 6902
rect 27382 6893 27434 6945
rect 32278 6967 32330 7019
rect 45622 6967 45674 7019
rect 46486 6967 46538 7019
rect 29398 6936 29450 6945
rect 29398 6902 29407 6936
rect 29407 6902 29441 6936
rect 29441 6902 29450 6936
rect 29398 6893 29450 6902
rect 29974 6893 30026 6945
rect 31414 6893 31466 6945
rect 32470 6893 32522 6945
rect 34006 6893 34058 6945
rect 35350 6893 35402 6945
rect 35542 6893 35594 6945
rect 36502 6893 36554 6945
rect 37078 6893 37130 6945
rect 23062 6745 23114 6797
rect 37270 6819 37322 6871
rect 37366 6819 37418 6871
rect 23926 6745 23978 6797
rect 34678 6745 34730 6797
rect 37654 6745 37706 6797
rect 39286 6893 39338 6945
rect 39862 6819 39914 6871
rect 41590 6893 41642 6945
rect 43798 6936 43850 6945
rect 43798 6902 43807 6936
rect 43807 6902 43841 6936
rect 43841 6902 43850 6936
rect 43798 6893 43850 6902
rect 42742 6819 42794 6871
rect 43606 6745 43658 6797
rect 45814 6893 45866 6945
rect 54742 7010 54794 7019
rect 45718 6819 45770 6871
rect 47254 6819 47306 6871
rect 50134 6893 50186 6945
rect 51286 6893 51338 6945
rect 52822 6936 52874 6945
rect 52822 6902 52831 6936
rect 52831 6902 52865 6936
rect 52865 6902 52874 6936
rect 52822 6893 52874 6902
rect 54742 6976 54751 7010
rect 54751 6976 54785 7010
rect 54785 6976 54794 7010
rect 54742 6967 54794 6976
rect 55414 6967 55466 7019
rect 58486 6967 58538 7019
rect 56278 6893 56330 6945
rect 49174 6745 49226 6797
rect 4294 6634 4346 6686
rect 4358 6634 4410 6686
rect 4422 6634 4474 6686
rect 4486 6634 4538 6686
rect 35014 6634 35066 6686
rect 35078 6634 35130 6686
rect 35142 6634 35194 6686
rect 35206 6634 35258 6686
rect 6166 6523 6218 6575
rect 12118 6523 12170 6575
rect 19030 6523 19082 6575
rect 33142 6566 33194 6575
rect 33142 6532 33151 6566
rect 33151 6532 33185 6566
rect 33185 6532 33194 6566
rect 33142 6523 33194 6532
rect 36694 6523 36746 6575
rect 38422 6523 38474 6575
rect 39286 6523 39338 6575
rect 50710 6523 50762 6575
rect 7126 6418 7178 6427
rect 7126 6384 7135 6418
rect 7135 6384 7169 6418
rect 7169 6384 7178 6418
rect 7126 6375 7178 6384
rect 8470 6375 8522 6427
rect 13942 6418 13994 6427
rect 13942 6384 13951 6418
rect 13951 6384 13985 6418
rect 13985 6384 13994 6418
rect 13942 6375 13994 6384
rect 14710 6418 14762 6427
rect 14710 6384 14719 6418
rect 14719 6384 14753 6418
rect 14753 6384 14762 6418
rect 14710 6375 14762 6384
rect 15478 6418 15530 6427
rect 15478 6384 15487 6418
rect 15487 6384 15521 6418
rect 15521 6384 15530 6418
rect 15478 6375 15530 6384
rect 1558 6344 1610 6353
rect 1558 6310 1567 6344
rect 1567 6310 1601 6344
rect 1601 6310 1610 6344
rect 1558 6301 1610 6310
rect 2038 6301 2090 6353
rect 3190 6344 3242 6353
rect 3190 6310 3199 6344
rect 3199 6310 3233 6344
rect 3233 6310 3242 6344
rect 3190 6301 3242 6310
rect 3862 6301 3914 6353
rect 4630 6301 4682 6353
rect 8758 6301 8810 6353
rect 10102 6344 10154 6353
rect 10102 6310 10111 6344
rect 10111 6310 10145 6344
rect 10145 6310 10154 6344
rect 10102 6301 10154 6310
rect 10870 6344 10922 6353
rect 10870 6310 10879 6344
rect 10879 6310 10913 6344
rect 10913 6310 10922 6344
rect 10870 6301 10922 6310
rect 11638 6301 11690 6353
rect 12310 6301 12362 6353
rect 16438 6375 16490 6427
rect 18454 6418 18506 6427
rect 18454 6384 18463 6418
rect 18463 6384 18497 6418
rect 18497 6384 18506 6418
rect 18454 6375 18506 6384
rect 19030 6375 19082 6427
rect 19990 6418 20042 6427
rect 19990 6384 19999 6418
rect 19999 6384 20033 6418
rect 20033 6384 20042 6418
rect 19990 6375 20042 6384
rect 20950 6375 21002 6427
rect 21526 6418 21578 6427
rect 21526 6384 21535 6418
rect 21535 6384 21569 6418
rect 21569 6384 21578 6418
rect 21526 6375 21578 6384
rect 22966 6418 23018 6427
rect 22966 6384 22975 6418
rect 22975 6384 23009 6418
rect 23009 6384 23018 6418
rect 22966 6375 23018 6384
rect 23254 6375 23306 6427
rect 24502 6418 24554 6427
rect 24502 6384 24511 6418
rect 24511 6384 24545 6418
rect 24545 6384 24554 6418
rect 24502 6375 24554 6384
rect 28534 6375 28586 6427
rect 29014 6418 29066 6427
rect 29014 6384 29023 6418
rect 29023 6384 29057 6418
rect 29057 6384 29066 6418
rect 29014 6375 29066 6384
rect 30646 6418 30698 6427
rect 30646 6384 30655 6418
rect 30655 6384 30689 6418
rect 30689 6384 30698 6418
rect 30646 6375 30698 6384
rect 32086 6375 32138 6427
rect 37270 6449 37322 6501
rect 42070 6449 42122 6501
rect 46966 6449 47018 6501
rect 47158 6449 47210 6501
rect 47350 6375 47402 6427
rect 51478 6375 51530 6427
rect 8566 6227 8618 6279
rect 16534 6301 16586 6353
rect 25654 6344 25706 6353
rect 25654 6310 25663 6344
rect 25663 6310 25697 6344
rect 25697 6310 25706 6344
rect 25654 6301 25706 6310
rect 26806 6344 26858 6353
rect 26806 6310 26815 6344
rect 26815 6310 26849 6344
rect 26849 6310 26858 6344
rect 26806 6301 26858 6310
rect 29686 6344 29738 6353
rect 29686 6310 29695 6344
rect 29695 6310 29729 6344
rect 29729 6310 29738 6344
rect 29686 6301 29738 6310
rect 31222 6344 31274 6353
rect 31222 6310 31231 6344
rect 31231 6310 31265 6344
rect 31265 6310 31274 6344
rect 31222 6301 31274 6310
rect 32566 6301 32618 6353
rect 36310 6344 36362 6353
rect 36310 6310 36319 6344
rect 36319 6310 36353 6344
rect 36353 6310 36362 6344
rect 36310 6301 36362 6310
rect 17686 6270 17738 6279
rect 17686 6236 17695 6270
rect 17695 6236 17729 6270
rect 17729 6236 17738 6270
rect 17686 6227 17738 6236
rect 18070 6227 18122 6279
rect 6934 6153 6986 6205
rect 5494 6079 5546 6131
rect 6262 6079 6314 6131
rect 7990 6153 8042 6205
rect 14134 6153 14186 6205
rect 13270 6079 13322 6131
rect 13942 6079 13994 6131
rect 17494 6153 17546 6205
rect 16726 6079 16778 6131
rect 33142 6227 33194 6279
rect 34294 6270 34346 6279
rect 34294 6236 34303 6270
rect 34303 6236 34337 6270
rect 34337 6236 34346 6270
rect 34294 6227 34346 6236
rect 22294 6153 22346 6205
rect 19318 6079 19370 6131
rect 19990 6079 20042 6131
rect 21430 6122 21482 6131
rect 21430 6088 21439 6122
rect 21439 6088 21473 6122
rect 21473 6088 21482 6122
rect 21430 6079 21482 6088
rect 22870 6122 22922 6131
rect 22870 6088 22879 6122
rect 22879 6088 22913 6122
rect 22913 6088 22922 6122
rect 22870 6079 22922 6088
rect 31798 6153 31850 6205
rect 35734 6227 35786 6279
rect 38902 6344 38954 6353
rect 38902 6310 38911 6344
rect 38911 6310 38945 6344
rect 38945 6310 38954 6344
rect 38902 6301 38954 6310
rect 40342 6344 40394 6353
rect 40342 6310 40351 6344
rect 40351 6310 40385 6344
rect 40385 6310 40394 6344
rect 40342 6301 40394 6310
rect 41494 6344 41546 6353
rect 41494 6310 41503 6344
rect 41503 6310 41537 6344
rect 41537 6310 41546 6344
rect 41494 6301 41546 6310
rect 41878 6301 41930 6353
rect 43318 6301 43370 6353
rect 44758 6344 44810 6353
rect 44758 6310 44767 6344
rect 44767 6310 44801 6344
rect 44801 6310 44810 6344
rect 44758 6301 44810 6310
rect 45526 6344 45578 6353
rect 45526 6310 45535 6344
rect 45535 6310 45569 6344
rect 45569 6310 45578 6344
rect 45526 6301 45578 6310
rect 46966 6344 47018 6353
rect 46966 6310 46975 6344
rect 46975 6310 47009 6344
rect 47009 6310 47018 6344
rect 46966 6301 47018 6310
rect 47734 6344 47786 6353
rect 47734 6310 47743 6344
rect 47743 6310 47777 6344
rect 47777 6310 47786 6344
rect 47734 6301 47786 6310
rect 48790 6301 48842 6353
rect 49558 6301 49610 6353
rect 51574 6301 51626 6353
rect 56854 6375 56906 6427
rect 53974 6301 54026 6353
rect 54646 6301 54698 6353
rect 36694 6227 36746 6279
rect 51190 6227 51242 6279
rect 55126 6227 55178 6279
rect 58102 6301 58154 6353
rect 58870 6227 58922 6279
rect 24310 6079 24362 6131
rect 27574 6079 27626 6131
rect 29302 6079 29354 6131
rect 29782 6079 29834 6131
rect 30646 6079 30698 6131
rect 45334 6153 45386 6205
rect 33526 6079 33578 6131
rect 49750 6079 49802 6131
rect 51094 6079 51146 6131
rect 19654 5968 19706 6020
rect 19718 5968 19770 6020
rect 19782 5968 19834 6020
rect 19846 5968 19898 6020
rect 50374 5968 50426 6020
rect 50438 5968 50490 6020
rect 50502 5968 50554 6020
rect 50566 5968 50618 6020
rect 5686 5783 5738 5835
rect 36214 5857 36266 5909
rect 54934 5857 54986 5909
rect 23350 5783 23402 5835
rect 24118 5783 24170 5835
rect 43030 5783 43082 5835
rect 56278 5783 56330 5835
rect 57718 5783 57770 5835
rect 6070 5752 6122 5761
rect 6070 5718 6079 5752
rect 6079 5718 6113 5752
rect 6113 5718 6122 5752
rect 6070 5709 6122 5718
rect 7510 5709 7562 5761
rect 34294 5709 34346 5761
rect 1078 5635 1130 5687
rect 2902 5678 2954 5687
rect 2902 5644 2911 5678
rect 2911 5644 2945 5678
rect 2945 5644 2954 5678
rect 2902 5635 2954 5644
rect 4918 5635 4970 5687
rect 5110 5678 5162 5687
rect 5110 5644 5119 5678
rect 5119 5644 5153 5678
rect 5153 5644 5162 5678
rect 5110 5635 5162 5644
rect 7222 5678 7274 5687
rect 7222 5644 7231 5678
rect 7231 5644 7265 5678
rect 7265 5644 7274 5678
rect 7222 5635 7274 5644
rect 7894 5635 7946 5687
rect 9046 5635 9098 5687
rect 10198 5635 10250 5687
rect 10486 5635 10538 5687
rect 12598 5678 12650 5687
rect 12598 5644 12607 5678
rect 12607 5644 12641 5678
rect 12641 5644 12650 5678
rect 12598 5635 12650 5644
rect 13366 5678 13418 5687
rect 13366 5644 13375 5678
rect 13375 5644 13409 5678
rect 13409 5644 13418 5678
rect 13366 5635 13418 5644
rect 14998 5678 15050 5687
rect 14998 5644 15007 5678
rect 15007 5644 15041 5678
rect 15041 5644 15050 5678
rect 14998 5635 15050 5644
rect 15862 5678 15914 5687
rect 15862 5644 15871 5678
rect 15871 5644 15905 5678
rect 15905 5644 15914 5678
rect 15862 5635 15914 5644
rect 16150 5635 16202 5687
rect 17974 5678 18026 5687
rect 17974 5644 17983 5678
rect 17983 5644 18017 5678
rect 18017 5644 18026 5678
rect 17974 5635 18026 5644
rect 18742 5678 18794 5687
rect 18742 5644 18751 5678
rect 18751 5644 18785 5678
rect 18785 5644 18794 5678
rect 18742 5635 18794 5644
rect 20182 5678 20234 5687
rect 20182 5644 20191 5678
rect 20191 5644 20225 5678
rect 20225 5644 20234 5678
rect 20182 5635 20234 5644
rect 20470 5635 20522 5687
rect 21718 5678 21770 5687
rect 21718 5644 21727 5678
rect 21727 5644 21761 5678
rect 21761 5644 21770 5678
rect 21718 5635 21770 5644
rect 22486 5678 22538 5687
rect 22486 5644 22495 5678
rect 22495 5644 22529 5678
rect 22529 5644 22538 5678
rect 22486 5635 22538 5644
rect 23062 5635 23114 5687
rect 23446 5635 23498 5687
rect 24598 5635 24650 5687
rect 26230 5678 26282 5687
rect 26230 5644 26239 5678
rect 26239 5644 26273 5678
rect 26273 5644 26282 5678
rect 26230 5635 26282 5644
rect 5974 5604 6026 5613
rect 5974 5570 5983 5604
rect 5983 5570 6017 5604
rect 6017 5570 6026 5604
rect 5974 5561 6026 5570
rect 26038 5561 26090 5613
rect 27190 5635 27242 5687
rect 27862 5635 27914 5687
rect 28822 5635 28874 5687
rect 30262 5635 30314 5687
rect 30838 5635 30890 5687
rect 31702 5635 31754 5687
rect 33142 5678 33194 5687
rect 33142 5644 33151 5678
rect 33151 5644 33185 5678
rect 33185 5644 33194 5678
rect 33142 5635 33194 5644
rect 34678 5678 34730 5687
rect 33238 5561 33290 5613
rect 34678 5644 34687 5678
rect 34687 5644 34721 5678
rect 34721 5644 34730 5678
rect 34678 5635 34730 5644
rect 36214 5635 36266 5687
rect 36406 5635 36458 5687
rect 37558 5678 37610 5687
rect 37558 5644 37567 5678
rect 37567 5644 37601 5678
rect 37601 5644 37610 5678
rect 37558 5635 37610 5644
rect 39094 5678 39146 5687
rect 37462 5561 37514 5613
rect 39094 5644 39103 5678
rect 39103 5644 39137 5678
rect 39137 5644 39146 5678
rect 39094 5635 39146 5644
rect 39286 5635 39338 5687
rect 40726 5635 40778 5687
rect 42598 5598 42650 5650
rect 42886 5598 42938 5650
rect 43510 5635 43562 5687
rect 44662 5678 44714 5687
rect 44662 5644 44671 5678
rect 44671 5644 44705 5678
rect 44705 5644 44714 5678
rect 44662 5635 44714 5644
rect 46102 5635 46154 5687
rect 46678 5635 46730 5687
rect 47542 5635 47594 5687
rect 48982 5678 49034 5687
rect 48982 5644 48991 5678
rect 48991 5644 49025 5678
rect 49025 5644 49034 5678
rect 48982 5635 49034 5644
rect 49654 5678 49706 5687
rect 49654 5644 49663 5678
rect 49663 5644 49697 5678
rect 49697 5644 49706 5678
rect 49654 5635 49706 5644
rect 50710 5635 50762 5687
rect 52150 5678 52202 5687
rect 52150 5644 52159 5678
rect 52159 5644 52193 5678
rect 52193 5644 52202 5678
rect 52150 5635 52202 5644
rect 52534 5635 52586 5687
rect 53686 5678 53738 5687
rect 53686 5644 53695 5678
rect 53695 5644 53729 5678
rect 53729 5644 53738 5678
rect 53686 5635 53738 5644
rect 57430 5678 57482 5687
rect 53590 5561 53642 5613
rect 57430 5644 57439 5678
rect 57439 5644 57473 5678
rect 57473 5644 57482 5678
rect 57430 5635 57482 5644
rect 59638 5561 59690 5613
rect 17686 5487 17738 5539
rect 12118 5456 12170 5465
rect 12118 5422 12127 5456
rect 12127 5422 12161 5456
rect 12161 5422 12170 5456
rect 12118 5413 12170 5422
rect 28438 5413 28490 5465
rect 37846 5413 37898 5465
rect 42598 5413 42650 5465
rect 4294 5302 4346 5354
rect 4358 5302 4410 5354
rect 4422 5302 4474 5354
rect 4486 5302 4538 5354
rect 35014 5302 35066 5354
rect 35078 5302 35130 5354
rect 35142 5302 35194 5354
rect 35206 5302 35258 5354
rect 18358 5191 18410 5243
rect 43798 5191 43850 5243
rect 12118 5043 12170 5095
rect 47062 5043 47114 5095
rect 310 4969 362 5021
rect 1846 4969 1898 5021
rect 3094 5012 3146 5021
rect 3094 4978 3103 5012
rect 3103 4978 3137 5012
rect 3137 4978 3146 5012
rect 3094 4969 3146 4978
rect 4150 5012 4202 5021
rect 4150 4978 4159 5012
rect 4159 4978 4193 5012
rect 4193 4978 4202 5012
rect 4150 4969 4202 4978
rect 5398 5012 5450 5021
rect 5398 4978 5407 5012
rect 5407 4978 5441 5012
rect 5441 4978 5450 5012
rect 5398 4969 5450 4978
rect 6070 4969 6122 5021
rect 7702 5012 7754 5021
rect 7702 4978 7711 5012
rect 7711 4978 7745 5012
rect 7745 4978 7754 5012
rect 7702 4969 7754 4978
rect 9238 5012 9290 5021
rect 7606 4895 7658 4947
rect 9238 4978 9247 5012
rect 9247 4978 9281 5012
rect 9281 4978 9290 5012
rect 9238 4969 9290 4978
rect 10294 4969 10346 5021
rect 10678 4969 10730 5021
rect 11830 4969 11882 5021
rect 12982 5012 13034 5021
rect 12982 4978 12991 5012
rect 12991 4978 13025 5012
rect 13025 4978 13034 5012
rect 13942 5012 13994 5021
rect 12982 4969 13034 4978
rect 13942 4978 13951 5012
rect 13951 4978 13985 5012
rect 13985 4978 13994 5012
rect 13942 4969 13994 4978
rect 14422 4969 14474 5021
rect 14806 4969 14858 5021
rect 16438 4969 16490 5021
rect 17302 4969 17354 5021
rect 17590 4969 17642 5021
rect 19030 5012 19082 5021
rect 19030 4978 19039 5012
rect 19039 4978 19073 5012
rect 19073 4978 19082 5012
rect 19030 4969 19082 4978
rect 19222 4969 19274 5021
rect 20566 5012 20618 5021
rect 20566 4978 20575 5012
rect 20575 4978 20609 5012
rect 20609 4978 20618 5012
rect 20566 4969 20618 4978
rect 21238 4969 21290 5021
rect 22774 5012 22826 5021
rect 22774 4978 22783 5012
rect 22783 4978 22817 5012
rect 22817 4978 22826 5012
rect 22774 4969 22826 4978
rect 23158 4969 23210 5021
rect 23830 4969 23882 5021
rect 24406 4969 24458 5021
rect 25846 5012 25898 5021
rect 25846 4978 25855 5012
rect 25855 4978 25889 5012
rect 25889 4978 25898 5012
rect 25846 4969 25898 4978
rect 26614 5012 26666 5021
rect 26614 4978 26623 5012
rect 26623 4978 26657 5012
rect 26657 4978 26666 5012
rect 26614 4969 26666 4978
rect 28918 5012 28970 5021
rect 28918 4978 28927 5012
rect 28927 4978 28961 5012
rect 28961 4978 28970 5012
rect 28918 4969 28970 4978
rect 29014 4969 29066 5021
rect 30358 5012 30410 5021
rect 30358 4978 30367 5012
rect 30367 4978 30401 5012
rect 30401 4978 30410 5012
rect 30358 4969 30410 4978
rect 31126 5012 31178 5021
rect 31126 4978 31135 5012
rect 31135 4978 31169 5012
rect 31169 4978 31178 5012
rect 31126 4969 31178 4978
rect 31894 5012 31946 5021
rect 31894 4978 31903 5012
rect 31903 4978 31937 5012
rect 31937 4978 31946 5012
rect 31894 4969 31946 4978
rect 33334 5012 33386 5021
rect 33334 4978 33343 5012
rect 33343 4978 33377 5012
rect 33377 4978 33386 5012
rect 33334 4969 33386 4978
rect 33430 4969 33482 5021
rect 34870 5012 34922 5021
rect 34870 4978 34879 5012
rect 34879 4978 34913 5012
rect 34913 4978 34922 5012
rect 34870 4969 34922 4978
rect 35638 5012 35690 5021
rect 35638 4978 35647 5012
rect 35647 4978 35681 5012
rect 35681 4978 35690 5012
rect 35638 4969 35690 4978
rect 36118 4969 36170 5021
rect 36886 4969 36938 5021
rect 38614 5012 38666 5021
rect 38614 4978 38623 5012
rect 38623 4978 38657 5012
rect 38657 4978 38666 5012
rect 38614 4969 38666 4978
rect 39382 5012 39434 5021
rect 39382 4978 39391 5012
rect 39391 4978 39425 5012
rect 39425 4978 39434 5012
rect 39382 4969 39434 4978
rect 40150 5012 40202 5021
rect 40150 4978 40159 5012
rect 40159 4978 40193 5012
rect 40193 4978 40202 5012
rect 40150 4969 40202 4978
rect 40918 5012 40970 5021
rect 40918 4978 40927 5012
rect 40927 4978 40961 5012
rect 40961 4978 40970 5012
rect 40918 4969 40970 4978
rect 41302 4969 41354 5021
rect 42454 5012 42506 5021
rect 42454 4978 42463 5012
rect 42463 4978 42497 5012
rect 42497 4978 42506 5012
rect 42454 4969 42506 4978
rect 43894 5012 43946 5021
rect 43894 4978 43903 5012
rect 43903 4978 43937 5012
rect 43937 4978 43946 5012
rect 43894 4969 43946 4978
rect 43990 4969 44042 5021
rect 44854 4969 44906 5021
rect 45622 4969 45674 5021
rect 46486 4969 46538 5021
rect 47926 4969 47978 5021
rect 49366 5012 49418 5021
rect 49366 4978 49375 5012
rect 49375 4978 49409 5012
rect 49409 4978 49418 5012
rect 49366 4969 49418 4978
rect 50422 5012 50474 5021
rect 50422 4978 50431 5012
rect 50431 4978 50465 5012
rect 50465 4978 50474 5012
rect 50422 4969 50474 4978
rect 50902 4969 50954 5021
rect 51862 5012 51914 5021
rect 51862 4978 51871 5012
rect 51871 4978 51905 5012
rect 51905 4978 51914 5012
rect 51862 4969 51914 4978
rect 51958 4969 52010 5021
rect 53302 4969 53354 5021
rect 59254 5117 59306 5169
rect 57814 5043 57866 5095
rect 57046 5012 57098 5021
rect 57046 4978 57055 5012
rect 57055 4978 57089 5012
rect 57089 4978 57098 5012
rect 57046 4969 57098 4978
rect 8566 4821 8618 4873
rect 26422 4821 26474 4873
rect 15766 4747 15818 4799
rect 37846 4747 37898 4799
rect 19654 4636 19706 4688
rect 19718 4636 19770 4688
rect 19782 4636 19834 4688
rect 19846 4636 19898 4688
rect 50374 4636 50426 4688
rect 50438 4636 50490 4688
rect 50502 4636 50554 4688
rect 50566 4636 50618 4688
rect 15766 4568 15818 4577
rect 15766 4534 15775 4568
rect 15775 4534 15809 4568
rect 15809 4534 15818 4568
rect 15766 4525 15818 4534
rect 19126 4568 19178 4577
rect 19126 4534 19135 4568
rect 19135 4534 19169 4568
rect 19169 4534 19178 4568
rect 19126 4525 19178 4534
rect 23926 4525 23978 4577
rect 24406 4525 24458 4577
rect 34198 4525 34250 4577
rect 790 4377 842 4429
rect 1174 4303 1226 4355
rect 1366 4229 1418 4281
rect 3766 4229 3818 4281
rect 4726 4451 4778 4503
rect 42934 4451 42986 4503
rect 43030 4377 43082 4429
rect 4726 4303 4778 4355
rect 5014 4229 5066 4281
rect 7414 4346 7466 4355
rect 5686 4229 5738 4281
rect 7414 4312 7423 4346
rect 7423 4312 7457 4346
rect 7457 4312 7466 4346
rect 7414 4303 7466 4312
rect 9622 4346 9674 4355
rect 6166 4155 6218 4207
rect 6454 4155 6506 4207
rect 9622 4312 9631 4346
rect 9631 4312 9665 4346
rect 9665 4312 9674 4346
rect 9622 4303 9674 4312
rect 10390 4346 10442 4355
rect 10390 4312 10399 4346
rect 10399 4312 10433 4346
rect 10433 4312 10442 4346
rect 10390 4303 10442 4312
rect 10774 4303 10826 4355
rect 13558 4346 13610 4355
rect 11158 4155 11210 4207
rect 11446 4081 11498 4133
rect 13558 4312 13567 4346
rect 13567 4312 13601 4346
rect 13601 4312 13610 4346
rect 13558 4303 13610 4312
rect 15478 4346 15530 4355
rect 15478 4312 15487 4346
rect 15487 4312 15521 4346
rect 15521 4312 15530 4346
rect 15478 4303 15530 4312
rect 15958 4303 16010 4355
rect 18838 4346 18890 4355
rect 16246 4155 16298 4207
rect 18838 4312 18847 4346
rect 18847 4312 18881 4346
rect 18881 4312 18890 4346
rect 18838 4303 18890 4312
rect 21046 4346 21098 4355
rect 16918 4081 16970 4133
rect 19510 4229 19562 4281
rect 21046 4312 21055 4346
rect 21055 4312 21089 4346
rect 21089 4312 21098 4346
rect 21046 4303 21098 4312
rect 21814 4346 21866 4355
rect 21814 4312 21823 4346
rect 21823 4312 21857 4346
rect 21857 4312 21866 4346
rect 21814 4303 21866 4312
rect 23254 4346 23306 4355
rect 23254 4312 23263 4346
rect 23263 4312 23297 4346
rect 23297 4312 23306 4346
rect 23254 4303 23306 4312
rect 24022 4346 24074 4355
rect 24022 4312 24031 4346
rect 24031 4312 24065 4346
rect 24065 4312 24074 4346
rect 24022 4303 24074 4312
rect 25462 4346 25514 4355
rect 25462 4312 25471 4346
rect 25471 4312 25505 4346
rect 25505 4312 25514 4346
rect 25462 4303 25514 4312
rect 26134 4303 26186 4355
rect 26518 4303 26570 4355
rect 28342 4346 28394 4355
rect 28342 4312 28351 4346
rect 28351 4312 28385 4346
rect 28385 4312 28394 4346
rect 28342 4303 28394 4312
rect 29110 4346 29162 4355
rect 29110 4312 29119 4346
rect 29119 4312 29153 4346
rect 29153 4312 29162 4346
rect 29110 4303 29162 4312
rect 30934 4346 30986 4355
rect 30934 4312 30943 4346
rect 30943 4312 30977 4346
rect 30977 4312 30986 4346
rect 30934 4303 30986 4312
rect 31702 4346 31754 4355
rect 31702 4312 31711 4346
rect 31711 4312 31745 4346
rect 31745 4312 31754 4346
rect 31702 4303 31754 4312
rect 32758 4346 32810 4355
rect 32758 4312 32767 4346
rect 32767 4312 32801 4346
rect 32801 4312 32810 4346
rect 32758 4303 32810 4312
rect 33910 4346 33962 4355
rect 33910 4312 33919 4346
rect 33919 4312 33953 4346
rect 33953 4312 33962 4346
rect 33910 4303 33962 4312
rect 34582 4303 34634 4355
rect 20950 4229 21002 4281
rect 21718 4229 21770 4281
rect 28054 4229 28106 4281
rect 28534 4229 28586 4281
rect 29398 4229 29450 4281
rect 20086 4155 20138 4207
rect 21430 4155 21482 4207
rect 21526 4155 21578 4207
rect 22870 4155 22922 4207
rect 24118 4155 24170 4207
rect 24502 4155 24554 4207
rect 25558 4155 25610 4207
rect 25942 4155 25994 4207
rect 26998 4155 27050 4207
rect 27382 4155 27434 4207
rect 28246 4155 28298 4207
rect 29014 4155 29066 4207
rect 18262 4081 18314 4133
rect 34198 4229 34250 4281
rect 36790 4346 36842 4355
rect 36790 4312 36799 4346
rect 36799 4312 36833 4346
rect 36833 4312 36842 4346
rect 36790 4303 36842 4312
rect 38998 4346 39050 4355
rect 37174 4229 37226 4281
rect 38998 4312 39007 4346
rect 39007 4312 39041 4346
rect 39041 4312 39050 4346
rect 38998 4303 39050 4312
rect 39766 4346 39818 4355
rect 39766 4312 39775 4346
rect 39775 4312 39809 4346
rect 39809 4312 39818 4346
rect 39766 4303 39818 4312
rect 41974 4346 42026 4355
rect 41974 4312 41983 4346
rect 41983 4312 42017 4346
rect 42017 4312 42026 4346
rect 41974 4303 42026 4312
rect 42262 4303 42314 4355
rect 43414 4303 43466 4355
rect 44950 4346 45002 4355
rect 44950 4312 44959 4346
rect 44959 4312 44993 4346
rect 44993 4312 45002 4346
rect 44950 4303 45002 4312
rect 46774 4346 46826 4355
rect 46774 4312 46783 4346
rect 46783 4312 46817 4346
rect 46817 4312 46826 4346
rect 46774 4303 46826 4312
rect 41398 4229 41450 4281
rect 41590 4229 41642 4281
rect 42070 4229 42122 4281
rect 43126 4229 43178 4281
rect 44086 4229 44138 4281
rect 44662 4229 44714 4281
rect 47446 4229 47498 4281
rect 47830 4303 47882 4355
rect 48598 4229 48650 4281
rect 49174 4303 49226 4355
rect 52630 4346 52682 4355
rect 48118 4155 48170 4207
rect 48982 4155 49034 4207
rect 49846 4155 49898 4207
rect 50998 4229 51050 4281
rect 52630 4312 52639 4346
rect 52639 4312 52673 4346
rect 52673 4312 52682 4346
rect 52630 4303 52682 4312
rect 53014 4229 53066 4281
rect 54070 4303 54122 4355
rect 55606 4346 55658 4355
rect 55606 4312 55615 4346
rect 55615 4312 55649 4346
rect 55649 4312 55658 4346
rect 55606 4303 55658 4312
rect 56662 4303 56714 4355
rect 54838 4229 54890 4281
rect 57142 4155 57194 4207
rect 58294 4229 58346 4281
rect 33814 4081 33866 4133
rect 34678 4081 34730 4133
rect 36694 4081 36746 4133
rect 37558 4081 37610 4133
rect 38518 4081 38570 4133
rect 40150 4081 40202 4133
rect 43798 4081 43850 4133
rect 47158 4081 47210 4133
rect 48502 4081 48554 4133
rect 49654 4081 49706 4133
rect 56566 4081 56618 4133
rect 59158 4081 59210 4133
rect 4294 3970 4346 4022
rect 4358 3970 4410 4022
rect 4422 3970 4474 4022
rect 4486 3970 4538 4022
rect 35014 3970 35066 4022
rect 35078 3970 35130 4022
rect 35142 3970 35194 4022
rect 35206 3970 35258 4022
rect 1942 3859 1994 3911
rect 3382 3859 3434 3911
rect 8758 3859 8810 3911
rect 10294 3859 10346 3911
rect 15382 3859 15434 3911
rect 16438 3859 16490 3911
rect 18358 3859 18410 3911
rect 19030 3859 19082 3911
rect 21334 3859 21386 3911
rect 22774 3859 22826 3911
rect 24502 3859 24554 3911
rect 24886 3859 24938 3911
rect 25366 3859 25418 3911
rect 26230 3859 26282 3911
rect 27478 3859 27530 3911
rect 28918 3859 28970 3911
rect 29014 3859 29066 3911
rect 30358 3859 30410 3911
rect 34486 3859 34538 3911
rect 35638 3859 35690 3911
rect 38134 3859 38186 3911
rect 39094 3859 39146 3911
rect 39670 3859 39722 3911
rect 40918 3859 40970 3911
rect 41206 3859 41258 3911
rect 502 3785 554 3837
rect 1654 3785 1706 3837
rect 2326 3785 2378 3837
rect 3094 3785 3146 3837
rect 8278 3785 8330 3837
rect 9238 3785 9290 3837
rect 12022 3785 12074 3837
rect 13366 3785 13418 3837
rect 13654 3785 13706 3837
rect 18262 3785 18314 3837
rect 22390 3785 22442 3837
rect 24214 3785 24266 3837
rect 25846 3785 25898 3837
rect 25942 3785 25994 3837
rect 27094 3785 27146 3837
rect 28054 3785 28106 3837
rect 35446 3785 35498 3837
rect 36022 3785 36074 3837
rect 36406 3785 36458 3837
rect 37078 3785 37130 3837
rect 38614 3785 38666 3837
rect 42550 3785 42602 3837
rect 43510 3785 43562 3837
rect 43702 3859 43754 3911
rect 44854 3859 44906 3911
rect 46294 3859 46346 3911
rect 47926 3859 47978 3911
rect 49270 3859 49322 3911
rect 50710 3859 50762 3911
rect 51382 3859 51434 3911
rect 51862 3859 51914 3911
rect 55990 3859 56042 3911
rect 43798 3785 43850 3837
rect 44470 3785 44522 3837
rect 45622 3785 45674 3837
rect 56758 3785 56810 3837
rect 57142 3785 57194 3837
rect 57910 3785 57962 3837
rect 982 3711 1034 3763
rect 2422 3711 2474 3763
rect 3382 3711 3434 3763
rect 118 3637 170 3689
rect 1654 3637 1706 3689
rect 2710 3637 2762 3689
rect 10294 3711 10346 3763
rect 11062 3711 11114 3763
rect 14230 3711 14282 3763
rect 14422 3711 14474 3763
rect 17782 3711 17834 3763
rect 18550 3754 18602 3763
rect 18550 3720 18559 3754
rect 18559 3720 18593 3754
rect 18593 3720 18602 3754
rect 18550 3711 18602 3720
rect 19414 3711 19466 3763
rect 20566 3711 20618 3763
rect 22102 3711 22154 3763
rect 24022 3711 24074 3763
rect 26326 3711 26378 3763
rect 27574 3711 27626 3763
rect 28726 3711 28778 3763
rect 5590 3680 5642 3689
rect 214 3563 266 3615
rect 1750 3563 1802 3615
rect 3094 3489 3146 3541
rect 5590 3646 5599 3680
rect 5599 3646 5633 3680
rect 5633 3646 5642 3680
rect 5590 3637 5642 3646
rect 6358 3637 6410 3689
rect 7030 3637 7082 3689
rect 7798 3637 7850 3689
rect 8566 3637 8618 3689
rect 9334 3637 9386 3689
rect 10006 3489 10058 3541
rect 13174 3637 13226 3689
rect 13366 3637 13418 3689
rect 13654 3563 13706 3615
rect 15190 3637 15242 3689
rect 17398 3637 17450 3689
rect 18262 3637 18314 3689
rect 18454 3563 18506 3615
rect 20278 3637 20330 3689
rect 20566 3563 20618 3615
rect 22678 3637 22730 3689
rect 22870 3637 22922 3689
rect 23638 3637 23690 3689
rect 24406 3637 24458 3689
rect 22966 3563 23018 3615
rect 24694 3563 24746 3615
rect 21718 3489 21770 3541
rect 22582 3489 22634 3541
rect 23542 3489 23594 3541
rect 24310 3489 24362 3541
rect 25846 3489 25898 3541
rect 27286 3637 27338 3689
rect 32662 3711 32714 3763
rect 33430 3711 33482 3763
rect 45238 3711 45290 3763
rect 28054 3489 28106 3541
rect 29494 3563 29546 3615
rect 30454 3637 30506 3689
rect 31318 3637 31370 3689
rect 32470 3637 32522 3689
rect 33526 3637 33578 3689
rect 34294 3637 34346 3689
rect 34966 3637 35018 3689
rect 35734 3637 35786 3689
rect 36502 3637 36554 3689
rect 37942 3637 37994 3689
rect 38710 3637 38762 3689
rect 39478 3637 39530 3689
rect 40246 3637 40298 3689
rect 41014 3637 41066 3689
rect 35350 3563 35402 3615
rect 36214 3563 36266 3615
rect 40054 3563 40106 3615
rect 41302 3563 41354 3615
rect 41590 3563 41642 3615
rect 42742 3637 42794 3689
rect 55894 3711 55946 3763
rect 43798 3563 43850 3615
rect 30454 3489 30506 3541
rect 31894 3489 31946 3541
rect 37846 3489 37898 3541
rect 39382 3489 39434 3541
rect 44566 3489 44618 3541
rect 46006 3563 46058 3615
rect 47158 3637 47210 3689
rect 48214 3637 48266 3689
rect 50710 3637 50762 3689
rect 50806 3637 50858 3689
rect 49078 3489 49130 3541
rect 50038 3489 50090 3541
rect 51190 3489 51242 3541
rect 52054 3637 52106 3689
rect 53398 3637 53450 3689
rect 54358 3563 54410 3615
rect 52054 3489 52106 3541
rect 52822 3489 52874 3541
rect 55222 3489 55274 3541
rect 56278 3563 56330 3615
rect 58198 3637 58250 3689
rect 59734 3637 59786 3689
rect 56374 3489 56426 3541
rect 56758 3489 56810 3541
rect 3958 3415 4010 3467
rect 5110 3415 5162 3467
rect 14038 3415 14090 3467
rect 19894 3415 19946 3467
rect 20182 3415 20234 3467
rect 23062 3415 23114 3467
rect 23830 3415 23882 3467
rect 24982 3415 25034 3467
rect 26614 3415 26666 3467
rect 27382 3415 27434 3467
rect 29302 3415 29354 3467
rect 29398 3415 29450 3467
rect 31126 3415 31178 3467
rect 33430 3415 33482 3467
rect 34870 3415 34922 3467
rect 56566 3415 56618 3467
rect 57334 3415 57386 3467
rect 19654 3304 19706 3356
rect 19718 3304 19770 3356
rect 19782 3304 19834 3356
rect 19846 3304 19898 3356
rect 50374 3304 50426 3356
rect 50438 3304 50490 3356
rect 50502 3304 50554 3356
rect 50566 3304 50618 3356
rect 598 3193 650 3245
rect 1462 3193 1514 3245
rect 2422 3193 2474 3245
rect 5206 3193 5258 3245
rect 9430 3193 9482 3245
rect 10678 3193 10730 3245
rect 12214 3193 12266 3245
rect 12982 3193 13034 3245
rect 19702 3193 19754 3245
rect 20374 3193 20426 3245
rect 21622 3236 21674 3245
rect 21622 3202 21631 3236
rect 21631 3202 21665 3236
rect 21665 3202 21674 3236
rect 21622 3193 21674 3202
rect 21718 3193 21770 3245
rect 41206 3193 41258 3245
rect 42166 3193 42218 3245
rect 43894 3193 43946 3245
rect 45142 3193 45194 3245
rect 46486 3193 46538 3245
rect 56854 3193 56906 3245
rect 58006 3193 58058 3245
rect 3478 3119 3530 3171
rect 4918 3119 4970 3171
rect 5110 3119 5162 3171
rect 5974 3119 6026 3171
rect 6166 3119 6218 3171
rect 1462 3045 1514 3097
rect 2134 3045 2186 3097
rect 6838 3045 6890 3097
rect 7702 3045 7754 3097
rect 8950 3045 9002 3097
rect 22 2971 74 3023
rect 694 2897 746 2949
rect 4918 3014 4970 3023
rect 2134 2897 2186 2949
rect 4918 2980 4927 3014
rect 4927 2980 4961 3014
rect 4961 2980 4970 3014
rect 4918 2971 4970 2980
rect 5206 2971 5258 3023
rect 5974 2971 6026 3023
rect 6742 2897 6794 2949
rect 8182 2971 8234 3023
rect 7702 2897 7754 2949
rect 7990 2897 8042 2949
rect 9814 2897 9866 2949
rect 10198 2897 10250 2949
rect 11542 2897 11594 2949
rect 22390 3119 22442 3171
rect 23158 3119 23210 3171
rect 18934 3045 18986 3097
rect 13078 2971 13130 3023
rect 14038 2971 14090 3023
rect 14806 2971 14858 3023
rect 16630 3014 16682 3023
rect 16630 2980 16639 3014
rect 16639 2980 16673 3014
rect 16673 2980 16682 3014
rect 16630 2971 16682 2980
rect 17014 2971 17066 3023
rect 13750 2897 13802 2949
rect 17782 2897 17834 2949
rect 17686 2823 17738 2875
rect 18934 2823 18986 2875
rect 19318 2897 19370 2949
rect 19318 2749 19370 2801
rect 21622 3045 21674 3097
rect 22486 3045 22538 3097
rect 31894 3045 31946 3097
rect 33334 3045 33386 3097
rect 42454 3045 42506 3097
rect 42934 3045 42986 3097
rect 43990 3045 44042 3097
rect 44374 3045 44426 3097
rect 45334 3045 45386 3097
rect 20662 2940 20714 2949
rect 20662 2906 20671 2940
rect 20671 2906 20705 2940
rect 20705 2906 20714 2940
rect 20662 2897 20714 2906
rect 21430 2897 21482 2949
rect 22486 2897 22538 2949
rect 24022 2971 24074 3023
rect 25078 2897 25130 2949
rect 26902 2971 26954 3023
rect 27670 2897 27722 2949
rect 29878 2971 29930 3023
rect 28918 2823 28970 2875
rect 29782 2897 29834 2949
rect 30550 2897 30602 2949
rect 32086 2971 32138 3023
rect 32278 2897 32330 2949
rect 33142 2897 33194 2949
rect 33334 2897 33386 2949
rect 35446 2971 35498 3023
rect 36214 2897 36266 2949
rect 37558 2971 37610 3023
rect 38326 2897 38378 2949
rect 40534 2971 40586 3023
rect 41110 2940 41162 2949
rect 41110 2906 41119 2940
rect 41119 2906 41153 2940
rect 41153 2906 41162 2940
rect 41110 2897 41162 2906
rect 41206 2897 41258 2949
rect 43030 2971 43082 3023
rect 43894 2897 43946 2949
rect 44182 2897 44234 2949
rect 45622 2971 45674 3023
rect 46390 2897 46442 2949
rect 49654 2971 49706 3023
rect 49942 2897 49994 2949
rect 51478 2971 51530 3023
rect 52246 2897 52298 2949
rect 53782 2971 53834 3023
rect 52918 2897 52970 2949
rect 53686 2897 53738 2949
rect 54838 2897 54890 2949
rect 57718 2897 57770 2949
rect 59446 2897 59498 2949
rect 35638 2823 35690 2875
rect 36886 2823 36938 2875
rect 37270 2823 37322 2875
rect 19894 2749 19946 2801
rect 24886 2792 24938 2801
rect 24886 2758 24895 2792
rect 24895 2758 24929 2792
rect 24929 2758 24938 2792
rect 24886 2749 24938 2758
rect 35254 2749 35306 2801
rect 42454 2749 42506 2801
rect 44662 2749 44714 2801
rect 45046 2749 45098 2801
rect 54454 2792 54506 2801
rect 54454 2758 54463 2792
rect 54463 2758 54497 2792
rect 54497 2758 54506 2792
rect 54454 2749 54506 2758
rect 4294 2638 4346 2690
rect 4358 2638 4410 2690
rect 4422 2638 4474 2690
rect 4486 2638 4538 2690
rect 35014 2638 35066 2690
rect 35078 2638 35130 2690
rect 35142 2638 35194 2690
rect 35206 2638 35258 2690
rect 3958 2527 4010 2579
rect 4246 2527 4298 2579
rect 4342 2527 4394 2579
rect 4822 2527 4874 2579
rect 20182 2527 20234 2579
rect 21238 2527 21290 2579
rect 35158 2527 35210 2579
rect 35542 2527 35594 2579
rect 42454 2527 42506 2579
rect 54454 2527 54506 2579
rect 24886 2453 24938 2505
rect 52822 2453 52874 2505
rect 34102 2379 34154 2431
rect 37270 2379 37322 2431
rect 45046 2379 45098 2431
rect 45814 2379 45866 2431
rect 4726 2009 4778 2061
rect 5302 2009 5354 2061
rect 4534 1861 4586 1913
rect 4822 1861 4874 1913
rect 18070 1861 18122 1913
rect 18262 1861 18314 1913
rect 13078 1713 13130 1765
rect 13270 1713 13322 1765
rect 30358 1713 30410 1765
rect 30646 1713 30698 1765
rect 34870 1713 34922 1765
rect 35926 1713 35978 1765
rect 39958 1713 40010 1765
rect 40246 1713 40298 1765
rect 50710 1713 50762 1765
rect 50902 1713 50954 1765
rect 54358 1713 54410 1765
rect 54646 1713 54698 1765
rect 50518 1639 50570 1691
rect 51094 1639 51146 1691
rect 20470 1565 20522 1617
rect 20854 1565 20906 1617
rect 22102 1565 22154 1617
rect 22678 1565 22730 1617
rect 50902 1565 50954 1617
rect 51574 1565 51626 1617
rect 36310 1491 36362 1543
rect 19318 1417 19370 1469
rect 19990 1417 20042 1469
rect 33238 1417 33290 1469
rect 33718 1417 33770 1469
rect 36310 1121 36362 1173
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 226 56975 254 59200
rect 214 56969 266 56975
rect 214 56911 266 56917
rect 706 56531 734 59200
rect 694 56525 746 56531
rect 694 56467 746 56473
rect 1186 55717 1214 59200
rect 1762 56975 1790 59200
rect 1750 56969 1802 56975
rect 1750 56911 1802 56917
rect 1750 56229 1802 56235
rect 1750 56171 1802 56177
rect 1174 55711 1226 55717
rect 1174 55653 1226 55659
rect 1762 30927 1790 56171
rect 2242 56161 2270 59200
rect 2818 56531 2846 59200
rect 3298 56975 3326 59200
rect 3286 56969 3338 56975
rect 3286 56911 3338 56917
rect 3874 56531 3902 59200
rect 4354 57614 4382 59200
rect 4354 57586 4670 57614
rect 4268 57304 4564 57324
rect 4324 57302 4348 57304
rect 4404 57302 4428 57304
rect 4484 57302 4508 57304
rect 4346 57250 4348 57302
rect 4410 57250 4422 57302
rect 4484 57250 4486 57302
rect 4324 57248 4348 57250
rect 4404 57248 4428 57250
rect 4484 57248 4508 57250
rect 4268 57228 4564 57248
rect 2806 56525 2858 56531
rect 2806 56467 2858 56473
rect 3862 56525 3914 56531
rect 3862 56467 3914 56473
rect 2998 56229 3050 56235
rect 2998 56171 3050 56177
rect 2230 56155 2282 56161
rect 2230 56097 2282 56103
rect 2038 55415 2090 55421
rect 2038 55357 2090 55363
rect 2050 55051 2078 55357
rect 2038 55045 2090 55051
rect 2038 54987 2090 54993
rect 2134 52085 2186 52091
rect 2134 52027 2186 52033
rect 1942 36101 1994 36107
rect 1942 36043 1994 36049
rect 1750 30921 1802 30927
rect 1750 30863 1802 30869
rect 1954 23749 1982 36043
rect 1942 23743 1994 23749
rect 1942 23685 1994 23691
rect 2146 8579 2174 52027
rect 3010 30409 3038 56171
rect 4268 55972 4564 55992
rect 4324 55970 4348 55972
rect 4404 55970 4428 55972
rect 4484 55970 4508 55972
rect 4346 55918 4348 55970
rect 4410 55918 4422 55970
rect 4484 55918 4486 55970
rect 4324 55916 4348 55918
rect 4404 55916 4428 55918
rect 4484 55916 4508 55918
rect 4268 55896 4564 55916
rect 4642 55717 4670 57586
rect 4930 56975 4958 59200
rect 4918 56969 4970 56975
rect 4918 56911 4970 56917
rect 4822 56747 4874 56753
rect 4822 56689 4874 56695
rect 5206 56747 5258 56753
rect 5206 56689 5258 56695
rect 4726 56229 4778 56235
rect 4726 56171 4778 56177
rect 4630 55711 4682 55717
rect 4630 55653 4682 55659
rect 4268 54640 4564 54660
rect 4324 54638 4348 54640
rect 4404 54638 4428 54640
rect 4484 54638 4508 54640
rect 4346 54586 4348 54638
rect 4410 54586 4422 54638
rect 4484 54586 4486 54638
rect 4324 54584 4348 54586
rect 4404 54584 4428 54586
rect 4484 54584 4508 54586
rect 4268 54564 4564 54584
rect 4268 53308 4564 53328
rect 4324 53306 4348 53308
rect 4404 53306 4428 53308
rect 4484 53306 4508 53308
rect 4346 53254 4348 53306
rect 4410 53254 4422 53306
rect 4484 53254 4486 53306
rect 4324 53252 4348 53254
rect 4404 53252 4428 53254
rect 4484 53252 4508 53254
rect 4268 53232 4564 53252
rect 4268 51976 4564 51996
rect 4324 51974 4348 51976
rect 4404 51974 4428 51976
rect 4484 51974 4508 51976
rect 4346 51922 4348 51974
rect 4410 51922 4422 51974
rect 4484 51922 4486 51974
rect 4324 51920 4348 51922
rect 4404 51920 4428 51922
rect 4484 51920 4508 51922
rect 4268 51900 4564 51920
rect 4268 50644 4564 50664
rect 4324 50642 4348 50644
rect 4404 50642 4428 50644
rect 4484 50642 4508 50644
rect 4346 50590 4348 50642
rect 4410 50590 4422 50642
rect 4484 50590 4486 50642
rect 4324 50588 4348 50590
rect 4404 50588 4428 50590
rect 4484 50588 4508 50590
rect 4268 50568 4564 50588
rect 4268 49312 4564 49332
rect 4324 49310 4348 49312
rect 4404 49310 4428 49312
rect 4484 49310 4508 49312
rect 4346 49258 4348 49310
rect 4410 49258 4422 49310
rect 4484 49258 4486 49310
rect 4324 49256 4348 49258
rect 4404 49256 4428 49258
rect 4484 49256 4508 49258
rect 4268 49236 4564 49256
rect 4268 47980 4564 48000
rect 4324 47978 4348 47980
rect 4404 47978 4428 47980
rect 4484 47978 4508 47980
rect 4346 47926 4348 47978
rect 4410 47926 4422 47978
rect 4484 47926 4486 47978
rect 4324 47924 4348 47926
rect 4404 47924 4428 47926
rect 4484 47924 4508 47926
rect 4268 47904 4564 47924
rect 4738 47534 4766 56171
rect 4834 48465 4862 56689
rect 4822 48459 4874 48465
rect 4822 48401 4874 48407
rect 4642 47506 4766 47534
rect 4268 46648 4564 46668
rect 4324 46646 4348 46648
rect 4404 46646 4428 46648
rect 4484 46646 4508 46648
rect 4346 46594 4348 46646
rect 4410 46594 4422 46646
rect 4484 46594 4486 46646
rect 4324 46592 4348 46594
rect 4404 46592 4428 46594
rect 4484 46592 4508 46594
rect 4268 46572 4564 46592
rect 4268 45316 4564 45336
rect 4324 45314 4348 45316
rect 4404 45314 4428 45316
rect 4484 45314 4508 45316
rect 4346 45262 4348 45314
rect 4410 45262 4422 45314
rect 4484 45262 4486 45314
rect 4324 45260 4348 45262
rect 4404 45260 4428 45262
rect 4484 45260 4508 45262
rect 4268 45240 4564 45260
rect 4268 43984 4564 44004
rect 4324 43982 4348 43984
rect 4404 43982 4428 43984
rect 4484 43982 4508 43984
rect 4346 43930 4348 43982
rect 4410 43930 4422 43982
rect 4484 43930 4486 43982
rect 4324 43928 4348 43930
rect 4404 43928 4428 43930
rect 4484 43928 4508 43930
rect 4268 43908 4564 43928
rect 4268 42652 4564 42672
rect 4324 42650 4348 42652
rect 4404 42650 4428 42652
rect 4484 42650 4508 42652
rect 4346 42598 4348 42650
rect 4410 42598 4422 42650
rect 4484 42598 4486 42650
rect 4324 42596 4348 42598
rect 4404 42596 4428 42598
rect 4484 42596 4508 42598
rect 4268 42576 4564 42596
rect 4268 41320 4564 41340
rect 4324 41318 4348 41320
rect 4404 41318 4428 41320
rect 4484 41318 4508 41320
rect 4346 41266 4348 41318
rect 4410 41266 4422 41318
rect 4484 41266 4486 41318
rect 4324 41264 4348 41266
rect 4404 41264 4428 41266
rect 4484 41264 4508 41266
rect 4268 41244 4564 41264
rect 4268 39988 4564 40008
rect 4324 39986 4348 39988
rect 4404 39986 4428 39988
rect 4484 39986 4508 39988
rect 4346 39934 4348 39986
rect 4410 39934 4422 39986
rect 4484 39934 4486 39986
rect 4324 39932 4348 39934
rect 4404 39932 4428 39934
rect 4484 39932 4508 39934
rect 4268 39912 4564 39932
rect 4268 38656 4564 38676
rect 4324 38654 4348 38656
rect 4404 38654 4428 38656
rect 4484 38654 4508 38656
rect 4346 38602 4348 38654
rect 4410 38602 4422 38654
rect 4484 38602 4486 38654
rect 4324 38600 4348 38602
rect 4404 38600 4428 38602
rect 4484 38600 4508 38602
rect 4268 38580 4564 38600
rect 4268 37324 4564 37344
rect 4324 37322 4348 37324
rect 4404 37322 4428 37324
rect 4484 37322 4508 37324
rect 4346 37270 4348 37322
rect 4410 37270 4422 37322
rect 4484 37270 4486 37322
rect 4324 37268 4348 37270
rect 4404 37268 4428 37270
rect 4484 37268 4508 37270
rect 4268 37248 4564 37268
rect 4268 35992 4564 36012
rect 4324 35990 4348 35992
rect 4404 35990 4428 35992
rect 4484 35990 4508 35992
rect 4346 35938 4348 35990
rect 4410 35938 4422 35990
rect 4484 35938 4486 35990
rect 4324 35936 4348 35938
rect 4404 35936 4428 35938
rect 4484 35936 4508 35938
rect 4268 35916 4564 35936
rect 4534 35657 4586 35663
rect 4534 35599 4586 35605
rect 4546 35071 4574 35599
rect 4534 35065 4586 35071
rect 4534 35007 4586 35013
rect 4268 34660 4564 34680
rect 4324 34658 4348 34660
rect 4404 34658 4428 34660
rect 4484 34658 4508 34660
rect 4346 34606 4348 34658
rect 4410 34606 4422 34658
rect 4484 34606 4486 34658
rect 4324 34604 4348 34606
rect 4404 34604 4428 34606
rect 4484 34604 4508 34606
rect 4268 34584 4564 34604
rect 4268 33328 4564 33348
rect 4324 33326 4348 33328
rect 4404 33326 4428 33328
rect 4484 33326 4508 33328
rect 4346 33274 4348 33326
rect 4410 33274 4422 33326
rect 4484 33274 4486 33326
rect 4324 33272 4348 33274
rect 4404 33272 4428 33274
rect 4484 33272 4508 33274
rect 4268 33252 4564 33272
rect 4268 31996 4564 32016
rect 4324 31994 4348 31996
rect 4404 31994 4428 31996
rect 4484 31994 4508 31996
rect 4346 31942 4348 31994
rect 4410 31942 4422 31994
rect 4484 31942 4486 31994
rect 4324 31940 4348 31942
rect 4404 31940 4428 31942
rect 4484 31940 4508 31942
rect 4268 31920 4564 31940
rect 4268 30664 4564 30684
rect 4324 30662 4348 30664
rect 4404 30662 4428 30664
rect 4484 30662 4508 30664
rect 4346 30610 4348 30662
rect 4410 30610 4422 30662
rect 4484 30610 4486 30662
rect 4324 30608 4348 30610
rect 4404 30608 4428 30610
rect 4484 30608 4508 30610
rect 4268 30588 4564 30608
rect 2998 30403 3050 30409
rect 2998 30345 3050 30351
rect 3574 29515 3626 29521
rect 3574 29457 3626 29463
rect 2134 8573 2186 8579
rect 2134 8515 2186 8521
rect 1654 8277 1706 8283
rect 1654 8219 1706 8225
rect 2134 8277 2186 8283
rect 2134 8219 2186 8225
rect 2998 8277 3050 8283
rect 2998 8219 3050 8225
rect 1462 7685 1514 7691
rect 1462 7627 1514 7633
rect 1078 5687 1130 5693
rect 1078 5629 1130 5635
rect 310 5021 362 5027
rect 310 4963 362 4969
rect 118 3689 170 3695
rect 118 3631 170 3637
rect 22 3023 74 3029
rect 22 2965 74 2971
rect 34 800 62 2965
rect 130 800 158 3631
rect 214 3615 266 3621
rect 214 3557 266 3563
rect 226 800 254 3557
rect 322 800 350 4963
rect 790 4429 842 4435
rect 790 4371 842 4377
rect 502 3837 554 3843
rect 502 3779 554 3785
rect 514 800 542 3779
rect 598 3245 650 3251
rect 598 3187 650 3193
rect 610 800 638 3187
rect 694 2949 746 2955
rect 694 2891 746 2897
rect 706 800 734 2891
rect 802 800 830 4371
rect 982 3763 1034 3769
rect 982 3705 1034 3711
rect 994 800 1022 3705
rect 1090 800 1118 5629
rect 1174 4355 1226 4361
rect 1174 4297 1226 4303
rect 1186 800 1214 4297
rect 1366 4281 1418 4287
rect 1366 4223 1418 4229
rect 1378 800 1406 4223
rect 1474 3251 1502 7627
rect 1666 7214 1694 8219
rect 1666 7186 1790 7214
rect 1654 7019 1706 7025
rect 1654 6961 1706 6967
rect 1558 6353 1610 6359
rect 1558 6295 1610 6301
rect 1462 3245 1514 3251
rect 1462 3187 1514 3193
rect 1462 3097 1514 3103
rect 1462 3039 1514 3045
rect 1474 800 1502 3039
rect 1570 800 1598 6295
rect 1666 3843 1694 6961
rect 1654 3837 1706 3843
rect 1654 3779 1706 3785
rect 1654 3689 1706 3695
rect 1654 3631 1706 3637
rect 1666 800 1694 3631
rect 1762 3621 1790 7186
rect 2038 6353 2090 6359
rect 2038 6295 2090 6301
rect 1846 5021 1898 5027
rect 1846 4963 1898 4969
rect 1750 3615 1802 3621
rect 1750 3557 1802 3563
rect 1858 800 1886 4963
rect 1942 3911 1994 3917
rect 1942 3853 1994 3859
rect 1954 800 1982 3853
rect 2050 800 2078 6295
rect 2146 3103 2174 8219
rect 2422 7463 2474 7469
rect 2422 7405 2474 7411
rect 2326 3837 2378 3843
rect 2326 3779 2378 3785
rect 2134 3097 2186 3103
rect 2134 3039 2186 3045
rect 2134 2949 2186 2955
rect 2134 2891 2186 2897
rect 2146 800 2174 2891
rect 2338 800 2366 3779
rect 2434 3769 2462 7405
rect 2518 7019 2570 7025
rect 2518 6961 2570 6967
rect 2422 3763 2474 3769
rect 2422 3705 2474 3711
rect 2422 3245 2474 3251
rect 2422 3187 2474 3193
rect 2434 800 2462 3187
rect 2530 800 2558 6961
rect 2902 5687 2954 5693
rect 2902 5629 2954 5635
rect 2710 3689 2762 3695
rect 2710 3631 2762 3637
rect 2722 800 2750 3631
rect 2914 2900 2942 5629
rect 2818 2872 2942 2900
rect 2818 800 2846 2872
rect 3010 2752 3038 8219
rect 3286 7759 3338 7765
rect 3286 7701 3338 7707
rect 3190 6353 3242 6359
rect 3190 6295 3242 6301
rect 3094 5021 3146 5027
rect 3094 4963 3146 4969
rect 3106 3843 3134 4963
rect 3094 3837 3146 3843
rect 3094 3779 3146 3785
rect 3094 3541 3146 3547
rect 3094 3483 3146 3489
rect 2914 2724 3038 2752
rect 2914 800 2942 2724
rect 3106 1864 3134 3483
rect 3010 1836 3134 1864
rect 3010 800 3038 1836
rect 3202 800 3230 6295
rect 3298 800 3326 7701
rect 3586 7691 3614 29457
rect 4268 29332 4564 29352
rect 4324 29330 4348 29332
rect 4404 29330 4428 29332
rect 4484 29330 4508 29332
rect 4346 29278 4348 29330
rect 4410 29278 4422 29330
rect 4484 29278 4486 29330
rect 4324 29276 4348 29278
rect 4404 29276 4428 29278
rect 4484 29276 4508 29278
rect 4268 29256 4564 29276
rect 3670 28331 3722 28337
rect 3670 28273 3722 28279
rect 3682 8209 3710 28273
rect 4268 28000 4564 28020
rect 4324 27998 4348 28000
rect 4404 27998 4428 28000
rect 4484 27998 4508 28000
rect 4346 27946 4348 27998
rect 4410 27946 4422 27998
rect 4484 27946 4486 27998
rect 4324 27944 4348 27946
rect 4404 27944 4428 27946
rect 4484 27944 4508 27946
rect 4268 27924 4564 27944
rect 4268 26668 4564 26688
rect 4324 26666 4348 26668
rect 4404 26666 4428 26668
rect 4484 26666 4508 26668
rect 4346 26614 4348 26666
rect 4410 26614 4422 26666
rect 4484 26614 4486 26666
rect 4324 26612 4348 26614
rect 4404 26612 4428 26614
rect 4484 26612 4508 26614
rect 4268 26592 4564 26612
rect 4268 25336 4564 25356
rect 4324 25334 4348 25336
rect 4404 25334 4428 25336
rect 4484 25334 4508 25336
rect 4346 25282 4348 25334
rect 4410 25282 4422 25334
rect 4484 25282 4486 25334
rect 4324 25280 4348 25282
rect 4404 25280 4428 25282
rect 4484 25280 4508 25282
rect 4268 25260 4564 25280
rect 4268 24004 4564 24024
rect 4324 24002 4348 24004
rect 4404 24002 4428 24004
rect 4484 24002 4508 24004
rect 4346 23950 4348 24002
rect 4410 23950 4422 24002
rect 4484 23950 4486 24002
rect 4324 23948 4348 23950
rect 4404 23948 4428 23950
rect 4484 23948 4508 23950
rect 4268 23928 4564 23948
rect 4268 22672 4564 22692
rect 4324 22670 4348 22672
rect 4404 22670 4428 22672
rect 4484 22670 4508 22672
rect 4346 22618 4348 22670
rect 4410 22618 4422 22670
rect 4484 22618 4486 22670
rect 4324 22616 4348 22618
rect 4404 22616 4428 22618
rect 4484 22616 4508 22618
rect 4268 22596 4564 22616
rect 4268 21340 4564 21360
rect 4324 21338 4348 21340
rect 4404 21338 4428 21340
rect 4484 21338 4508 21340
rect 4346 21286 4348 21338
rect 4410 21286 4422 21338
rect 4484 21286 4486 21338
rect 4324 21284 4348 21286
rect 4404 21284 4428 21286
rect 4484 21284 4508 21286
rect 4268 21264 4564 21284
rect 4268 20008 4564 20028
rect 4324 20006 4348 20008
rect 4404 20006 4428 20008
rect 4484 20006 4508 20008
rect 4346 19954 4348 20006
rect 4410 19954 4422 20006
rect 4484 19954 4486 20006
rect 4324 19952 4348 19954
rect 4404 19952 4428 19954
rect 4484 19952 4508 19954
rect 4268 19932 4564 19952
rect 4150 19599 4202 19605
rect 4150 19541 4202 19547
rect 4162 17294 4190 19541
rect 4268 18676 4564 18696
rect 4324 18674 4348 18676
rect 4404 18674 4428 18676
rect 4484 18674 4508 18676
rect 4346 18622 4348 18674
rect 4410 18622 4422 18674
rect 4484 18622 4486 18674
rect 4324 18620 4348 18622
rect 4404 18620 4428 18622
rect 4484 18620 4508 18622
rect 4268 18600 4564 18620
rect 4066 17266 4190 17294
rect 4268 17344 4564 17364
rect 4324 17342 4348 17344
rect 4404 17342 4428 17344
rect 4484 17342 4508 17344
rect 4346 17290 4348 17342
rect 4410 17290 4422 17342
rect 4484 17290 4486 17342
rect 4324 17288 4348 17290
rect 4404 17288 4428 17290
rect 4484 17288 4508 17290
rect 4268 17268 4564 17288
rect 4066 10947 4094 17266
rect 4268 16012 4564 16032
rect 4324 16010 4348 16012
rect 4404 16010 4428 16012
rect 4484 16010 4508 16012
rect 4346 15958 4348 16010
rect 4410 15958 4422 16010
rect 4484 15958 4486 16010
rect 4324 15956 4348 15958
rect 4404 15956 4428 15958
rect 4484 15956 4508 15958
rect 4268 15936 4564 15956
rect 4268 14680 4564 14700
rect 4324 14678 4348 14680
rect 4404 14678 4428 14680
rect 4484 14678 4508 14680
rect 4346 14626 4348 14678
rect 4410 14626 4422 14678
rect 4484 14626 4486 14678
rect 4324 14624 4348 14626
rect 4404 14624 4428 14626
rect 4484 14624 4508 14626
rect 4268 14604 4564 14624
rect 4150 13457 4202 13463
rect 4150 13399 4202 13405
rect 4054 10941 4106 10947
rect 4054 10883 4106 10889
rect 3670 8203 3722 8209
rect 3670 8145 3722 8151
rect 4054 7759 4106 7765
rect 4054 7701 4106 7707
rect 3574 7685 3626 7691
rect 3574 7627 3626 7633
rect 3382 7463 3434 7469
rect 3382 7405 3434 7411
rect 3394 3917 3422 7405
rect 3670 6871 3722 6877
rect 3670 6813 3722 6819
rect 3382 3911 3434 3917
rect 3382 3853 3434 3859
rect 3382 3763 3434 3769
rect 3382 3705 3434 3711
rect 3394 800 3422 3705
rect 3478 3171 3530 3177
rect 3478 3113 3530 3119
rect 3490 800 3518 3113
rect 3682 800 3710 6813
rect 3862 6353 3914 6359
rect 3862 6295 3914 6301
rect 3766 4281 3818 4287
rect 3766 4223 3818 4229
rect 3778 800 3806 4223
rect 3874 800 3902 6295
rect 3958 3467 4010 3473
rect 3958 3409 4010 3415
rect 3970 2585 3998 3409
rect 3958 2579 4010 2585
rect 3958 2521 4010 2527
rect 4066 800 4094 7701
rect 4162 7617 4190 13399
rect 4268 13348 4564 13368
rect 4324 13346 4348 13348
rect 4404 13346 4428 13348
rect 4484 13346 4508 13348
rect 4346 13294 4348 13346
rect 4410 13294 4422 13346
rect 4484 13294 4486 13346
rect 4324 13292 4348 13294
rect 4404 13292 4428 13294
rect 4484 13292 4508 13294
rect 4268 13272 4564 13292
rect 4268 12016 4564 12036
rect 4324 12014 4348 12016
rect 4404 12014 4428 12016
rect 4484 12014 4508 12016
rect 4346 11962 4348 12014
rect 4410 11962 4422 12014
rect 4484 11962 4486 12014
rect 4324 11960 4348 11962
rect 4404 11960 4428 11962
rect 4484 11960 4508 11962
rect 4268 11940 4564 11960
rect 4268 10684 4564 10704
rect 4324 10682 4348 10684
rect 4404 10682 4428 10684
rect 4484 10682 4508 10684
rect 4346 10630 4348 10682
rect 4410 10630 4422 10682
rect 4484 10630 4486 10682
rect 4324 10628 4348 10630
rect 4404 10628 4428 10630
rect 4484 10628 4508 10630
rect 4268 10608 4564 10628
rect 4268 9352 4564 9372
rect 4324 9350 4348 9352
rect 4404 9350 4428 9352
rect 4484 9350 4508 9352
rect 4346 9298 4348 9350
rect 4410 9298 4422 9350
rect 4484 9298 4486 9350
rect 4324 9296 4348 9298
rect 4404 9296 4428 9298
rect 4484 9296 4508 9298
rect 4268 9276 4564 9296
rect 4268 8020 4564 8040
rect 4324 8018 4348 8020
rect 4404 8018 4428 8020
rect 4484 8018 4508 8020
rect 4346 7966 4348 8018
rect 4410 7966 4422 8018
rect 4484 7966 4486 8018
rect 4324 7964 4348 7966
rect 4404 7964 4428 7966
rect 4484 7964 4508 7966
rect 4268 7944 4564 7964
rect 4150 7611 4202 7617
rect 4150 7553 4202 7559
rect 4268 6688 4564 6708
rect 4324 6686 4348 6688
rect 4404 6686 4428 6688
rect 4484 6686 4508 6688
rect 4346 6634 4348 6686
rect 4410 6634 4422 6686
rect 4484 6634 4486 6686
rect 4324 6632 4348 6634
rect 4404 6632 4428 6634
rect 4484 6632 4508 6634
rect 4268 6612 4564 6632
rect 4642 6452 4670 47506
rect 5218 41435 5246 56689
rect 5410 56531 5438 59200
rect 5782 56747 5834 56753
rect 5782 56689 5834 56695
rect 5398 56525 5450 56531
rect 5398 56467 5450 56473
rect 5590 56229 5642 56235
rect 5590 56171 5642 56177
rect 5398 55563 5450 55569
rect 5398 55505 5450 55511
rect 5410 48539 5438 55505
rect 5602 50167 5630 56171
rect 5794 56161 5822 56689
rect 5986 56531 6014 59200
rect 6466 56975 6494 59200
rect 6454 56969 6506 56975
rect 6454 56911 6506 56917
rect 6070 56821 6122 56827
rect 6070 56763 6122 56769
rect 5974 56525 6026 56531
rect 5974 56467 6026 56473
rect 5782 56155 5834 56161
rect 5782 56097 5834 56103
rect 5590 50161 5642 50167
rect 5590 50103 5642 50109
rect 5398 48533 5450 48539
rect 5398 48475 5450 48481
rect 6082 48465 6110 56763
rect 7042 56531 7070 59200
rect 7318 56747 7370 56753
rect 7318 56689 7370 56695
rect 7030 56525 7082 56531
rect 7030 56467 7082 56473
rect 6358 56229 6410 56235
rect 6358 56171 6410 56177
rect 7222 56229 7274 56235
rect 7222 56171 7274 56177
rect 6070 48459 6122 48465
rect 6070 48401 6122 48407
rect 6370 44099 6398 56171
rect 6934 48755 6986 48761
rect 6934 48697 6986 48703
rect 6358 44093 6410 44099
rect 6358 44035 6410 44041
rect 5206 41429 5258 41435
rect 5206 41371 5258 41377
rect 6838 32549 6890 32555
rect 6838 32491 6890 32497
rect 6550 32401 6602 32407
rect 6550 32343 6602 32349
rect 6562 31889 6590 32343
rect 6550 31883 6602 31889
rect 6550 31825 6602 31831
rect 6850 31815 6878 32491
rect 6838 31809 6890 31815
rect 6838 31751 6890 31757
rect 6262 28109 6314 28115
rect 6262 28051 6314 28057
rect 5398 25445 5450 25451
rect 5398 25387 5450 25393
rect 5410 25155 5438 25387
rect 5398 25149 5450 25155
rect 5398 25091 5450 25097
rect 5974 20117 6026 20123
rect 5974 20059 6026 20065
rect 5878 19451 5930 19457
rect 5878 19393 5930 19399
rect 5890 19328 5918 19393
rect 5842 19300 5918 19328
rect 5842 19161 5870 19300
rect 5986 19235 6014 20059
rect 6166 19747 6218 19753
rect 6166 19689 6218 19695
rect 6178 19328 6206 19689
rect 6130 19300 6206 19328
rect 5974 19229 6026 19235
rect 5974 19171 6026 19177
rect 6130 19161 6158 19300
rect 5830 19155 5882 19161
rect 5830 19097 5882 19103
rect 6118 19155 6170 19161
rect 6118 19097 6170 19103
rect 6070 12421 6122 12427
rect 6070 12363 6122 12369
rect 5494 9757 5546 9763
rect 5494 9699 5546 9705
rect 5506 9171 5534 9699
rect 5494 9165 5546 9171
rect 5494 9107 5546 9113
rect 4822 8277 4874 8283
rect 4822 8219 4874 8225
rect 4642 6424 4766 6452
rect 4630 6353 4682 6359
rect 4630 6295 4682 6301
rect 4268 5356 4564 5376
rect 4324 5354 4348 5356
rect 4404 5354 4428 5356
rect 4484 5354 4508 5356
rect 4346 5302 4348 5354
rect 4410 5302 4422 5354
rect 4484 5302 4486 5354
rect 4324 5300 4348 5302
rect 4404 5300 4428 5302
rect 4484 5300 4508 5302
rect 4268 5280 4564 5300
rect 4150 5021 4202 5027
rect 4150 4963 4202 4969
rect 4162 800 4190 4963
rect 4642 4676 4670 6295
rect 4546 4648 4670 4676
rect 4546 4232 4574 4648
rect 4738 4509 4766 6424
rect 4726 4503 4778 4509
rect 4726 4445 4778 4451
rect 4726 4355 4778 4361
rect 4726 4297 4778 4303
rect 4546 4204 4670 4232
rect 4268 4024 4564 4044
rect 4324 4022 4348 4024
rect 4404 4022 4428 4024
rect 4484 4022 4508 4024
rect 4346 3970 4348 4022
rect 4410 3970 4422 4022
rect 4484 3970 4486 4022
rect 4324 3968 4348 3970
rect 4404 3968 4428 3970
rect 4484 3968 4508 3970
rect 4268 3948 4564 3968
rect 4268 2692 4564 2712
rect 4324 2690 4348 2692
rect 4404 2690 4428 2692
rect 4484 2690 4508 2692
rect 4346 2638 4348 2690
rect 4410 2638 4422 2690
rect 4484 2638 4486 2690
rect 4324 2636 4348 2638
rect 4404 2636 4428 2638
rect 4484 2636 4508 2638
rect 4268 2616 4564 2636
rect 4246 2579 4298 2585
rect 4246 2521 4298 2527
rect 4342 2579 4394 2585
rect 4342 2521 4394 2527
rect 4258 800 4286 2521
rect 4354 800 4382 2521
rect 4642 2456 4670 4204
rect 4450 2428 4670 2456
rect 4450 2012 4478 2428
rect 4738 2160 4766 4297
rect 4834 2585 4862 8219
rect 5302 7463 5354 7469
rect 5302 7405 5354 7411
rect 5110 6945 5162 6951
rect 5162 6905 5246 6933
rect 5110 6887 5162 6893
rect 4918 5687 4970 5693
rect 4918 5629 4970 5635
rect 5110 5687 5162 5693
rect 5110 5629 5162 5635
rect 4930 3177 4958 5629
rect 5014 4281 5066 4287
rect 5014 4223 5066 4229
rect 4918 3171 4970 3177
rect 4918 3113 4970 3119
rect 4918 3023 4970 3029
rect 4918 2965 4970 2971
rect 4822 2579 4874 2585
rect 4822 2521 4874 2527
rect 4738 2132 4862 2160
rect 4726 2061 4778 2067
rect 4450 1984 4670 2012
rect 4726 2003 4778 2009
rect 4534 1913 4586 1919
rect 4534 1855 4586 1861
rect 4546 800 4574 1855
rect 4642 800 4670 1984
rect 4738 800 4766 2003
rect 4834 1919 4862 2132
rect 4822 1913 4874 1919
rect 4822 1855 4874 1861
rect 4930 800 4958 2965
rect 5026 800 5054 4223
rect 5122 3473 5150 5629
rect 5110 3467 5162 3473
rect 5110 3409 5162 3415
rect 5218 3251 5246 6905
rect 5206 3245 5258 3251
rect 5206 3187 5258 3193
rect 5110 3171 5162 3177
rect 5110 3113 5162 3119
rect 5122 800 5150 3113
rect 5206 3023 5258 3029
rect 5206 2965 5258 2971
rect 5218 800 5246 2965
rect 5314 2067 5342 7405
rect 5686 6945 5738 6951
rect 5686 6887 5738 6893
rect 5878 6945 5930 6951
rect 5878 6887 5930 6893
rect 5494 6131 5546 6137
rect 5494 6073 5546 6079
rect 5398 5021 5450 5027
rect 5398 4963 5450 4969
rect 5302 2061 5354 2067
rect 5302 2003 5354 2009
rect 5410 800 5438 4963
rect 5506 800 5534 6073
rect 5698 5841 5726 6887
rect 5686 5835 5738 5841
rect 5686 5777 5738 5783
rect 5686 4281 5738 4287
rect 5686 4223 5738 4229
rect 5590 3689 5642 3695
rect 5590 3631 5642 3637
rect 5602 800 5630 3631
rect 5698 800 5726 4223
rect 5890 800 5918 6887
rect 6082 5767 6110 12363
rect 6274 12353 6302 28051
rect 6550 26851 6602 26857
rect 6550 26793 6602 26799
rect 6454 19525 6506 19531
rect 6454 19467 6506 19473
rect 6466 19328 6494 19467
rect 6418 19300 6494 19328
rect 6418 19161 6446 19300
rect 6406 19155 6458 19161
rect 6406 19097 6458 19103
rect 6562 17294 6590 26793
rect 6946 17294 6974 48697
rect 7234 40399 7262 56171
rect 7330 41583 7358 56689
rect 7522 55717 7550 59200
rect 8098 56975 8126 59200
rect 8086 56969 8138 56975
rect 8086 56911 8138 56917
rect 7894 56895 7946 56901
rect 7894 56837 7946 56843
rect 7510 55711 7562 55717
rect 7510 55653 7562 55659
rect 7702 55563 7754 55569
rect 7702 55505 7754 55511
rect 7606 43797 7658 43803
rect 7606 43739 7658 43745
rect 7318 41577 7370 41583
rect 7318 41519 7370 41525
rect 7222 40393 7274 40399
rect 7222 40335 7274 40341
rect 7126 23447 7178 23453
rect 7126 23389 7178 23395
rect 6466 17266 6590 17294
rect 6850 17266 6974 17294
rect 6262 12347 6314 12353
rect 6262 12289 6314 12295
rect 6466 7173 6494 17266
rect 6850 7543 6878 17266
rect 6934 10793 6986 10799
rect 6934 10735 6986 10741
rect 6946 10503 6974 10735
rect 6934 10497 6986 10503
rect 6934 10439 6986 10445
rect 6838 7537 6890 7543
rect 6838 7479 6890 7485
rect 6454 7167 6506 7173
rect 6454 7109 6506 7115
rect 6166 6945 6218 6951
rect 6166 6887 6218 6893
rect 6550 6945 6602 6951
rect 6550 6887 6602 6893
rect 6178 6581 6206 6887
rect 6166 6575 6218 6581
rect 6166 6517 6218 6523
rect 6262 6131 6314 6137
rect 6262 6073 6314 6079
rect 6070 5761 6122 5767
rect 6070 5703 6122 5709
rect 5974 5613 6026 5619
rect 5974 5555 6026 5561
rect 5986 3177 6014 5555
rect 6070 5021 6122 5027
rect 6070 4963 6122 4969
rect 5974 3171 6026 3177
rect 5974 3113 6026 3119
rect 5974 3023 6026 3029
rect 5974 2965 6026 2971
rect 5986 800 6014 2965
rect 6082 800 6110 4963
rect 6166 4207 6218 4213
rect 6166 4149 6218 4155
rect 6178 3177 6206 4149
rect 6166 3171 6218 3177
rect 6166 3113 6218 3119
rect 6274 800 6302 6073
rect 6454 4207 6506 4213
rect 6454 4149 6506 4155
rect 6358 3689 6410 3695
rect 6358 3631 6410 3637
rect 6370 800 6398 3631
rect 6466 800 6494 4149
rect 6562 800 6590 6887
rect 7138 6433 7166 23389
rect 7510 8129 7562 8135
rect 7510 8071 7562 8077
rect 7318 6945 7370 6951
rect 7318 6887 7370 6893
rect 7126 6427 7178 6433
rect 7126 6369 7178 6375
rect 6934 6205 6986 6211
rect 6934 6147 6986 6153
rect 6838 3097 6890 3103
rect 6838 3039 6890 3045
rect 6742 2949 6794 2955
rect 6742 2891 6794 2897
rect 6754 800 6782 2891
rect 6850 800 6878 3039
rect 6946 800 6974 6147
rect 7222 5687 7274 5693
rect 7222 5629 7274 5635
rect 7030 3689 7082 3695
rect 7030 3631 7082 3637
rect 7042 800 7070 3631
rect 7234 800 7262 5629
rect 7330 800 7358 6887
rect 7522 5767 7550 8071
rect 7618 7099 7646 43739
rect 7714 11909 7742 55505
rect 7906 22343 7934 56837
rect 8578 56531 8606 59200
rect 9046 56821 9098 56827
rect 9046 56763 9098 56769
rect 8566 56525 8618 56531
rect 8566 56467 8618 56473
rect 8566 56229 8618 56235
rect 8566 56171 8618 56177
rect 8578 40991 8606 56171
rect 8566 40985 8618 40991
rect 8566 40927 8618 40933
rect 7990 36101 8042 36107
rect 7990 36043 8042 36049
rect 7894 22337 7946 22343
rect 7894 22279 7946 22285
rect 7702 11903 7754 11909
rect 7702 11845 7754 11851
rect 8002 7173 8030 36043
rect 9058 33240 9086 56763
rect 9154 55717 9182 59200
rect 9634 56975 9662 59200
rect 9622 56969 9674 56975
rect 9622 56911 9674 56917
rect 10006 56747 10058 56753
rect 10006 56689 10058 56695
rect 9142 55711 9194 55717
rect 9142 55653 9194 55659
rect 9334 55563 9386 55569
rect 9334 55505 9386 55511
rect 9346 41509 9374 55505
rect 9334 41503 9386 41509
rect 9334 41445 9386 41451
rect 9334 33881 9386 33887
rect 9334 33823 9386 33829
rect 9010 33212 9086 33240
rect 9010 33073 9038 33212
rect 8998 33067 9050 33073
rect 8998 33009 9050 33015
rect 8854 32771 8906 32777
rect 8854 32713 8906 32719
rect 8866 32555 8894 32713
rect 8854 32549 8906 32555
rect 8854 32491 8906 32497
rect 8566 23595 8618 23601
rect 8566 23537 8618 23543
rect 8578 22491 8606 23537
rect 8758 22781 8810 22787
rect 8758 22723 8810 22729
rect 8566 22485 8618 22491
rect 8566 22427 8618 22433
rect 7990 7167 8042 7173
rect 7990 7109 8042 7115
rect 7606 7093 7658 7099
rect 7606 7035 7658 7041
rect 8086 6945 8138 6951
rect 8086 6887 8138 6893
rect 7990 6205 8042 6211
rect 7990 6147 8042 6153
rect 7510 5761 7562 5767
rect 7510 5703 7562 5709
rect 7894 5687 7946 5693
rect 7894 5629 7946 5635
rect 7702 5021 7754 5027
rect 7702 4963 7754 4969
rect 7606 4947 7658 4953
rect 7606 4889 7658 4895
rect 7414 4355 7466 4361
rect 7414 4297 7466 4303
rect 7426 800 7454 4297
rect 7618 800 7646 4889
rect 7714 3103 7742 4963
rect 7798 3689 7850 3695
rect 7798 3631 7850 3637
rect 7702 3097 7754 3103
rect 7702 3039 7754 3045
rect 7702 2949 7754 2955
rect 7702 2891 7754 2897
rect 7714 800 7742 2891
rect 7810 800 7838 3631
rect 7906 800 7934 5629
rect 8002 2955 8030 6147
rect 7990 2949 8042 2955
rect 7990 2891 8042 2897
rect 8098 800 8126 6887
rect 8470 6427 8522 6433
rect 8470 6369 8522 6375
rect 8278 3837 8330 3843
rect 8278 3779 8330 3785
rect 8182 3023 8234 3029
rect 8182 2965 8234 2971
rect 8194 800 8222 2965
rect 8290 800 8318 3779
rect 8482 800 8510 6369
rect 8770 6359 8798 22723
rect 9346 8431 9374 33823
rect 10018 33147 10046 56689
rect 10210 56531 10238 59200
rect 10690 56531 10718 59200
rect 11266 56975 11294 59200
rect 11254 56969 11306 56975
rect 11254 56911 11306 56917
rect 11746 56531 11774 59200
rect 12322 56531 12350 59200
rect 12802 56975 12830 59200
rect 12790 56969 12842 56975
rect 12790 56911 12842 56917
rect 13078 56747 13130 56753
rect 13078 56689 13130 56695
rect 10198 56525 10250 56531
rect 10198 56467 10250 56473
rect 10678 56525 10730 56531
rect 10678 56467 10730 56473
rect 11734 56525 11786 56531
rect 11734 56467 11786 56473
rect 12310 56525 12362 56531
rect 12310 56467 12362 56473
rect 10102 56229 10154 56235
rect 10102 56171 10154 56177
rect 11158 56229 11210 56235
rect 11158 56171 11210 56177
rect 11926 56229 11978 56235
rect 11926 56171 11978 56177
rect 12310 56229 12362 56235
rect 12310 56171 12362 56177
rect 10006 33141 10058 33147
rect 10006 33083 10058 33089
rect 9430 21449 9482 21455
rect 9430 21391 9482 21397
rect 9442 14203 9470 21391
rect 9430 14197 9482 14203
rect 9430 14139 9482 14145
rect 10114 14129 10142 56171
rect 11170 54533 11198 56171
rect 11158 54527 11210 54533
rect 11158 54469 11210 54475
rect 11062 50827 11114 50833
rect 11062 50769 11114 50775
rect 10870 25593 10922 25599
rect 10870 25535 10922 25541
rect 10198 16787 10250 16793
rect 10198 16729 10250 16735
rect 10102 14123 10154 14129
rect 10102 14065 10154 14071
rect 9334 8425 9386 8431
rect 9334 8367 9386 8373
rect 10210 7765 10238 16729
rect 10774 10127 10826 10133
rect 10774 10069 10826 10075
rect 10786 8431 10814 10069
rect 10774 8425 10826 8431
rect 10774 8367 10826 8373
rect 10582 8277 10634 8283
rect 10582 8219 10634 8225
rect 10198 7759 10250 7765
rect 10198 7701 10250 7707
rect 9142 7463 9194 7469
rect 9142 7405 9194 7411
rect 9910 7463 9962 7469
rect 9910 7405 9962 7411
rect 8854 6945 8906 6951
rect 8854 6887 8906 6893
rect 8758 6353 8810 6359
rect 8758 6295 8810 6301
rect 8566 6279 8618 6285
rect 8566 6221 8618 6227
rect 8578 4879 8606 6221
rect 8566 4873 8618 4879
rect 8566 4815 8618 4821
rect 8758 3911 8810 3917
rect 8758 3853 8810 3859
rect 8566 3689 8618 3695
rect 8770 3640 8798 3853
rect 8566 3631 8618 3637
rect 8578 800 8606 3631
rect 8674 3612 8798 3640
rect 8674 800 8702 3612
rect 8866 3492 8894 6887
rect 9046 5687 9098 5693
rect 9046 5629 9098 5635
rect 8770 3464 8894 3492
rect 8770 800 8798 3464
rect 8950 3097 9002 3103
rect 8950 3039 9002 3045
rect 8962 800 8990 3039
rect 9058 800 9086 5629
rect 9154 800 9182 7405
rect 9526 6871 9578 6877
rect 9526 6813 9578 6819
rect 9238 5021 9290 5027
rect 9238 4963 9290 4969
rect 9250 3843 9278 4963
rect 9238 3837 9290 3843
rect 9238 3779 9290 3785
rect 9334 3689 9386 3695
rect 9250 3649 9334 3677
rect 9250 800 9278 3649
rect 9334 3631 9386 3637
rect 9430 3245 9482 3251
rect 9430 3187 9482 3193
rect 9442 800 9470 3187
rect 9538 800 9566 6813
rect 9622 4355 9674 4361
rect 9622 4297 9674 4303
rect 9634 800 9662 4297
rect 9814 2949 9866 2955
rect 9814 2891 9866 2897
rect 9826 800 9854 2891
rect 9922 800 9950 7405
rect 10102 6353 10154 6359
rect 10102 6295 10154 6301
rect 10006 3541 10058 3547
rect 10006 3483 10058 3489
rect 10018 800 10046 3483
rect 10114 800 10142 6295
rect 10198 5687 10250 5693
rect 10198 5629 10250 5635
rect 10486 5687 10538 5693
rect 10486 5629 10538 5635
rect 10210 2955 10238 5629
rect 10294 5021 10346 5027
rect 10294 4963 10346 4969
rect 10306 3917 10334 4963
rect 10390 4355 10442 4361
rect 10390 4297 10442 4303
rect 10294 3911 10346 3917
rect 10294 3853 10346 3859
rect 10294 3763 10346 3769
rect 10294 3705 10346 3711
rect 10198 2949 10250 2955
rect 10198 2891 10250 2897
rect 10306 800 10334 3705
rect 10402 800 10430 4297
rect 10498 800 10526 5629
rect 10594 800 10622 8219
rect 10882 7765 10910 25535
rect 11074 17294 11102 50769
rect 11938 17607 11966 56171
rect 12214 49421 12266 49427
rect 12214 49363 12266 49369
rect 11926 17601 11978 17607
rect 11926 17543 11978 17549
rect 12226 17294 12254 49363
rect 11074 17266 11486 17294
rect 10966 8277 11018 8283
rect 10966 8219 11018 8225
rect 10870 7759 10922 7765
rect 10870 7701 10922 7707
rect 10870 6353 10922 6359
rect 10870 6295 10922 6301
rect 10678 5021 10730 5027
rect 10678 4963 10730 4969
rect 10690 3251 10718 4963
rect 10774 4355 10826 4361
rect 10774 4297 10826 4303
rect 10678 3245 10730 3251
rect 10678 3187 10730 3193
rect 10786 800 10814 4297
rect 10882 800 10910 6295
rect 10978 800 11006 8219
rect 11350 7759 11402 7765
rect 11350 7701 11402 7707
rect 11062 7463 11114 7469
rect 11062 7405 11114 7411
rect 11074 3769 11102 7405
rect 11254 7019 11306 7025
rect 11254 6961 11306 6967
rect 11158 4207 11210 4213
rect 11158 4149 11210 4155
rect 11062 3763 11114 3769
rect 11062 3705 11114 3711
rect 11170 800 11198 4149
rect 11266 800 11294 6961
rect 11362 800 11390 7701
rect 11458 4232 11486 17266
rect 12130 17266 12254 17294
rect 12322 17294 12350 56171
rect 12406 55563 12458 55569
rect 12406 55505 12458 55511
rect 12418 55199 12446 55505
rect 12406 55193 12458 55199
rect 12406 55135 12458 55141
rect 12790 46165 12842 46171
rect 12790 46107 12842 46113
rect 12322 17266 12542 17294
rect 11542 14567 11594 14573
rect 11542 14509 11594 14515
rect 11554 8431 11582 14509
rect 11542 8425 11594 8431
rect 11542 8367 11594 8373
rect 11734 8277 11786 8283
rect 11734 8219 11786 8225
rect 11638 6353 11690 6359
rect 11638 6295 11690 6301
rect 11458 4204 11582 4232
rect 11446 4133 11498 4139
rect 11446 4075 11498 4081
rect 11458 800 11486 4075
rect 11554 2955 11582 4204
rect 11542 2949 11594 2955
rect 11542 2891 11594 2897
rect 11650 800 11678 6295
rect 11746 800 11774 8219
rect 12130 6581 12158 17266
rect 12514 9467 12542 17266
rect 12598 14271 12650 14277
rect 12598 14213 12650 14219
rect 12610 13833 12638 14213
rect 12598 13827 12650 13833
rect 12598 13769 12650 13775
rect 12502 9461 12554 9467
rect 12502 9403 12554 9409
rect 12310 9091 12362 9097
rect 12310 9033 12362 9039
rect 12322 8431 12350 9033
rect 12310 8425 12362 8431
rect 12310 8367 12362 8373
rect 12502 8277 12554 8283
rect 12502 8219 12554 8225
rect 12406 8129 12458 8135
rect 12406 8071 12458 8077
rect 12418 7913 12446 8071
rect 12406 7907 12458 7913
rect 12406 7849 12458 7855
rect 12418 7765 12446 7849
rect 12406 7759 12458 7765
rect 12406 7701 12458 7707
rect 12214 7463 12266 7469
rect 12214 7405 12266 7411
rect 12118 6575 12170 6581
rect 12118 6517 12170 6523
rect 12118 5465 12170 5471
rect 12118 5407 12170 5413
rect 12130 5101 12158 5407
rect 12118 5095 12170 5101
rect 12118 5037 12170 5043
rect 11830 5021 11882 5027
rect 11830 4963 11882 4969
rect 11842 800 11870 4963
rect 12022 3837 12074 3843
rect 12022 3779 12074 3785
rect 12034 800 12062 3779
rect 12226 3640 12254 7405
rect 12310 6353 12362 6359
rect 12310 6295 12362 6301
rect 12130 3612 12254 3640
rect 12130 800 12158 3612
rect 12214 3245 12266 3251
rect 12214 3187 12266 3193
rect 12226 800 12254 3187
rect 12322 800 12350 6295
rect 12514 800 12542 8219
rect 12802 7932 12830 46107
rect 13090 33073 13118 56689
rect 13378 56531 13406 59200
rect 13654 56747 13706 56753
rect 13654 56689 13706 56695
rect 13366 56525 13418 56531
rect 13366 56467 13418 56473
rect 13558 56229 13610 56235
rect 13558 56171 13610 56177
rect 13570 38401 13598 56171
rect 13558 38395 13610 38401
rect 13558 38337 13610 38343
rect 13078 33067 13130 33073
rect 13078 33009 13130 33015
rect 13078 32105 13130 32111
rect 13078 32047 13130 32053
rect 13090 21011 13118 32047
rect 13666 28263 13694 56689
rect 13858 55717 13886 59200
rect 14434 56975 14462 59200
rect 14422 56969 14474 56975
rect 14422 56911 14474 56917
rect 14914 56531 14942 59200
rect 15394 56531 15422 59200
rect 15970 57049 15998 59200
rect 16450 57123 16478 59200
rect 16438 57117 16490 57123
rect 16438 57059 16490 57065
rect 15958 57043 16010 57049
rect 15958 56985 16010 56991
rect 16054 56747 16106 56753
rect 16054 56689 16106 56695
rect 14902 56525 14954 56531
rect 14902 56467 14954 56473
rect 15382 56525 15434 56531
rect 15382 56467 15434 56473
rect 15190 56229 15242 56235
rect 15190 56171 15242 56177
rect 15286 56229 15338 56235
rect 15286 56171 15338 56177
rect 13846 55711 13898 55717
rect 13846 55653 13898 55659
rect 13846 55415 13898 55421
rect 13846 55357 13898 55363
rect 13750 46165 13802 46171
rect 13750 46107 13802 46113
rect 13654 28257 13706 28263
rect 13654 28199 13706 28205
rect 13558 25223 13610 25229
rect 13558 25165 13610 25171
rect 13078 21005 13130 21011
rect 13078 20947 13130 20953
rect 12982 14493 13034 14499
rect 12982 14435 13034 14441
rect 12994 10133 13022 14435
rect 12982 10127 13034 10133
rect 12982 10069 13034 10075
rect 12802 7913 12926 7932
rect 13570 7913 13598 25165
rect 13654 23595 13706 23601
rect 13654 23537 13706 23543
rect 13666 22417 13694 23537
rect 13654 22411 13706 22417
rect 13654 22353 13706 22359
rect 13762 8135 13790 46107
rect 13858 25747 13886 55357
rect 14998 50827 15050 50833
rect 14998 50769 15050 50775
rect 14038 50753 14090 50759
rect 14038 50695 14090 50701
rect 13846 25741 13898 25747
rect 13846 25683 13898 25689
rect 13942 19599 13994 19605
rect 13942 19541 13994 19547
rect 13954 18125 13982 19541
rect 13942 18119 13994 18125
rect 13942 18061 13994 18067
rect 13942 12495 13994 12501
rect 13942 12437 13994 12443
rect 13846 11163 13898 11169
rect 13846 11105 13898 11111
rect 13750 8129 13802 8135
rect 13750 8071 13802 8077
rect 12790 7907 12926 7913
rect 12842 7904 12926 7907
rect 12790 7849 12842 7855
rect 12790 7759 12842 7765
rect 12790 7701 12842 7707
rect 12694 7019 12746 7025
rect 12694 6961 12746 6967
rect 12598 5687 12650 5693
rect 12598 5629 12650 5635
rect 12610 800 12638 5629
rect 12706 800 12734 6961
rect 12802 800 12830 7701
rect 12898 7617 12926 7904
rect 13558 7907 13610 7913
rect 13558 7849 13610 7855
rect 13570 7765 13598 7849
rect 13558 7759 13610 7765
rect 13558 7701 13610 7707
rect 12886 7611 12938 7617
rect 12886 7553 12938 7559
rect 13462 6945 13514 6951
rect 13462 6887 13514 6893
rect 13654 6945 13706 6951
rect 13654 6887 13706 6893
rect 13270 6131 13322 6137
rect 13270 6073 13322 6079
rect 12982 5021 13034 5027
rect 12982 4963 13034 4969
rect 12994 3251 13022 4963
rect 13174 3689 13226 3695
rect 13174 3631 13226 3637
rect 12982 3245 13034 3251
rect 12982 3187 13034 3193
rect 12994 3029 13118 3048
rect 12994 3023 13130 3029
rect 12994 3020 13078 3023
rect 12994 800 13022 3020
rect 13078 2965 13130 2971
rect 13186 2894 13214 3631
rect 13090 2866 13214 2894
rect 13090 1864 13118 2866
rect 13090 1836 13214 1864
rect 13078 1765 13130 1771
rect 13078 1707 13130 1713
rect 13090 800 13118 1707
rect 13186 800 13214 1836
rect 13282 1771 13310 6073
rect 13366 5687 13418 5693
rect 13366 5629 13418 5635
rect 13378 3843 13406 5629
rect 13366 3837 13418 3843
rect 13366 3779 13418 3785
rect 13366 3689 13418 3695
rect 13366 3631 13418 3637
rect 13270 1765 13322 1771
rect 13270 1707 13322 1713
rect 13378 800 13406 3631
rect 13474 800 13502 6887
rect 13558 4355 13610 4361
rect 13558 4297 13610 4303
rect 13570 800 13598 4297
rect 13666 3843 13694 6887
rect 13858 5268 13886 11105
rect 13954 6433 13982 12437
rect 13942 6427 13994 6433
rect 13942 6369 13994 6375
rect 13942 6131 13994 6137
rect 13942 6073 13994 6079
rect 13762 5240 13886 5268
rect 13654 3837 13706 3843
rect 13654 3779 13706 3785
rect 13654 3615 13706 3621
rect 13654 3557 13706 3563
rect 13666 800 13694 3557
rect 13762 2955 13790 5240
rect 13954 5120 13982 6073
rect 13858 5092 13982 5120
rect 13750 2949 13802 2955
rect 13750 2891 13802 2897
rect 13858 800 13886 5092
rect 13942 5021 13994 5027
rect 13942 4963 13994 4969
rect 13954 800 13982 4963
rect 14050 3473 14078 50695
rect 14614 11607 14666 11613
rect 14614 11549 14666 11555
rect 14230 10423 14282 10429
rect 14230 10365 14282 10371
rect 14134 6205 14186 6211
rect 14134 6147 14186 6153
rect 14038 3467 14090 3473
rect 14038 3409 14090 3415
rect 14038 3023 14090 3029
rect 14038 2965 14090 2971
rect 14050 800 14078 2965
rect 14146 800 14174 6147
rect 14242 3769 14270 10365
rect 14626 9837 14654 11549
rect 14614 9831 14666 9837
rect 14614 9773 14666 9779
rect 14710 8943 14762 8949
rect 14710 8885 14762 8891
rect 14518 6945 14570 6951
rect 14518 6887 14570 6893
rect 14422 5021 14474 5027
rect 14422 4963 14474 4969
rect 14434 3936 14462 4963
rect 14338 3908 14462 3936
rect 14230 3763 14282 3769
rect 14230 3705 14282 3711
rect 14338 800 14366 3908
rect 14422 3763 14474 3769
rect 14422 3705 14474 3711
rect 14434 800 14462 3705
rect 14530 800 14558 6887
rect 14722 6433 14750 8885
rect 15010 7913 15038 50769
rect 15202 38179 15230 56171
rect 15190 38173 15242 38179
rect 15190 38115 15242 38121
rect 15298 32555 15326 56171
rect 15286 32549 15338 32555
rect 15286 32491 15338 32497
rect 15190 28109 15242 28115
rect 15190 28051 15242 28057
rect 15094 22263 15146 22269
rect 15094 22205 15146 22211
rect 15106 15757 15134 22205
rect 15094 15751 15146 15757
rect 15094 15693 15146 15699
rect 14998 7907 15050 7913
rect 14998 7849 15050 7855
rect 15010 7765 15038 7849
rect 14998 7759 15050 7765
rect 14998 7701 15050 7707
rect 15202 7099 15230 28051
rect 16066 19161 16094 56689
rect 17026 56531 17054 59200
rect 17506 57049 17534 59200
rect 18082 57614 18110 59200
rect 18082 57586 18206 57614
rect 17494 57043 17546 57049
rect 17494 56985 17546 56991
rect 17878 56747 17930 56753
rect 17878 56689 17930 56695
rect 17014 56525 17066 56531
rect 17014 56467 17066 56473
rect 16822 56229 16874 56235
rect 16822 56171 16874 56177
rect 16342 52751 16394 52757
rect 16342 52693 16394 52699
rect 16054 19155 16106 19161
rect 16054 19097 16106 19103
rect 16354 17294 16382 52693
rect 16438 37433 16490 37439
rect 16438 37375 16490 37381
rect 16258 17266 16382 17294
rect 15862 15899 15914 15905
rect 15862 15841 15914 15847
rect 15478 15529 15530 15535
rect 15478 15471 15530 15477
rect 15286 7463 15338 7469
rect 15286 7405 15338 7411
rect 15190 7093 15242 7099
rect 15190 7035 15242 7041
rect 15094 6945 15146 6951
rect 14914 6905 15094 6933
rect 14710 6427 14762 6433
rect 14710 6369 14762 6375
rect 14806 5021 14858 5027
rect 14806 4963 14858 4969
rect 14818 3936 14846 4963
rect 14626 3908 14846 3936
rect 14626 2604 14654 3908
rect 14806 3023 14858 3029
rect 14806 2965 14858 2971
rect 14626 2576 14750 2604
rect 14722 800 14750 2576
rect 14818 800 14846 2965
rect 14914 800 14942 6905
rect 15094 6887 15146 6893
rect 14998 5687 15050 5693
rect 14998 5629 15050 5635
rect 15010 800 15038 5629
rect 15190 3689 15242 3695
rect 15190 3631 15242 3637
rect 15202 800 15230 3631
rect 15298 800 15326 7405
rect 15490 6433 15518 15471
rect 15874 15165 15902 15841
rect 15862 15159 15914 15165
rect 15862 15101 15914 15107
rect 16150 10497 16202 10503
rect 16150 10439 16202 10445
rect 16162 8431 16190 10439
rect 16150 8425 16202 8431
rect 16150 8367 16202 8373
rect 16054 8277 16106 8283
rect 16054 8219 16106 8225
rect 15766 8129 15818 8135
rect 15766 8071 15818 8077
rect 15670 7463 15722 7469
rect 15670 7405 15722 7411
rect 15478 6427 15530 6433
rect 15478 6369 15530 6375
rect 15478 4355 15530 4361
rect 15478 4297 15530 4303
rect 15382 3911 15434 3917
rect 15382 3853 15434 3859
rect 15394 800 15422 3853
rect 15490 800 15518 4297
rect 15682 800 15710 7405
rect 15778 7099 15806 8071
rect 15766 7093 15818 7099
rect 15766 7035 15818 7041
rect 15862 5687 15914 5693
rect 15862 5629 15914 5635
rect 15766 4799 15818 4805
rect 15766 4741 15818 4747
rect 15778 4583 15806 4741
rect 15766 4577 15818 4583
rect 15766 4519 15818 4525
rect 15874 2894 15902 5629
rect 15958 4355 16010 4361
rect 15958 4297 16010 4303
rect 15778 2866 15902 2894
rect 15778 800 15806 2866
rect 15970 2160 15998 4297
rect 15874 2132 15998 2160
rect 15874 800 15902 2132
rect 16066 800 16094 8219
rect 16258 7765 16286 17266
rect 16342 8277 16394 8283
rect 16342 8219 16394 8225
rect 16246 7759 16298 7765
rect 16246 7701 16298 7707
rect 16150 5687 16202 5693
rect 16150 5629 16202 5635
rect 16162 800 16190 5629
rect 16246 4207 16298 4213
rect 16246 4149 16298 4155
rect 16258 800 16286 4149
rect 16354 800 16382 8219
rect 16450 6433 16478 37375
rect 16534 16935 16586 16941
rect 16534 16877 16586 16883
rect 16546 7099 16574 16877
rect 16834 9763 16862 56171
rect 17014 52825 17066 52831
rect 17014 52767 17066 52773
rect 16822 9757 16874 9763
rect 16822 9699 16874 9705
rect 17026 8431 17054 52767
rect 17782 34769 17834 34775
rect 17782 34711 17834 34717
rect 17794 34109 17822 34711
rect 17782 34103 17834 34109
rect 17782 34045 17834 34051
rect 17890 19457 17918 56689
rect 18070 56229 18122 56235
rect 18070 56171 18122 56177
rect 17974 42539 18026 42545
rect 17974 42481 18026 42487
rect 17878 19451 17930 19457
rect 17878 19393 17930 19399
rect 17986 14573 18014 42481
rect 18082 40325 18110 56171
rect 18178 56161 18206 57586
rect 18562 56531 18590 59200
rect 19138 57049 19166 59200
rect 19618 57614 19646 59200
rect 19618 57586 20030 57614
rect 19126 57043 19178 57049
rect 19126 56985 19178 56991
rect 19222 56747 19274 56753
rect 19222 56689 19274 56695
rect 18550 56525 18602 56531
rect 18550 56467 18602 56473
rect 18166 56155 18218 56161
rect 18166 56097 18218 56103
rect 18070 40319 18122 40325
rect 18070 40261 18122 40267
rect 19126 34917 19178 34923
rect 19126 34859 19178 34865
rect 18838 30847 18890 30853
rect 18838 30789 18890 30795
rect 18550 15455 18602 15461
rect 18550 15397 18602 15403
rect 18070 15233 18122 15239
rect 18070 15175 18122 15181
rect 17974 14567 18026 14573
rect 17974 14509 18026 14515
rect 17974 13679 18026 13685
rect 17974 13621 18026 13627
rect 17590 11015 17642 11021
rect 17590 10957 17642 10963
rect 17302 10201 17354 10207
rect 17302 10143 17354 10149
rect 17014 8425 17066 8431
rect 17014 8367 17066 8373
rect 17110 7167 17162 7173
rect 17110 7109 17162 7115
rect 16534 7093 16586 7099
rect 16534 7035 16586 7041
rect 16438 6427 16490 6433
rect 16438 6369 16490 6375
rect 16534 6353 16586 6359
rect 16534 6295 16586 6301
rect 16438 5021 16490 5027
rect 16438 4963 16490 4969
rect 16450 3917 16478 4963
rect 16438 3911 16490 3917
rect 16438 3853 16490 3859
rect 16546 800 16574 6295
rect 16726 6131 16778 6137
rect 16726 6073 16778 6079
rect 16630 3023 16682 3029
rect 16630 2965 16682 2971
rect 16642 800 16670 2965
rect 16738 800 16766 6073
rect 16918 4133 16970 4139
rect 16918 4075 16970 4081
rect 16930 800 16958 4075
rect 17014 3023 17066 3029
rect 17014 2965 17066 2971
rect 17026 800 17054 2965
rect 17122 800 17150 7109
rect 17314 6951 17342 10143
rect 17302 6945 17354 6951
rect 17302 6887 17354 6893
rect 17494 6205 17546 6211
rect 17494 6147 17546 6153
rect 17302 5021 17354 5027
rect 17302 4963 17354 4969
rect 17314 2894 17342 4963
rect 17398 3689 17450 3695
rect 17398 3631 17450 3637
rect 17218 2866 17342 2894
rect 17218 800 17246 2866
rect 17410 800 17438 3631
rect 17506 800 17534 6147
rect 17602 5120 17630 10957
rect 17782 10867 17834 10873
rect 17782 10809 17834 10815
rect 17686 6279 17738 6285
rect 17686 6221 17738 6227
rect 17698 5545 17726 6221
rect 17686 5539 17738 5545
rect 17686 5481 17738 5487
rect 17602 5092 17726 5120
rect 17590 5021 17642 5027
rect 17590 4963 17642 4969
rect 17602 800 17630 4963
rect 17698 3196 17726 5092
rect 17794 3769 17822 10809
rect 17986 7913 18014 13621
rect 17974 7907 18026 7913
rect 17974 7849 18026 7855
rect 18082 7099 18110 15175
rect 18454 10127 18506 10133
rect 18454 10069 18506 10075
rect 18358 7611 18410 7617
rect 18358 7553 18410 7559
rect 18070 7093 18122 7099
rect 18070 7035 18122 7041
rect 17878 6945 17930 6951
rect 17878 6887 17930 6893
rect 17782 3763 17834 3769
rect 17782 3705 17834 3711
rect 17698 3168 17822 3196
rect 17794 2955 17822 3168
rect 17782 2949 17834 2955
rect 17782 2891 17834 2897
rect 17686 2875 17738 2881
rect 17686 2817 17738 2823
rect 17698 800 17726 2817
rect 17890 800 17918 6887
rect 18070 6279 18122 6285
rect 18070 6221 18122 6227
rect 17974 5687 18026 5693
rect 17974 5629 18026 5635
rect 17986 800 18014 5629
rect 18082 2012 18110 6221
rect 18370 5249 18398 7553
rect 18466 6433 18494 10069
rect 18454 6427 18506 6433
rect 18454 6369 18506 6375
rect 18358 5243 18410 5249
rect 18358 5185 18410 5191
rect 18262 4133 18314 4139
rect 18262 4075 18314 4081
rect 18274 3843 18302 4075
rect 18358 3911 18410 3917
rect 18358 3853 18410 3859
rect 18262 3837 18314 3843
rect 18262 3779 18314 3785
rect 18262 3689 18314 3695
rect 18262 3631 18314 3637
rect 18082 1984 18206 2012
rect 18070 1913 18122 1919
rect 18070 1855 18122 1861
rect 18082 800 18110 1855
rect 18178 1716 18206 1984
rect 18274 1919 18302 3631
rect 18262 1913 18314 1919
rect 18262 1855 18314 1861
rect 18178 1688 18302 1716
rect 18274 800 18302 1688
rect 18370 800 18398 3853
rect 18562 3769 18590 15397
rect 18850 7099 18878 30789
rect 19030 16565 19082 16571
rect 19030 16507 19082 16513
rect 18934 15603 18986 15609
rect 18934 15545 18986 15551
rect 18838 7093 18890 7099
rect 18838 7035 18890 7041
rect 18646 6945 18698 6951
rect 18646 6887 18698 6893
rect 18550 3763 18602 3769
rect 18550 3705 18602 3711
rect 18454 3615 18506 3621
rect 18454 3557 18506 3563
rect 18466 800 18494 3557
rect 18658 2894 18686 6887
rect 18742 5687 18794 5693
rect 18742 5629 18794 5635
rect 18562 2866 18686 2894
rect 18562 800 18590 2866
rect 18754 800 18782 5629
rect 18838 4355 18890 4361
rect 18838 4297 18890 4303
rect 18850 800 18878 4297
rect 18946 3103 18974 15545
rect 19042 6581 19070 16507
rect 19030 6575 19082 6581
rect 19030 6517 19082 6523
rect 19042 6433 19070 6517
rect 19030 6427 19082 6433
rect 19030 6369 19082 6375
rect 19030 5021 19082 5027
rect 19030 4963 19082 4969
rect 19042 3917 19070 4963
rect 19138 4583 19166 34859
rect 19234 19827 19262 56689
rect 19628 56638 19924 56658
rect 19684 56636 19708 56638
rect 19764 56636 19788 56638
rect 19844 56636 19868 56638
rect 19706 56584 19708 56636
rect 19770 56584 19782 56636
rect 19844 56584 19846 56636
rect 19684 56582 19708 56584
rect 19764 56582 19788 56584
rect 19844 56582 19868 56584
rect 19628 56562 19924 56582
rect 20002 56531 20030 57586
rect 19990 56525 20042 56531
rect 19990 56467 20042 56473
rect 20194 55717 20222 59200
rect 20674 56975 20702 59200
rect 20662 56969 20714 56975
rect 20662 56911 20714 56917
rect 20854 56895 20906 56901
rect 20854 56837 20906 56843
rect 20374 56229 20426 56235
rect 20374 56171 20426 56177
rect 20182 55711 20234 55717
rect 20182 55653 20234 55659
rect 19628 55306 19924 55326
rect 19684 55304 19708 55306
rect 19764 55304 19788 55306
rect 19844 55304 19868 55306
rect 19706 55252 19708 55304
rect 19770 55252 19782 55304
rect 19844 55252 19846 55304
rect 19684 55250 19708 55252
rect 19764 55250 19788 55252
rect 19844 55250 19868 55252
rect 19628 55230 19924 55250
rect 19628 53974 19924 53994
rect 19684 53972 19708 53974
rect 19764 53972 19788 53974
rect 19844 53972 19868 53974
rect 19706 53920 19708 53972
rect 19770 53920 19782 53972
rect 19844 53920 19846 53972
rect 19684 53918 19708 53920
rect 19764 53918 19788 53920
rect 19844 53918 19868 53920
rect 19628 53898 19924 53918
rect 19628 52642 19924 52662
rect 19684 52640 19708 52642
rect 19764 52640 19788 52642
rect 19844 52640 19868 52642
rect 19706 52588 19708 52640
rect 19770 52588 19782 52640
rect 19844 52588 19846 52640
rect 19684 52586 19708 52588
rect 19764 52586 19788 52588
rect 19844 52586 19868 52588
rect 19628 52566 19924 52586
rect 19628 51310 19924 51330
rect 19684 51308 19708 51310
rect 19764 51308 19788 51310
rect 19844 51308 19868 51310
rect 19706 51256 19708 51308
rect 19770 51256 19782 51308
rect 19844 51256 19846 51308
rect 19684 51254 19708 51256
rect 19764 51254 19788 51256
rect 19844 51254 19868 51256
rect 19628 51234 19924 51254
rect 19628 49978 19924 49998
rect 19684 49976 19708 49978
rect 19764 49976 19788 49978
rect 19844 49976 19868 49978
rect 19706 49924 19708 49976
rect 19770 49924 19782 49976
rect 19844 49924 19846 49976
rect 19684 49922 19708 49924
rect 19764 49922 19788 49924
rect 19844 49922 19868 49924
rect 19628 49902 19924 49922
rect 19628 48646 19924 48666
rect 19684 48644 19708 48646
rect 19764 48644 19788 48646
rect 19844 48644 19868 48646
rect 19706 48592 19708 48644
rect 19770 48592 19782 48644
rect 19844 48592 19846 48644
rect 19684 48590 19708 48592
rect 19764 48590 19788 48592
rect 19844 48590 19868 48592
rect 19628 48570 19924 48590
rect 19628 47314 19924 47334
rect 19684 47312 19708 47314
rect 19764 47312 19788 47314
rect 19844 47312 19868 47314
rect 19706 47260 19708 47312
rect 19770 47260 19782 47312
rect 19844 47260 19846 47312
rect 19684 47258 19708 47260
rect 19764 47258 19788 47260
rect 19844 47258 19868 47260
rect 19628 47238 19924 47258
rect 19628 45982 19924 46002
rect 19684 45980 19708 45982
rect 19764 45980 19788 45982
rect 19844 45980 19868 45982
rect 19706 45928 19708 45980
rect 19770 45928 19782 45980
rect 19844 45928 19846 45980
rect 19684 45926 19708 45928
rect 19764 45926 19788 45928
rect 19844 45926 19868 45928
rect 19628 45906 19924 45926
rect 19628 44650 19924 44670
rect 19684 44648 19708 44650
rect 19764 44648 19788 44650
rect 19844 44648 19868 44650
rect 19706 44596 19708 44648
rect 19770 44596 19782 44648
rect 19844 44596 19846 44648
rect 19684 44594 19708 44596
rect 19764 44594 19788 44596
rect 19844 44594 19868 44596
rect 19628 44574 19924 44594
rect 19628 43318 19924 43338
rect 19684 43316 19708 43318
rect 19764 43316 19788 43318
rect 19844 43316 19868 43318
rect 19706 43264 19708 43316
rect 19770 43264 19782 43316
rect 19844 43264 19846 43316
rect 19684 43262 19708 43264
rect 19764 43262 19788 43264
rect 19844 43262 19868 43264
rect 19628 43242 19924 43262
rect 19628 41986 19924 42006
rect 19684 41984 19708 41986
rect 19764 41984 19788 41986
rect 19844 41984 19868 41986
rect 19706 41932 19708 41984
rect 19770 41932 19782 41984
rect 19844 41932 19846 41984
rect 19684 41930 19708 41932
rect 19764 41930 19788 41932
rect 19844 41930 19868 41932
rect 19628 41910 19924 41930
rect 19628 40654 19924 40674
rect 19684 40652 19708 40654
rect 19764 40652 19788 40654
rect 19844 40652 19868 40654
rect 19706 40600 19708 40652
rect 19770 40600 19782 40652
rect 19844 40600 19846 40652
rect 19684 40598 19708 40600
rect 19764 40598 19788 40600
rect 19844 40598 19868 40600
rect 19628 40578 19924 40598
rect 19628 39322 19924 39342
rect 19684 39320 19708 39322
rect 19764 39320 19788 39322
rect 19844 39320 19868 39322
rect 19706 39268 19708 39320
rect 19770 39268 19782 39320
rect 19844 39268 19846 39320
rect 19684 39266 19708 39268
rect 19764 39266 19788 39268
rect 19844 39266 19868 39268
rect 19628 39246 19924 39266
rect 19628 37990 19924 38010
rect 19684 37988 19708 37990
rect 19764 37988 19788 37990
rect 19844 37988 19868 37990
rect 19706 37936 19708 37988
rect 19770 37936 19782 37988
rect 19844 37936 19846 37988
rect 19684 37934 19708 37936
rect 19764 37934 19788 37936
rect 19844 37934 19868 37936
rect 19628 37914 19924 37934
rect 19628 36658 19924 36678
rect 19684 36656 19708 36658
rect 19764 36656 19788 36658
rect 19844 36656 19868 36658
rect 19706 36604 19708 36656
rect 19770 36604 19782 36656
rect 19844 36604 19846 36656
rect 19684 36602 19708 36604
rect 19764 36602 19788 36604
rect 19844 36602 19868 36604
rect 19628 36582 19924 36602
rect 20386 36255 20414 56171
rect 20470 55563 20522 55569
rect 20470 55505 20522 55511
rect 20482 46319 20510 55505
rect 20470 46313 20522 46319
rect 20470 46255 20522 46261
rect 20374 36249 20426 36255
rect 20374 36191 20426 36197
rect 20470 35583 20522 35589
rect 20470 35525 20522 35531
rect 19628 35326 19924 35346
rect 19684 35324 19708 35326
rect 19764 35324 19788 35326
rect 19844 35324 19868 35326
rect 19706 35272 19708 35324
rect 19770 35272 19782 35324
rect 19844 35272 19846 35324
rect 19684 35270 19708 35272
rect 19764 35270 19788 35272
rect 19844 35270 19868 35272
rect 19628 35250 19924 35270
rect 19990 34843 20042 34849
rect 19990 34785 20042 34791
rect 19628 33994 19924 34014
rect 19684 33992 19708 33994
rect 19764 33992 19788 33994
rect 19844 33992 19868 33994
rect 19706 33940 19708 33992
rect 19770 33940 19782 33992
rect 19844 33940 19846 33992
rect 19684 33938 19708 33940
rect 19764 33938 19788 33940
rect 19844 33938 19868 33940
rect 19628 33918 19924 33938
rect 19628 32662 19924 32682
rect 19684 32660 19708 32662
rect 19764 32660 19788 32662
rect 19844 32660 19868 32662
rect 19706 32608 19708 32660
rect 19770 32608 19782 32660
rect 19844 32608 19846 32660
rect 19684 32606 19708 32608
rect 19764 32606 19788 32608
rect 19844 32606 19868 32608
rect 19628 32586 19924 32606
rect 19628 31330 19924 31350
rect 19684 31328 19708 31330
rect 19764 31328 19788 31330
rect 19844 31328 19868 31330
rect 19706 31276 19708 31328
rect 19770 31276 19782 31328
rect 19844 31276 19846 31328
rect 19684 31274 19708 31276
rect 19764 31274 19788 31276
rect 19844 31274 19868 31276
rect 19628 31254 19924 31274
rect 19628 29998 19924 30018
rect 19684 29996 19708 29998
rect 19764 29996 19788 29998
rect 19844 29996 19868 29998
rect 19706 29944 19708 29996
rect 19770 29944 19782 29996
rect 19844 29944 19846 29996
rect 19684 29942 19708 29944
rect 19764 29942 19788 29944
rect 19844 29942 19868 29944
rect 19628 29922 19924 29942
rect 19628 28666 19924 28686
rect 19684 28664 19708 28666
rect 19764 28664 19788 28666
rect 19844 28664 19868 28666
rect 19706 28612 19708 28664
rect 19770 28612 19782 28664
rect 19844 28612 19846 28664
rect 19684 28610 19708 28612
rect 19764 28610 19788 28612
rect 19844 28610 19868 28612
rect 19628 28590 19924 28610
rect 19628 27334 19924 27354
rect 19684 27332 19708 27334
rect 19764 27332 19788 27334
rect 19844 27332 19868 27334
rect 19706 27280 19708 27332
rect 19770 27280 19782 27332
rect 19844 27280 19846 27332
rect 19684 27278 19708 27280
rect 19764 27278 19788 27280
rect 19844 27278 19868 27280
rect 19628 27258 19924 27278
rect 19628 26002 19924 26022
rect 19684 26000 19708 26002
rect 19764 26000 19788 26002
rect 19844 26000 19868 26002
rect 19706 25948 19708 26000
rect 19770 25948 19782 26000
rect 19844 25948 19846 26000
rect 19684 25946 19708 25948
rect 19764 25946 19788 25948
rect 19844 25946 19868 25948
rect 19628 25926 19924 25946
rect 19628 24670 19924 24690
rect 19684 24668 19708 24670
rect 19764 24668 19788 24670
rect 19844 24668 19868 24670
rect 19706 24616 19708 24668
rect 19770 24616 19782 24668
rect 19844 24616 19846 24668
rect 19684 24614 19708 24616
rect 19764 24614 19788 24616
rect 19844 24614 19868 24616
rect 19628 24594 19924 24614
rect 19628 23338 19924 23358
rect 19684 23336 19708 23338
rect 19764 23336 19788 23338
rect 19844 23336 19868 23338
rect 19706 23284 19708 23336
rect 19770 23284 19782 23336
rect 19844 23284 19846 23336
rect 19684 23282 19708 23284
rect 19764 23282 19788 23284
rect 19844 23282 19868 23284
rect 19628 23262 19924 23282
rect 19414 22781 19466 22787
rect 19414 22723 19466 22729
rect 19222 19821 19274 19827
rect 19222 19763 19274 19769
rect 19426 10133 19454 22723
rect 19628 22006 19924 22026
rect 19684 22004 19708 22006
rect 19764 22004 19788 22006
rect 19844 22004 19868 22006
rect 19706 21952 19708 22004
rect 19770 21952 19782 22004
rect 19844 21952 19846 22004
rect 19684 21950 19708 21952
rect 19764 21950 19788 21952
rect 19844 21950 19868 21952
rect 19628 21930 19924 21950
rect 19628 20674 19924 20694
rect 19684 20672 19708 20674
rect 19764 20672 19788 20674
rect 19844 20672 19868 20674
rect 19706 20620 19708 20672
rect 19770 20620 19782 20672
rect 19844 20620 19846 20672
rect 19684 20618 19708 20620
rect 19764 20618 19788 20620
rect 19844 20618 19868 20620
rect 19628 20598 19924 20618
rect 19628 19342 19924 19362
rect 19684 19340 19708 19342
rect 19764 19340 19788 19342
rect 19844 19340 19868 19342
rect 19706 19288 19708 19340
rect 19770 19288 19782 19340
rect 19844 19288 19846 19340
rect 19684 19286 19708 19288
rect 19764 19286 19788 19288
rect 19844 19286 19868 19288
rect 19628 19266 19924 19286
rect 19628 18010 19924 18030
rect 19684 18008 19708 18010
rect 19764 18008 19788 18010
rect 19844 18008 19868 18010
rect 19706 17956 19708 18008
rect 19770 17956 19782 18008
rect 19844 17956 19846 18008
rect 19684 17954 19708 17956
rect 19764 17954 19788 17956
rect 19844 17954 19868 17956
rect 19628 17934 19924 17954
rect 19628 16678 19924 16698
rect 19684 16676 19708 16678
rect 19764 16676 19788 16678
rect 19844 16676 19868 16678
rect 19706 16624 19708 16676
rect 19770 16624 19782 16676
rect 19844 16624 19846 16676
rect 19684 16622 19708 16624
rect 19764 16622 19788 16624
rect 19844 16622 19868 16624
rect 19628 16602 19924 16622
rect 19628 15346 19924 15366
rect 19684 15344 19708 15346
rect 19764 15344 19788 15346
rect 19844 15344 19868 15346
rect 19706 15292 19708 15344
rect 19770 15292 19782 15344
rect 19844 15292 19846 15344
rect 19684 15290 19708 15292
rect 19764 15290 19788 15292
rect 19844 15290 19868 15292
rect 19628 15270 19924 15290
rect 19628 14014 19924 14034
rect 19684 14012 19708 14014
rect 19764 14012 19788 14014
rect 19844 14012 19868 14014
rect 19706 13960 19708 14012
rect 19770 13960 19782 14012
rect 19844 13960 19846 14012
rect 19684 13958 19708 13960
rect 19764 13958 19788 13960
rect 19844 13958 19868 13960
rect 19628 13938 19924 13958
rect 19628 12682 19924 12702
rect 19684 12680 19708 12682
rect 19764 12680 19788 12682
rect 19844 12680 19868 12682
rect 19706 12628 19708 12680
rect 19770 12628 19782 12680
rect 19844 12628 19846 12680
rect 19684 12626 19708 12628
rect 19764 12626 19788 12628
rect 19844 12626 19868 12628
rect 19628 12606 19924 12626
rect 19628 11350 19924 11370
rect 19684 11348 19708 11350
rect 19764 11348 19788 11350
rect 19844 11348 19868 11350
rect 19706 11296 19708 11348
rect 19770 11296 19782 11348
rect 19844 11296 19846 11348
rect 19684 11294 19708 11296
rect 19764 11294 19788 11296
rect 19844 11294 19868 11296
rect 19628 11274 19924 11294
rect 19414 10127 19466 10133
rect 19414 10069 19466 10075
rect 19628 10018 19924 10038
rect 19684 10016 19708 10018
rect 19764 10016 19788 10018
rect 19844 10016 19868 10018
rect 19706 9964 19708 10016
rect 19770 9964 19782 10016
rect 19844 9964 19846 10016
rect 19684 9962 19708 9964
rect 19764 9962 19788 9964
rect 19844 9962 19868 9964
rect 19628 9942 19924 9962
rect 19628 8686 19924 8706
rect 19684 8684 19708 8686
rect 19764 8684 19788 8686
rect 19844 8684 19868 8686
rect 19706 8632 19708 8684
rect 19770 8632 19782 8684
rect 19844 8632 19846 8684
rect 19684 8630 19708 8632
rect 19764 8630 19788 8632
rect 19844 8630 19868 8632
rect 19628 8610 19924 8630
rect 19628 7354 19924 7374
rect 19684 7352 19708 7354
rect 19764 7352 19788 7354
rect 19844 7352 19868 7354
rect 19706 7300 19708 7352
rect 19770 7300 19782 7352
rect 19844 7300 19846 7352
rect 19684 7298 19708 7300
rect 19764 7298 19788 7300
rect 19844 7298 19868 7300
rect 19628 7278 19924 7298
rect 20002 6433 20030 34785
rect 20374 34769 20426 34775
rect 20374 34711 20426 34717
rect 20386 7099 20414 34711
rect 20482 9023 20510 35525
rect 20866 19753 20894 56837
rect 21250 56531 21278 59200
rect 21622 56895 21674 56901
rect 21622 56837 21674 56843
rect 21238 56525 21290 56531
rect 21238 56467 21290 56473
rect 21430 56229 21482 56235
rect 21430 56171 21482 56177
rect 21442 51203 21470 56171
rect 21430 51197 21482 51203
rect 21430 51139 21482 51145
rect 21634 47534 21662 56837
rect 21730 56531 21758 59200
rect 22306 56975 22334 59200
rect 22294 56969 22346 56975
rect 22294 56911 22346 56917
rect 21814 56747 21866 56753
rect 21814 56689 21866 56695
rect 22006 56747 22058 56753
rect 22006 56689 22058 56695
rect 21718 56525 21770 56531
rect 21718 56467 21770 56473
rect 21826 56161 21854 56689
rect 21814 56155 21866 56161
rect 21814 56097 21866 56103
rect 22018 48484 22046 56689
rect 22786 56531 22814 59200
rect 22774 56525 22826 56531
rect 22774 56467 22826 56473
rect 22870 56303 22922 56309
rect 22870 56245 22922 56251
rect 22102 56229 22154 56235
rect 22102 56171 22154 56177
rect 22678 56229 22730 56235
rect 22678 56171 22730 56177
rect 21970 48465 22046 48484
rect 21958 48459 22046 48465
rect 22010 48456 22046 48459
rect 21958 48401 22010 48407
rect 22114 47534 22142 56171
rect 22198 52085 22250 52091
rect 22198 52027 22250 52033
rect 21634 47506 21758 47534
rect 21334 38765 21386 38771
rect 21334 38707 21386 38713
rect 20854 19747 20906 19753
rect 20854 19689 20906 19695
rect 20758 17823 20810 17829
rect 20758 17765 20810 17771
rect 20770 17294 20798 17765
rect 20770 17266 20894 17294
rect 20866 12974 20894 17266
rect 20866 12946 20990 12974
rect 20662 10349 20714 10355
rect 20662 10291 20714 10297
rect 20470 9017 20522 9023
rect 20470 8959 20522 8965
rect 20374 7093 20426 7099
rect 20374 7035 20426 7041
rect 20374 6945 20426 6951
rect 20374 6887 20426 6893
rect 19990 6427 20042 6433
rect 19990 6369 20042 6375
rect 19318 6131 19370 6137
rect 19318 6073 19370 6079
rect 19990 6131 20042 6137
rect 19990 6073 20042 6079
rect 19222 5021 19274 5027
rect 19222 4963 19274 4969
rect 19126 4577 19178 4583
rect 19126 4519 19178 4525
rect 19030 3911 19082 3917
rect 19030 3853 19082 3859
rect 18934 3097 18986 3103
rect 18934 3039 18986 3045
rect 18934 2875 18986 2881
rect 18934 2817 18986 2823
rect 18946 800 18974 2817
rect 19234 2604 19262 4963
rect 19330 2955 19358 6073
rect 19628 6022 19924 6042
rect 19684 6020 19708 6022
rect 19764 6020 19788 6022
rect 19844 6020 19868 6022
rect 19706 5968 19708 6020
rect 19770 5968 19782 6020
rect 19844 5968 19846 6020
rect 19684 5966 19708 5968
rect 19764 5966 19788 5968
rect 19844 5966 19868 5968
rect 19628 5946 19924 5966
rect 19628 4690 19924 4710
rect 19684 4688 19708 4690
rect 19764 4688 19788 4690
rect 19844 4688 19868 4690
rect 19706 4636 19708 4688
rect 19770 4636 19782 4688
rect 19844 4636 19846 4688
rect 19684 4634 19708 4636
rect 19764 4634 19788 4636
rect 19844 4634 19868 4636
rect 19628 4614 19924 4634
rect 19510 4281 19562 4287
rect 19510 4223 19562 4229
rect 19414 3763 19466 3769
rect 19414 3705 19466 3711
rect 19318 2949 19370 2955
rect 19318 2891 19370 2897
rect 19318 2801 19370 2807
rect 19318 2743 19370 2749
rect 19042 2576 19262 2604
rect 19042 800 19070 2576
rect 19330 1568 19358 2743
rect 19234 1540 19358 1568
rect 19234 800 19262 1540
rect 19318 1469 19370 1475
rect 19318 1411 19370 1417
rect 19330 800 19358 1411
rect 19426 800 19454 3705
rect 19522 2012 19550 4223
rect 19892 3506 19948 3515
rect 19892 3441 19894 3450
rect 19946 3441 19948 3450
rect 19894 3409 19946 3415
rect 19628 3358 19924 3378
rect 19684 3356 19708 3358
rect 19764 3356 19788 3358
rect 19844 3356 19868 3358
rect 19706 3304 19708 3356
rect 19770 3304 19782 3356
rect 19844 3304 19846 3356
rect 19684 3302 19708 3304
rect 19764 3302 19788 3304
rect 19844 3302 19868 3304
rect 19628 3282 19924 3302
rect 19702 3245 19754 3251
rect 19702 3187 19754 3193
rect 19796 3210 19852 3219
rect 19522 1984 19646 2012
rect 19618 800 19646 1984
rect 19714 800 19742 3187
rect 19796 3145 19852 3154
rect 19810 800 19838 3145
rect 19894 2801 19946 2807
rect 19894 2743 19946 2749
rect 19906 800 19934 2743
rect 20002 1475 20030 6073
rect 20182 5687 20234 5693
rect 20182 5629 20234 5635
rect 20086 4207 20138 4213
rect 20086 4149 20138 4155
rect 19990 1469 20042 1475
rect 19990 1411 20042 1417
rect 20098 800 20126 4149
rect 20194 3473 20222 5629
rect 20278 3689 20330 3695
rect 20278 3631 20330 3637
rect 20182 3467 20234 3473
rect 20182 3409 20234 3415
rect 20182 2579 20234 2585
rect 20182 2521 20234 2527
rect 20194 800 20222 2521
rect 20290 800 20318 3631
rect 20386 3251 20414 6887
rect 20470 5687 20522 5693
rect 20470 5629 20522 5635
rect 20374 3245 20426 3251
rect 20374 3187 20426 3193
rect 20482 1716 20510 5629
rect 20566 5021 20618 5027
rect 20566 4963 20618 4969
rect 20578 3769 20606 4963
rect 20566 3763 20618 3769
rect 20566 3705 20618 3711
rect 20566 3615 20618 3621
rect 20566 3557 20618 3563
rect 20578 1864 20606 3557
rect 20674 2955 20702 10291
rect 20758 7463 20810 7469
rect 20758 7405 20810 7411
rect 20662 2949 20714 2955
rect 20662 2891 20714 2897
rect 20578 1836 20702 1864
rect 20482 1688 20606 1716
rect 20470 1617 20522 1623
rect 20470 1559 20522 1565
rect 20482 800 20510 1559
rect 20578 800 20606 1688
rect 20674 800 20702 1836
rect 20770 800 20798 7405
rect 20854 6945 20906 6951
rect 20854 6887 20906 6893
rect 20866 1623 20894 6887
rect 20962 6433 20990 12946
rect 21046 10127 21098 10133
rect 21046 10069 21098 10075
rect 21058 7765 21086 10069
rect 21346 8357 21374 38707
rect 21622 35139 21674 35145
rect 21622 35081 21674 35087
rect 21526 11237 21578 11243
rect 21526 11179 21578 11185
rect 21334 8351 21386 8357
rect 21334 8293 21386 8299
rect 21046 7759 21098 7765
rect 21046 7701 21098 7707
rect 21238 6945 21290 6951
rect 21154 6905 21238 6933
rect 20950 6427 21002 6433
rect 20950 6369 21002 6375
rect 21046 4355 21098 4361
rect 21046 4297 21098 4303
rect 20950 4281 21002 4287
rect 20950 4223 21002 4229
rect 20854 1617 20906 1623
rect 20854 1559 20906 1565
rect 20962 800 20990 4223
rect 21058 800 21086 4297
rect 21154 800 21182 6905
rect 21238 6887 21290 6893
rect 21538 6433 21566 11179
rect 21526 6427 21578 6433
rect 21526 6369 21578 6375
rect 21430 6131 21482 6137
rect 21430 6073 21482 6079
rect 21238 5021 21290 5027
rect 21238 4963 21290 4969
rect 21250 2585 21278 4963
rect 21442 4213 21470 6073
rect 21430 4207 21482 4213
rect 21430 4149 21482 4155
rect 21526 4207 21578 4213
rect 21526 4149 21578 4155
rect 21334 3911 21386 3917
rect 21334 3853 21386 3859
rect 21238 2579 21290 2585
rect 21238 2521 21290 2527
rect 21346 2456 21374 3853
rect 21430 2949 21482 2955
rect 21430 2891 21482 2897
rect 21250 2428 21374 2456
rect 21250 800 21278 2428
rect 21442 800 21470 2891
rect 21538 800 21566 4149
rect 21634 3251 21662 35081
rect 21730 16127 21758 47506
rect 22018 47506 22142 47534
rect 22210 47534 22238 52027
rect 22210 47506 22334 47534
rect 22018 37454 22046 47506
rect 22018 37426 22142 37454
rect 22114 25525 22142 37426
rect 22102 25519 22154 25525
rect 22102 25461 22154 25467
rect 21718 16121 21770 16127
rect 21718 16063 21770 16069
rect 21910 13087 21962 13093
rect 21910 13029 21962 13035
rect 21922 7099 21950 13029
rect 22306 7173 22334 47506
rect 22690 35737 22718 56171
rect 22882 48539 22910 56245
rect 23362 55717 23390 59200
rect 23842 56975 23870 59200
rect 23830 56969 23882 56975
rect 23830 56911 23882 56917
rect 24418 56531 24446 59200
rect 24406 56525 24458 56531
rect 24406 56467 24458 56473
rect 24406 56229 24458 56235
rect 24406 56171 24458 56177
rect 23350 55711 23402 55717
rect 23350 55653 23402 55659
rect 23158 55415 23210 55421
rect 23158 55357 23210 55363
rect 22966 49495 23018 49501
rect 22966 49437 23018 49443
rect 22870 48533 22922 48539
rect 22870 48475 22922 48481
rect 22678 35731 22730 35737
rect 22678 35673 22730 35679
rect 22870 22263 22922 22269
rect 22870 22205 22922 22211
rect 22882 19457 22910 22205
rect 22870 19451 22922 19457
rect 22870 19393 22922 19399
rect 22486 15677 22538 15683
rect 22486 15619 22538 15625
rect 22498 12974 22526 15619
rect 22402 12946 22526 12974
rect 22294 7167 22346 7173
rect 22294 7109 22346 7115
rect 21910 7093 21962 7099
rect 21910 7035 21962 7041
rect 21910 6945 21962 6951
rect 21910 6887 21962 6893
rect 21718 5687 21770 5693
rect 21718 5629 21770 5635
rect 21730 4287 21758 5629
rect 21814 4355 21866 4361
rect 21814 4297 21866 4303
rect 21718 4281 21770 4287
rect 21718 4223 21770 4229
rect 21718 3541 21770 3547
rect 21718 3483 21770 3489
rect 21730 3251 21758 3483
rect 21622 3245 21674 3251
rect 21622 3187 21674 3193
rect 21718 3245 21770 3251
rect 21718 3187 21770 3193
rect 21622 3097 21674 3103
rect 21622 3039 21674 3045
rect 21634 800 21662 3039
rect 21826 800 21854 4297
rect 21922 800 21950 6887
rect 22294 6205 22346 6211
rect 22294 6147 22346 6153
rect 22102 3763 22154 3769
rect 22102 3705 22154 3711
rect 22114 2308 22142 3705
rect 22018 2280 22142 2308
rect 22018 800 22046 2280
rect 22102 1617 22154 1623
rect 22102 1559 22154 1565
rect 22114 800 22142 1559
rect 22306 800 22334 6147
rect 22402 3843 22430 12946
rect 22978 6433 23006 49437
rect 23062 49421 23114 49427
rect 23062 49363 23114 49369
rect 23074 7839 23102 49363
rect 23170 20123 23198 55357
rect 23254 51567 23306 51573
rect 23254 51509 23306 51515
rect 23158 20117 23210 20123
rect 23158 20059 23210 20065
rect 23266 17829 23294 51509
rect 24418 46097 24446 56171
rect 24898 55717 24926 59200
rect 25474 56975 25502 59200
rect 25462 56969 25514 56975
rect 25462 56911 25514 56917
rect 25954 56531 25982 59200
rect 26530 56531 26558 59200
rect 27010 56975 27038 59200
rect 26998 56969 27050 56975
rect 26998 56911 27050 56917
rect 27286 56747 27338 56753
rect 27286 56689 27338 56695
rect 25942 56525 25994 56531
rect 25942 56467 25994 56473
rect 26518 56525 26570 56531
rect 26518 56467 26570 56473
rect 27298 56457 27326 56689
rect 27586 56531 27614 59200
rect 28066 56531 28094 59200
rect 28642 56975 28670 59200
rect 29122 57049 29150 59200
rect 29110 57043 29162 57049
rect 29110 56985 29162 56991
rect 28630 56969 28682 56975
rect 28630 56911 28682 56917
rect 29698 56531 29726 59200
rect 30178 56975 30206 59200
rect 30166 56969 30218 56975
rect 30166 56911 30218 56917
rect 30658 56531 30686 59200
rect 31234 56531 31262 59200
rect 31714 56975 31742 59200
rect 31702 56969 31754 56975
rect 31702 56911 31754 56917
rect 32290 56531 32318 59200
rect 32566 56895 32618 56901
rect 32566 56837 32618 56843
rect 32470 56821 32522 56827
rect 32470 56763 32522 56769
rect 27574 56525 27626 56531
rect 27574 56467 27626 56473
rect 28054 56525 28106 56531
rect 28054 56467 28106 56473
rect 29686 56525 29738 56531
rect 29686 56467 29738 56473
rect 30646 56525 30698 56531
rect 30646 56467 30698 56473
rect 31222 56525 31274 56531
rect 31222 56467 31274 56473
rect 32278 56525 32330 56531
rect 32278 56467 32330 56473
rect 32482 56457 32510 56763
rect 27286 56451 27338 56457
rect 27286 56393 27338 56399
rect 32470 56451 32522 56457
rect 32470 56393 32522 56399
rect 26134 56229 26186 56235
rect 26134 56171 26186 56177
rect 27766 56229 27818 56235
rect 27766 56171 27818 56177
rect 28438 56229 28490 56235
rect 28438 56171 28490 56177
rect 29590 56229 29642 56235
rect 29590 56171 29642 56177
rect 30934 56229 30986 56235
rect 30934 56171 30986 56177
rect 32470 56229 32522 56235
rect 32470 56171 32522 56177
rect 24886 55711 24938 55717
rect 24886 55653 24938 55659
rect 25078 55563 25130 55569
rect 25078 55505 25130 55511
rect 24406 46091 24458 46097
rect 24406 46033 24458 46039
rect 24694 38247 24746 38253
rect 24694 38189 24746 38195
rect 24502 20191 24554 20197
rect 24502 20133 24554 20139
rect 23254 17823 23306 17829
rect 23254 17765 23306 17771
rect 23158 17453 23210 17459
rect 23158 17395 23210 17401
rect 23062 7833 23114 7839
rect 23062 7775 23114 7781
rect 23170 7691 23198 17395
rect 24214 14197 24266 14203
rect 24214 14139 24266 14145
rect 23446 12939 23498 12945
rect 23446 12881 23498 12887
rect 23458 11835 23486 12881
rect 23446 11829 23498 11835
rect 23446 11771 23498 11777
rect 23542 11755 23594 11761
rect 23542 11697 23594 11703
rect 23554 11632 23582 11697
rect 23266 11604 23582 11632
rect 23266 11539 23294 11604
rect 23254 11533 23306 11539
rect 23254 11475 23306 11481
rect 23926 11089 23978 11095
rect 23926 11031 23978 11037
rect 23254 10941 23306 10947
rect 23254 10883 23306 10889
rect 23158 7685 23210 7691
rect 23158 7627 23210 7633
rect 23062 7167 23114 7173
rect 23062 7109 23114 7115
rect 23074 6803 23102 7109
rect 23062 6797 23114 6803
rect 23062 6739 23114 6745
rect 23266 6433 23294 10883
rect 23446 10127 23498 10133
rect 23446 10069 23498 10075
rect 23458 7099 23486 10069
rect 23938 7765 23966 11031
rect 23926 7759 23978 7765
rect 23926 7701 23978 7707
rect 23734 7463 23786 7469
rect 23734 7405 23786 7411
rect 23446 7093 23498 7099
rect 23446 7035 23498 7041
rect 23638 7019 23690 7025
rect 23638 6961 23690 6967
rect 22966 6427 23018 6433
rect 22966 6369 23018 6375
rect 23254 6427 23306 6433
rect 23254 6369 23306 6375
rect 22870 6131 22922 6137
rect 22870 6073 22922 6079
rect 22486 5687 22538 5693
rect 22486 5629 22538 5635
rect 22390 3837 22442 3843
rect 22390 3779 22442 3785
rect 22390 3171 22442 3177
rect 22390 3113 22442 3119
rect 22402 800 22430 3113
rect 22498 3103 22526 5629
rect 22774 5021 22826 5027
rect 22774 4963 22826 4969
rect 22786 3917 22814 4963
rect 22882 4213 22910 6073
rect 23350 5835 23402 5841
rect 23350 5777 23402 5783
rect 23062 5687 23114 5693
rect 23062 5629 23114 5635
rect 22870 4207 22922 4213
rect 22870 4149 22922 4155
rect 22774 3911 22826 3917
rect 22774 3853 22826 3859
rect 23074 3788 23102 5629
rect 23158 5021 23210 5027
rect 23158 4963 23210 4969
rect 22786 3760 23102 3788
rect 22678 3689 22730 3695
rect 22678 3631 22730 3637
rect 22582 3541 22634 3547
rect 22582 3483 22634 3489
rect 22486 3097 22538 3103
rect 22486 3039 22538 3045
rect 22486 2949 22538 2955
rect 22486 2891 22538 2897
rect 22498 800 22526 2891
rect 22594 800 22622 3483
rect 22690 1623 22718 3631
rect 22678 1617 22730 1623
rect 22678 1559 22730 1565
rect 22786 800 22814 3760
rect 22870 3689 22922 3695
rect 22870 3631 22922 3637
rect 22882 800 22910 3631
rect 22966 3615 23018 3621
rect 22966 3557 23018 3563
rect 22978 800 23006 3557
rect 23062 3467 23114 3473
rect 23062 3409 23114 3415
rect 23074 2604 23102 3409
rect 23170 3177 23198 4963
rect 23254 4355 23306 4361
rect 23254 4297 23306 4303
rect 23158 3171 23210 3177
rect 23158 3113 23210 3119
rect 23074 2576 23198 2604
rect 23170 800 23198 2576
rect 23266 800 23294 4297
rect 23362 800 23390 5777
rect 23446 5687 23498 5693
rect 23446 5629 23498 5635
rect 23458 800 23486 5629
rect 23650 3788 23678 6961
rect 23554 3760 23678 3788
rect 23554 3547 23582 3760
rect 23638 3689 23690 3695
rect 23638 3631 23690 3637
rect 23542 3541 23594 3547
rect 23542 3483 23594 3489
rect 23650 800 23678 3631
rect 23746 800 23774 7405
rect 24226 7099 24254 14139
rect 24214 7093 24266 7099
rect 24214 7035 24266 7041
rect 23926 6945 23978 6951
rect 23926 6887 23978 6893
rect 24118 6945 24170 6951
rect 24118 6887 24170 6893
rect 23938 6803 23966 6887
rect 23926 6797 23978 6803
rect 23926 6739 23978 6745
rect 24130 5841 24158 6887
rect 24514 6433 24542 20133
rect 24706 7765 24734 38189
rect 25090 21085 25118 55505
rect 25558 53565 25610 53571
rect 25558 53507 25610 53513
rect 25570 49871 25598 53507
rect 25846 50309 25898 50315
rect 25846 50251 25898 50257
rect 25558 49865 25610 49871
rect 25558 49807 25610 49813
rect 25858 49797 25886 50251
rect 25846 49791 25898 49797
rect 25846 49733 25898 49739
rect 26146 49205 26174 56171
rect 26614 53417 26666 53423
rect 26614 53359 26666 53365
rect 26134 49199 26186 49205
rect 26134 49141 26186 49147
rect 25174 39579 25226 39585
rect 25174 39521 25226 39527
rect 25078 21079 25130 21085
rect 25078 21021 25130 21027
rect 25186 11169 25214 39521
rect 25270 39505 25322 39511
rect 25270 39447 25322 39453
rect 25174 11163 25226 11169
rect 25174 11105 25226 11111
rect 25282 10429 25310 39447
rect 25366 36767 25418 36773
rect 25366 36709 25418 36715
rect 25378 11243 25406 36709
rect 26518 31735 26570 31741
rect 26518 31677 26570 31683
rect 25462 28923 25514 28929
rect 25462 28865 25514 28871
rect 25474 13167 25502 28865
rect 26530 26931 26558 31677
rect 26518 26925 26570 26931
rect 26518 26867 26570 26873
rect 25558 22263 25610 22269
rect 25558 22205 25610 22211
rect 25462 13161 25514 13167
rect 25462 13103 25514 13109
rect 25366 11237 25418 11243
rect 25366 11179 25418 11185
rect 25270 10423 25322 10429
rect 25270 10365 25322 10371
rect 25570 10133 25598 22205
rect 26626 21677 26654 53359
rect 27778 50167 27806 56171
rect 28342 55193 28394 55199
rect 28342 55135 28394 55141
rect 27766 50161 27818 50167
rect 27766 50103 27818 50109
rect 27958 47571 28010 47577
rect 27958 47513 28010 47519
rect 26710 43427 26762 43433
rect 26710 43369 26762 43375
rect 26614 21671 26666 21677
rect 26614 21613 26666 21619
rect 26230 20931 26282 20937
rect 26230 20873 26282 20879
rect 25654 19673 25706 19679
rect 25654 19615 25706 19621
rect 25558 10127 25610 10133
rect 25558 10069 25610 10075
rect 24694 7759 24746 7765
rect 24694 7701 24746 7707
rect 24598 7463 24650 7469
rect 24598 7405 24650 7411
rect 24790 7463 24842 7469
rect 24790 7405 24842 7411
rect 24502 6427 24554 6433
rect 24502 6369 24554 6375
rect 24310 6131 24362 6137
rect 24310 6073 24362 6079
rect 24118 5835 24170 5841
rect 24118 5777 24170 5783
rect 23830 5021 23882 5027
rect 23830 4963 23882 4969
rect 23842 3473 23870 4963
rect 23926 4577 23978 4583
rect 23926 4519 23978 4525
rect 23830 3467 23882 3473
rect 23830 3409 23882 3415
rect 23938 2604 23966 4519
rect 24022 4355 24074 4361
rect 24022 4297 24074 4303
rect 24034 3769 24062 4297
rect 24118 4207 24170 4213
rect 24118 4149 24170 4155
rect 24022 3763 24074 3769
rect 24022 3705 24074 3711
rect 24022 3023 24074 3029
rect 24022 2965 24074 2971
rect 23842 2576 23966 2604
rect 23842 800 23870 2576
rect 24034 800 24062 2965
rect 24130 800 24158 4149
rect 24214 3837 24266 3843
rect 24214 3779 24266 3785
rect 24226 800 24254 3779
rect 24322 3547 24350 6073
rect 24610 5860 24638 7405
rect 24514 5832 24638 5860
rect 24406 5021 24458 5027
rect 24406 4963 24458 4969
rect 24418 4583 24446 4963
rect 24406 4577 24458 4583
rect 24406 4519 24458 4525
rect 24514 4213 24542 5832
rect 24598 5687 24650 5693
rect 24598 5629 24650 5635
rect 24502 4207 24554 4213
rect 24502 4149 24554 4155
rect 24502 3911 24554 3917
rect 24502 3853 24554 3859
rect 24406 3689 24458 3695
rect 24406 3631 24458 3637
rect 24310 3541 24362 3547
rect 24310 3483 24362 3489
rect 24418 1864 24446 3631
rect 24322 1836 24446 1864
rect 24322 800 24350 1836
rect 24514 800 24542 3853
rect 24610 800 24638 5629
rect 24694 3615 24746 3621
rect 24694 3557 24746 3563
rect 24706 800 24734 3557
rect 24802 800 24830 7405
rect 25666 7099 25694 19615
rect 25942 13013 25994 13019
rect 25942 12955 25994 12961
rect 25954 7765 25982 12955
rect 26242 7765 26270 20873
rect 26722 20197 26750 43369
rect 26806 40911 26858 40917
rect 26806 40853 26858 40859
rect 26818 28115 26846 40853
rect 27190 38765 27242 38771
rect 27190 38707 27242 38713
rect 27202 38549 27230 38707
rect 27190 38543 27242 38549
rect 27190 38485 27242 38491
rect 26806 28109 26858 28115
rect 26806 28051 26858 28057
rect 27190 27887 27242 27893
rect 27190 27829 27242 27835
rect 26998 23521 27050 23527
rect 26998 23463 27050 23469
rect 26710 20191 26762 20197
rect 26710 20133 26762 20139
rect 26422 15751 26474 15757
rect 26422 15693 26474 15699
rect 25942 7759 25994 7765
rect 25942 7701 25994 7707
rect 26230 7759 26282 7765
rect 26230 7701 26282 7707
rect 25942 7463 25994 7469
rect 25942 7405 25994 7411
rect 25654 7093 25706 7099
rect 25654 7035 25706 7041
rect 25174 7019 25226 7025
rect 25174 6961 25226 6967
rect 24886 6945 24938 6951
rect 24886 6887 24938 6893
rect 24898 3917 24926 6887
rect 24886 3911 24938 3917
rect 24886 3853 24938 3859
rect 24982 3467 25034 3473
rect 24982 3409 25034 3415
rect 24886 2801 24938 2807
rect 24886 2743 24938 2749
rect 24898 2511 24926 2743
rect 24886 2505 24938 2511
rect 24886 2447 24938 2453
rect 24994 800 25022 3409
rect 25078 2949 25130 2955
rect 25078 2891 25130 2897
rect 25090 800 25118 2891
rect 25186 800 25214 6961
rect 25654 6353 25706 6359
rect 25654 6295 25706 6301
rect 25462 4355 25514 4361
rect 25462 4297 25514 4303
rect 25366 3911 25418 3917
rect 25366 3853 25418 3859
rect 25378 800 25406 3853
rect 25474 800 25502 4297
rect 25558 4207 25610 4213
rect 25558 4149 25610 4155
rect 25570 800 25598 4149
rect 25666 800 25694 6295
rect 25846 5021 25898 5027
rect 25846 4963 25898 4969
rect 25858 3843 25886 4963
rect 25954 4213 25982 7405
rect 26434 7099 26462 15693
rect 27010 7765 27038 23463
rect 26998 7759 27050 7765
rect 26998 7701 27050 7707
rect 26710 7463 26762 7469
rect 26710 7405 26762 7411
rect 26422 7093 26474 7099
rect 26422 7035 26474 7041
rect 26230 5687 26282 5693
rect 26230 5629 26282 5635
rect 26038 5613 26090 5619
rect 26038 5555 26090 5561
rect 25942 4207 25994 4213
rect 25942 4149 25994 4155
rect 25846 3837 25898 3843
rect 25846 3779 25898 3785
rect 25942 3837 25994 3843
rect 25942 3779 25994 3785
rect 25846 3541 25898 3547
rect 25846 3483 25898 3489
rect 25858 800 25886 3483
rect 25954 800 25982 3779
rect 26050 800 26078 5555
rect 26134 4355 26186 4361
rect 26134 4297 26186 4303
rect 26146 800 26174 4297
rect 26242 3917 26270 5629
rect 26614 5021 26666 5027
rect 26614 4963 26666 4969
rect 26422 4873 26474 4879
rect 26422 4815 26474 4821
rect 26230 3911 26282 3917
rect 26230 3853 26282 3859
rect 26326 3763 26378 3769
rect 26326 3705 26378 3711
rect 26338 800 26366 3705
rect 26434 800 26462 4815
rect 26518 4355 26570 4361
rect 26518 4297 26570 4303
rect 26530 800 26558 4297
rect 26626 3473 26654 4963
rect 26614 3467 26666 3473
rect 26614 3409 26666 3415
rect 26722 800 26750 7405
rect 27202 7099 27230 27829
rect 27970 7913 27998 47513
rect 28246 45425 28298 45431
rect 28246 45367 28298 45373
rect 28258 45135 28286 45367
rect 28246 45129 28298 45135
rect 28246 45071 28298 45077
rect 28150 21671 28202 21677
rect 28150 21613 28202 21619
rect 28162 9763 28190 21613
rect 28246 19599 28298 19605
rect 28246 19541 28298 19547
rect 28150 9757 28202 9763
rect 28150 9699 28202 9705
rect 28258 9412 28286 19541
rect 28162 9384 28286 9412
rect 27958 7907 28010 7913
rect 27958 7849 28010 7855
rect 28162 7636 28190 9384
rect 28246 9239 28298 9245
rect 28246 9181 28298 9187
rect 28066 7608 28190 7636
rect 28066 7173 28094 7608
rect 28150 7463 28202 7469
rect 28150 7405 28202 7411
rect 28054 7167 28106 7173
rect 28054 7109 28106 7115
rect 27190 7093 27242 7099
rect 27190 7035 27242 7041
rect 27766 7019 27818 7025
rect 27766 6961 27818 6967
rect 27094 6945 27146 6951
rect 27094 6887 27146 6893
rect 27382 6945 27434 6951
rect 27382 6887 27434 6893
rect 26806 6353 26858 6359
rect 26806 6295 26858 6301
rect 26818 800 26846 6295
rect 26998 4207 27050 4213
rect 26998 4149 27050 4155
rect 26902 3023 26954 3029
rect 26902 2965 26954 2971
rect 26914 800 26942 2965
rect 27010 800 27038 4149
rect 27106 3843 27134 6887
rect 27190 5687 27242 5693
rect 27190 5629 27242 5635
rect 27094 3837 27146 3843
rect 27094 3779 27146 3785
rect 27202 800 27230 5629
rect 27394 4213 27422 6887
rect 27574 6131 27626 6137
rect 27574 6073 27626 6079
rect 27382 4207 27434 4213
rect 27382 4149 27434 4155
rect 27478 3911 27530 3917
rect 27478 3853 27530 3859
rect 27286 3689 27338 3695
rect 27286 3631 27338 3637
rect 27298 800 27326 3631
rect 27382 3467 27434 3473
rect 27382 3409 27434 3415
rect 27394 800 27422 3409
rect 27490 800 27518 3853
rect 27586 3769 27614 6073
rect 27574 3763 27626 3769
rect 27574 3705 27626 3711
rect 27670 2949 27722 2955
rect 27670 2891 27722 2897
rect 27682 800 27710 2891
rect 27778 800 27806 6961
rect 27862 5687 27914 5693
rect 27862 5629 27914 5635
rect 27874 800 27902 5629
rect 28054 4281 28106 4287
rect 28054 4223 28106 4229
rect 28066 3843 28094 4223
rect 28054 3837 28106 3843
rect 28054 3779 28106 3785
rect 28054 3541 28106 3547
rect 28054 3483 28106 3489
rect 28066 800 28094 3483
rect 28162 800 28190 7405
rect 28258 7099 28286 9181
rect 28354 7173 28382 55135
rect 28342 7167 28394 7173
rect 28342 7109 28394 7115
rect 28246 7093 28298 7099
rect 28246 7035 28298 7041
rect 28450 5471 28478 56171
rect 29014 46387 29066 46393
rect 29014 46329 29066 46335
rect 28822 18267 28874 18273
rect 28822 18209 28874 18215
rect 28834 16793 28862 18209
rect 28822 16787 28874 16793
rect 28822 16729 28874 16735
rect 28534 9757 28586 9763
rect 28534 9699 28586 9705
rect 28546 6433 28574 9699
rect 29026 6433 29054 46329
rect 29398 35213 29450 35219
rect 29398 35155 29450 35161
rect 29302 12421 29354 12427
rect 29302 12363 29354 12369
rect 29314 11835 29342 12363
rect 29302 11829 29354 11835
rect 29302 11771 29354 11777
rect 29410 7765 29438 35155
rect 29494 16861 29546 16867
rect 29494 16803 29546 16809
rect 29398 7759 29450 7765
rect 29398 7701 29450 7707
rect 29206 7463 29258 7469
rect 29206 7405 29258 7411
rect 28534 6427 28586 6433
rect 28534 6369 28586 6375
rect 29014 6427 29066 6433
rect 29014 6369 29066 6375
rect 28822 5687 28874 5693
rect 28822 5629 28874 5635
rect 28438 5465 28490 5471
rect 28438 5407 28490 5413
rect 28342 4355 28394 4361
rect 28342 4297 28394 4303
rect 28246 4207 28298 4213
rect 28246 4149 28298 4155
rect 28258 800 28286 4149
rect 28354 800 28382 4297
rect 28534 4281 28586 4287
rect 28834 4232 28862 5629
rect 28918 5021 28970 5027
rect 28918 4963 28970 4969
rect 29014 5021 29066 5027
rect 29014 4963 29066 4969
rect 28534 4223 28586 4229
rect 28546 800 28574 4223
rect 28642 4204 28862 4232
rect 28642 800 28670 4204
rect 28930 3917 28958 4963
rect 29026 4213 29054 4963
rect 29110 4355 29162 4361
rect 29110 4297 29162 4303
rect 29014 4207 29066 4213
rect 29014 4149 29066 4155
rect 28918 3911 28970 3917
rect 28918 3853 28970 3859
rect 29014 3911 29066 3917
rect 29014 3853 29066 3859
rect 28726 3763 28778 3769
rect 28726 3705 28778 3711
rect 28738 800 28766 3705
rect 28918 2875 28970 2881
rect 28918 2817 28970 2823
rect 28930 800 28958 2817
rect 29026 800 29054 3853
rect 29122 800 29150 4297
rect 29218 800 29246 7405
rect 29506 7099 29534 16803
rect 29602 12131 29630 56171
rect 30946 51647 30974 56171
rect 31222 54231 31274 54237
rect 31222 54173 31274 54179
rect 31126 54083 31178 54089
rect 31126 54025 31178 54031
rect 30934 51641 30986 51647
rect 30934 51583 30986 51589
rect 30838 46239 30890 46245
rect 30838 46181 30890 46187
rect 30166 45203 30218 45209
rect 30166 45145 30218 45151
rect 30070 42243 30122 42249
rect 30070 42185 30122 42191
rect 30082 42101 30110 42185
rect 30070 42095 30122 42101
rect 30070 42037 30122 42043
rect 30082 37454 30110 42037
rect 29986 37426 30110 37454
rect 29986 27374 30014 37426
rect 29986 27346 30110 27374
rect 30082 25599 30110 27346
rect 30070 25593 30122 25599
rect 30070 25535 30122 25541
rect 29590 12125 29642 12131
rect 29590 12067 29642 12073
rect 30178 7765 30206 45145
rect 30742 44093 30794 44099
rect 30742 44035 30794 44041
rect 30754 43877 30782 44035
rect 30742 43871 30794 43877
rect 30742 43813 30794 43819
rect 30262 38247 30314 38253
rect 30262 38189 30314 38195
rect 30274 37454 30302 38189
rect 30274 37426 30398 37454
rect 30370 27374 30398 37426
rect 30274 27346 30398 27374
rect 30274 18791 30302 27346
rect 30646 25001 30698 25007
rect 30646 24943 30698 24949
rect 30262 18785 30314 18791
rect 30262 18727 30314 18733
rect 30166 7759 30218 7765
rect 30166 7701 30218 7707
rect 29590 7463 29642 7469
rect 29590 7405 29642 7411
rect 29494 7093 29546 7099
rect 29494 7035 29546 7041
rect 29398 6945 29450 6951
rect 29398 6887 29450 6893
rect 29302 6131 29354 6137
rect 29302 6073 29354 6079
rect 29314 3473 29342 6073
rect 29410 4287 29438 6887
rect 29398 4281 29450 4287
rect 29398 4223 29450 4229
rect 29494 3615 29546 3621
rect 29494 3557 29546 3563
rect 29302 3467 29354 3473
rect 29302 3409 29354 3415
rect 29398 3467 29450 3473
rect 29398 3409 29450 3415
rect 29410 800 29438 3409
rect 29506 800 29534 3557
rect 29602 800 29630 7405
rect 29974 6945 30026 6951
rect 29974 6887 30026 6893
rect 29686 6353 29738 6359
rect 29686 6295 29738 6301
rect 29698 800 29726 6295
rect 29782 6131 29834 6137
rect 29782 6073 29834 6079
rect 29794 2955 29822 6073
rect 29878 3023 29930 3029
rect 29878 2965 29930 2971
rect 29782 2949 29834 2955
rect 29782 2891 29834 2897
rect 29890 800 29918 2965
rect 29986 800 30014 6887
rect 30658 6433 30686 24943
rect 30850 7913 30878 46181
rect 31138 10207 31166 54025
rect 31234 10355 31262 54173
rect 32482 38327 32510 56171
rect 32470 38321 32522 38327
rect 32470 38263 32522 38269
rect 32374 38173 32426 38179
rect 32374 38115 32426 38121
rect 31702 24927 31754 24933
rect 31702 24869 31754 24875
rect 31510 16935 31562 16941
rect 31510 16877 31562 16883
rect 31522 10503 31550 16877
rect 31510 10497 31562 10503
rect 31510 10439 31562 10445
rect 31222 10349 31274 10355
rect 31222 10291 31274 10297
rect 31126 10201 31178 10207
rect 31126 10143 31178 10149
rect 30838 7907 30890 7913
rect 30838 7849 30890 7855
rect 31030 7463 31082 7469
rect 31030 7405 31082 7411
rect 30742 7167 30794 7173
rect 30742 7109 30794 7115
rect 30646 6427 30698 6433
rect 30646 6369 30698 6375
rect 30646 6131 30698 6137
rect 30646 6073 30698 6079
rect 30262 5687 30314 5693
rect 30262 5629 30314 5635
rect 30274 2894 30302 5629
rect 30358 5021 30410 5027
rect 30358 4963 30410 4969
rect 30370 3917 30398 4963
rect 30358 3911 30410 3917
rect 30358 3853 30410 3859
rect 30454 3689 30506 3695
rect 30082 2866 30302 2894
rect 30370 3649 30454 3677
rect 30082 800 30110 2866
rect 30370 1864 30398 3649
rect 30454 3631 30506 3637
rect 30454 3541 30506 3547
rect 30454 3483 30506 3489
rect 30274 1836 30398 1864
rect 30274 800 30302 1836
rect 30358 1765 30410 1771
rect 30358 1707 30410 1713
rect 30370 800 30398 1707
rect 30466 800 30494 3483
rect 30550 2949 30602 2955
rect 30550 2891 30602 2897
rect 30562 800 30590 2891
rect 30658 1771 30686 6073
rect 30646 1765 30698 1771
rect 30646 1707 30698 1713
rect 30754 800 30782 7109
rect 30838 5687 30890 5693
rect 30838 5629 30890 5635
rect 30850 800 30878 5629
rect 30934 4355 30986 4361
rect 30934 4297 30986 4303
rect 30946 800 30974 4297
rect 31042 800 31070 7405
rect 31714 7099 31742 24869
rect 32278 14789 32330 14795
rect 32278 14731 32330 14737
rect 32086 10793 32138 10799
rect 32086 10735 32138 10741
rect 31702 7093 31754 7099
rect 31702 7035 31754 7041
rect 31414 6945 31466 6951
rect 31414 6887 31466 6893
rect 31222 6353 31274 6359
rect 31222 6295 31274 6301
rect 31126 5021 31178 5027
rect 31126 4963 31178 4969
rect 31138 3473 31166 4963
rect 31126 3467 31178 3473
rect 31126 3409 31178 3415
rect 31234 800 31262 6295
rect 31318 3689 31370 3695
rect 31318 3631 31370 3637
rect 31330 800 31358 3631
rect 31426 800 31454 6887
rect 32098 6433 32126 10735
rect 32290 7025 32318 14731
rect 32386 7913 32414 38115
rect 32578 35441 32606 56837
rect 32770 56531 32798 59200
rect 33346 56975 33374 59200
rect 33334 56969 33386 56975
rect 33334 56911 33386 56917
rect 33826 56531 33854 59200
rect 34402 57614 34430 59200
rect 34402 57586 34622 57614
rect 34102 56895 34154 56901
rect 34102 56837 34154 56843
rect 32758 56525 32810 56531
rect 32758 56467 32810 56473
rect 33814 56525 33866 56531
rect 33814 56467 33866 56473
rect 32662 52085 32714 52091
rect 32662 52027 32714 52033
rect 32566 35435 32618 35441
rect 32566 35377 32618 35383
rect 32470 34103 32522 34109
rect 32470 34045 32522 34051
rect 32374 7907 32426 7913
rect 32374 7849 32426 7855
rect 32482 7099 32510 34045
rect 32674 9763 32702 52027
rect 32758 44093 32810 44099
rect 32758 44035 32810 44041
rect 33142 44093 33194 44099
rect 33142 44035 33194 44041
rect 32770 43729 32798 44035
rect 33154 43803 33182 44035
rect 33142 43797 33194 43803
rect 33142 43739 33194 43745
rect 32758 43723 32810 43729
rect 32758 43665 32810 43671
rect 32758 37137 32810 37143
rect 32758 37079 32810 37085
rect 32770 26857 32798 37079
rect 33814 34251 33866 34257
rect 33814 34193 33866 34199
rect 32758 26851 32810 26857
rect 32758 26793 32810 26799
rect 33826 23009 33854 34193
rect 33814 23003 33866 23009
rect 33814 22945 33866 22951
rect 33238 22485 33290 22491
rect 33238 22427 33290 22433
rect 33142 13901 33194 13907
rect 33142 13843 33194 13849
rect 32662 9757 32714 9763
rect 32662 9699 32714 9705
rect 32950 7241 33002 7247
rect 32950 7183 33002 7189
rect 32470 7093 32522 7099
rect 32470 7035 32522 7041
rect 32278 7019 32330 7025
rect 32278 6961 32330 6967
rect 32470 6945 32522 6951
rect 32194 6905 32470 6933
rect 32086 6427 32138 6433
rect 32086 6369 32138 6375
rect 31798 6205 31850 6211
rect 31798 6147 31850 6153
rect 31702 5687 31754 5693
rect 31702 5629 31754 5635
rect 31714 4528 31742 5629
rect 31618 4500 31742 4528
rect 31618 800 31646 4500
rect 31702 4355 31754 4361
rect 31702 4297 31754 4303
rect 31714 800 31742 4297
rect 31810 800 31838 6147
rect 31894 5021 31946 5027
rect 31894 4963 31946 4969
rect 31906 3547 31934 4963
rect 31894 3541 31946 3547
rect 31894 3483 31946 3489
rect 31894 3097 31946 3103
rect 31894 3039 31946 3045
rect 31906 800 31934 3039
rect 32086 3023 32138 3029
rect 32086 2965 32138 2971
rect 32098 800 32126 2965
rect 32194 800 32222 6905
rect 32470 6887 32522 6893
rect 32566 6353 32618 6359
rect 32566 6295 32618 6301
rect 32470 3689 32522 3695
rect 32470 3631 32522 3637
rect 32278 2949 32330 2955
rect 32278 2891 32330 2897
rect 32290 800 32318 2891
rect 32482 800 32510 3631
rect 32578 800 32606 6295
rect 32758 4355 32810 4361
rect 32758 4297 32810 4303
rect 32662 3763 32714 3769
rect 32662 3705 32714 3711
rect 32674 800 32702 3705
rect 32770 800 32798 4297
rect 32962 800 32990 7183
rect 33154 6581 33182 13843
rect 33250 7099 33278 22427
rect 34114 14277 34142 56837
rect 34594 56531 34622 57586
rect 34882 56975 34910 59200
rect 34988 57304 35284 57324
rect 35044 57302 35068 57304
rect 35124 57302 35148 57304
rect 35204 57302 35228 57304
rect 35066 57250 35068 57302
rect 35130 57250 35142 57302
rect 35204 57250 35206 57302
rect 35044 57248 35068 57250
rect 35124 57248 35148 57250
rect 35204 57248 35228 57250
rect 34988 57228 35284 57248
rect 34870 56969 34922 56975
rect 34870 56911 34922 56917
rect 35458 56531 35486 59200
rect 34582 56525 34634 56531
rect 34582 56467 34634 56473
rect 35446 56525 35498 56531
rect 35446 56467 35498 56473
rect 35938 56439 35966 59200
rect 36514 56975 36542 59200
rect 36994 57614 37022 59200
rect 36994 57586 37118 57614
rect 36502 56969 36554 56975
rect 36502 56911 36554 56917
rect 36118 56747 36170 56753
rect 36118 56689 36170 56695
rect 36886 56747 36938 56753
rect 36886 56689 36938 56695
rect 36022 56451 36074 56457
rect 35938 56411 36022 56439
rect 36022 56393 36074 56399
rect 34198 56229 34250 56235
rect 34198 56171 34250 56177
rect 34390 56229 34442 56235
rect 34390 56171 34442 56177
rect 34102 14271 34154 14277
rect 34102 14213 34154 14219
rect 34006 13753 34058 13759
rect 34006 13695 34058 13701
rect 33622 7463 33674 7469
rect 33622 7405 33674 7411
rect 33238 7093 33290 7099
rect 33238 7035 33290 7041
rect 33142 6575 33194 6581
rect 33142 6517 33194 6523
rect 33154 6285 33182 6517
rect 33142 6279 33194 6285
rect 33142 6221 33194 6227
rect 33526 6131 33578 6137
rect 33526 6073 33578 6079
rect 33142 5687 33194 5693
rect 33142 5629 33194 5635
rect 33154 2955 33182 5629
rect 33238 5613 33290 5619
rect 33238 5555 33290 5561
rect 33142 2949 33194 2955
rect 33142 2891 33194 2897
rect 33250 2752 33278 5555
rect 33334 5021 33386 5027
rect 33334 4963 33386 4969
rect 33430 5021 33482 5027
rect 33430 4963 33482 4969
rect 33346 3103 33374 4963
rect 33442 3769 33470 4963
rect 33538 3811 33566 6073
rect 33524 3802 33580 3811
rect 33430 3763 33482 3769
rect 33524 3737 33580 3746
rect 33430 3705 33482 3711
rect 33526 3689 33578 3695
rect 33526 3631 33578 3637
rect 33430 3467 33482 3473
rect 33430 3409 33482 3415
rect 33334 3097 33386 3103
rect 33334 3039 33386 3045
rect 33334 2949 33386 2955
rect 33334 2891 33386 2897
rect 33058 2724 33278 2752
rect 33058 800 33086 2724
rect 33346 1568 33374 2891
rect 33154 1540 33374 1568
rect 33154 800 33182 1540
rect 33238 1469 33290 1475
rect 33238 1411 33290 1417
rect 33250 800 33278 1411
rect 33442 800 33470 3409
rect 33538 800 33566 3631
rect 33634 800 33662 7405
rect 34018 7099 34046 13695
rect 34102 7611 34154 7617
rect 34102 7553 34154 7559
rect 34006 7093 34058 7099
rect 34006 7035 34058 7041
rect 34006 6945 34058 6951
rect 34006 6887 34058 6893
rect 33910 4355 33962 4361
rect 33910 4297 33962 4303
rect 33814 4133 33866 4139
rect 33814 4075 33866 4081
rect 33716 3358 33772 3367
rect 33716 3293 33772 3302
rect 33730 1475 33758 3293
rect 33718 1469 33770 1475
rect 33718 1411 33770 1417
rect 33826 800 33854 4075
rect 33922 800 33950 4297
rect 34018 800 34046 6887
rect 34114 2437 34142 7553
rect 34210 4583 34238 56171
rect 34402 17015 34430 56171
rect 34988 55972 35284 55992
rect 35044 55970 35068 55972
rect 35124 55970 35148 55972
rect 35204 55970 35228 55972
rect 35066 55918 35068 55970
rect 35130 55918 35142 55970
rect 35204 55918 35206 55970
rect 35044 55916 35068 55918
rect 35124 55916 35148 55918
rect 35204 55916 35228 55918
rect 34988 55896 35284 55916
rect 36130 55865 36158 56689
rect 36214 56229 36266 56235
rect 36214 56171 36266 56177
rect 36598 56229 36650 56235
rect 36598 56171 36650 56177
rect 36118 55859 36170 55865
rect 36118 55801 36170 55807
rect 35830 54749 35882 54755
rect 35830 54691 35882 54697
rect 34988 54640 35284 54660
rect 35044 54638 35068 54640
rect 35124 54638 35148 54640
rect 35204 54638 35228 54640
rect 35066 54586 35068 54638
rect 35130 54586 35142 54638
rect 35204 54586 35206 54638
rect 35044 54584 35068 54586
rect 35124 54584 35148 54586
rect 35204 54584 35228 54586
rect 34988 54564 35284 54584
rect 34870 54083 34922 54089
rect 34870 54025 34922 54031
rect 34774 44093 34826 44099
rect 34774 44035 34826 44041
rect 34678 42761 34730 42767
rect 34678 42703 34730 42709
rect 34690 42545 34718 42703
rect 34678 42539 34730 42545
rect 34678 42481 34730 42487
rect 34786 17294 34814 44035
rect 34690 17266 34814 17294
rect 34390 17009 34442 17015
rect 34390 16951 34442 16957
rect 34582 14197 34634 14203
rect 34582 14139 34634 14145
rect 34594 7765 34622 14139
rect 34582 7759 34634 7765
rect 34582 7701 34634 7707
rect 34390 7463 34442 7469
rect 34390 7405 34442 7411
rect 34294 6279 34346 6285
rect 34294 6221 34346 6227
rect 34306 5767 34334 6221
rect 34294 5761 34346 5767
rect 34294 5703 34346 5709
rect 34198 4577 34250 4583
rect 34198 4519 34250 4525
rect 34198 4281 34250 4287
rect 34198 4223 34250 4229
rect 34102 2431 34154 2437
rect 34102 2373 34154 2379
rect 34210 2160 34238 4223
rect 34294 3689 34346 3695
rect 34294 3631 34346 3637
rect 34114 2132 34238 2160
rect 34114 800 34142 2132
rect 34306 800 34334 3631
rect 34402 800 34430 7405
rect 34690 6803 34718 17266
rect 34882 15683 34910 54025
rect 34988 53308 35284 53328
rect 35044 53306 35068 53308
rect 35124 53306 35148 53308
rect 35204 53306 35228 53308
rect 35066 53254 35068 53306
rect 35130 53254 35142 53306
rect 35204 53254 35206 53306
rect 35044 53252 35068 53254
rect 35124 53252 35148 53254
rect 35204 53252 35228 53254
rect 34988 53232 35284 53252
rect 34988 51976 35284 51996
rect 35044 51974 35068 51976
rect 35124 51974 35148 51976
rect 35204 51974 35228 51976
rect 35066 51922 35068 51974
rect 35130 51922 35142 51974
rect 35204 51922 35206 51974
rect 35044 51920 35068 51922
rect 35124 51920 35148 51922
rect 35204 51920 35228 51922
rect 34988 51900 35284 51920
rect 34988 50644 35284 50664
rect 35044 50642 35068 50644
rect 35124 50642 35148 50644
rect 35204 50642 35228 50644
rect 35066 50590 35068 50642
rect 35130 50590 35142 50642
rect 35204 50590 35206 50642
rect 35044 50588 35068 50590
rect 35124 50588 35148 50590
rect 35204 50588 35228 50590
rect 34988 50568 35284 50588
rect 34988 49312 35284 49332
rect 35044 49310 35068 49312
rect 35124 49310 35148 49312
rect 35204 49310 35228 49312
rect 35066 49258 35068 49310
rect 35130 49258 35142 49310
rect 35204 49258 35206 49310
rect 35044 49256 35068 49258
rect 35124 49256 35148 49258
rect 35204 49256 35228 49258
rect 34988 49236 35284 49256
rect 34988 47980 35284 48000
rect 35044 47978 35068 47980
rect 35124 47978 35148 47980
rect 35204 47978 35228 47980
rect 35066 47926 35068 47978
rect 35130 47926 35142 47978
rect 35204 47926 35206 47978
rect 35044 47924 35068 47926
rect 35124 47924 35148 47926
rect 35204 47924 35228 47926
rect 34988 47904 35284 47924
rect 34988 46648 35284 46668
rect 35044 46646 35068 46648
rect 35124 46646 35148 46648
rect 35204 46646 35228 46648
rect 35066 46594 35068 46646
rect 35130 46594 35142 46646
rect 35204 46594 35206 46646
rect 35044 46592 35068 46594
rect 35124 46592 35148 46594
rect 35204 46592 35228 46594
rect 34988 46572 35284 46592
rect 35842 46393 35870 54691
rect 35830 46387 35882 46393
rect 35830 46329 35882 46335
rect 34988 45316 35284 45336
rect 35044 45314 35068 45316
rect 35124 45314 35148 45316
rect 35204 45314 35228 45316
rect 35066 45262 35068 45314
rect 35130 45262 35142 45314
rect 35204 45262 35206 45314
rect 35044 45260 35068 45262
rect 35124 45260 35148 45262
rect 35204 45260 35228 45262
rect 34988 45240 35284 45260
rect 34988 43984 35284 44004
rect 35044 43982 35068 43984
rect 35124 43982 35148 43984
rect 35204 43982 35228 43984
rect 35066 43930 35068 43982
rect 35130 43930 35142 43982
rect 35204 43930 35206 43982
rect 35044 43928 35068 43930
rect 35124 43928 35148 43930
rect 35204 43928 35228 43930
rect 34988 43908 35284 43928
rect 34988 42652 35284 42672
rect 35044 42650 35068 42652
rect 35124 42650 35148 42652
rect 35204 42650 35228 42652
rect 35066 42598 35068 42650
rect 35130 42598 35142 42650
rect 35204 42598 35206 42650
rect 35044 42596 35068 42598
rect 35124 42596 35148 42598
rect 35204 42596 35228 42598
rect 34988 42576 35284 42596
rect 34988 41320 35284 41340
rect 35044 41318 35068 41320
rect 35124 41318 35148 41320
rect 35204 41318 35228 41320
rect 35066 41266 35068 41318
rect 35130 41266 35142 41318
rect 35204 41266 35206 41318
rect 35044 41264 35068 41266
rect 35124 41264 35148 41266
rect 35204 41264 35228 41266
rect 34988 41244 35284 41264
rect 34988 39988 35284 40008
rect 35044 39986 35068 39988
rect 35124 39986 35148 39988
rect 35204 39986 35228 39988
rect 35066 39934 35068 39986
rect 35130 39934 35142 39986
rect 35204 39934 35206 39986
rect 35044 39932 35068 39934
rect 35124 39932 35148 39934
rect 35204 39932 35228 39934
rect 34988 39912 35284 39932
rect 36226 38845 36254 56171
rect 36310 54083 36362 54089
rect 36310 54025 36362 54031
rect 36214 38839 36266 38845
rect 36214 38781 36266 38787
rect 34988 38656 35284 38676
rect 35044 38654 35068 38656
rect 35124 38654 35148 38656
rect 35204 38654 35228 38656
rect 35066 38602 35068 38654
rect 35130 38602 35142 38654
rect 35204 38602 35206 38654
rect 35044 38600 35068 38602
rect 35124 38600 35148 38602
rect 35204 38600 35228 38602
rect 34988 38580 35284 38600
rect 34988 37324 35284 37344
rect 35044 37322 35068 37324
rect 35124 37322 35148 37324
rect 35204 37322 35228 37324
rect 35066 37270 35068 37322
rect 35130 37270 35142 37322
rect 35204 37270 35206 37322
rect 35044 37268 35068 37270
rect 35124 37268 35148 37270
rect 35204 37268 35228 37270
rect 34988 37248 35284 37268
rect 34988 35992 35284 36012
rect 35044 35990 35068 35992
rect 35124 35990 35148 35992
rect 35204 35990 35228 35992
rect 35066 35938 35068 35990
rect 35130 35938 35142 35990
rect 35204 35938 35206 35990
rect 35044 35936 35068 35938
rect 35124 35936 35148 35938
rect 35204 35936 35228 35938
rect 34988 35916 35284 35936
rect 35926 35509 35978 35515
rect 35926 35451 35978 35457
rect 34988 34660 35284 34680
rect 35044 34658 35068 34660
rect 35124 34658 35148 34660
rect 35204 34658 35228 34660
rect 35066 34606 35068 34658
rect 35130 34606 35142 34658
rect 35204 34606 35206 34658
rect 35044 34604 35068 34606
rect 35124 34604 35148 34606
rect 35204 34604 35228 34606
rect 34988 34584 35284 34604
rect 34988 33328 35284 33348
rect 35044 33326 35068 33328
rect 35124 33326 35148 33328
rect 35204 33326 35228 33328
rect 35066 33274 35068 33326
rect 35130 33274 35142 33326
rect 35204 33274 35206 33326
rect 35044 33272 35068 33274
rect 35124 33272 35148 33274
rect 35204 33272 35228 33274
rect 34988 33252 35284 33272
rect 34988 31996 35284 32016
rect 35044 31994 35068 31996
rect 35124 31994 35148 31996
rect 35204 31994 35228 31996
rect 35066 31942 35068 31994
rect 35130 31942 35142 31994
rect 35204 31942 35206 31994
rect 35044 31940 35068 31942
rect 35124 31940 35148 31942
rect 35204 31940 35228 31942
rect 34988 31920 35284 31940
rect 34988 30664 35284 30684
rect 35044 30662 35068 30664
rect 35124 30662 35148 30664
rect 35204 30662 35228 30664
rect 35066 30610 35068 30662
rect 35130 30610 35142 30662
rect 35204 30610 35206 30662
rect 35044 30608 35068 30610
rect 35124 30608 35148 30610
rect 35204 30608 35228 30610
rect 34988 30588 35284 30608
rect 34988 29332 35284 29352
rect 35044 29330 35068 29332
rect 35124 29330 35148 29332
rect 35204 29330 35228 29332
rect 35066 29278 35068 29330
rect 35130 29278 35142 29330
rect 35204 29278 35206 29330
rect 35044 29276 35068 29278
rect 35124 29276 35148 29278
rect 35204 29276 35228 29278
rect 34988 29256 35284 29276
rect 34988 28000 35284 28020
rect 35044 27998 35068 28000
rect 35124 27998 35148 28000
rect 35204 27998 35228 28000
rect 35066 27946 35068 27998
rect 35130 27946 35142 27998
rect 35204 27946 35206 27998
rect 35044 27944 35068 27946
rect 35124 27944 35148 27946
rect 35204 27944 35228 27946
rect 34988 27924 35284 27944
rect 34988 26668 35284 26688
rect 35044 26666 35068 26668
rect 35124 26666 35148 26668
rect 35204 26666 35228 26668
rect 35066 26614 35068 26666
rect 35130 26614 35142 26666
rect 35204 26614 35206 26666
rect 35044 26612 35068 26614
rect 35124 26612 35148 26614
rect 35204 26612 35228 26614
rect 34988 26592 35284 26612
rect 34988 25336 35284 25356
rect 35044 25334 35068 25336
rect 35124 25334 35148 25336
rect 35204 25334 35228 25336
rect 35066 25282 35068 25334
rect 35130 25282 35142 25334
rect 35204 25282 35206 25334
rect 35044 25280 35068 25282
rect 35124 25280 35148 25282
rect 35204 25280 35228 25282
rect 34988 25260 35284 25280
rect 34988 24004 35284 24024
rect 35044 24002 35068 24004
rect 35124 24002 35148 24004
rect 35204 24002 35228 24004
rect 35066 23950 35068 24002
rect 35130 23950 35142 24002
rect 35204 23950 35206 24002
rect 35044 23948 35068 23950
rect 35124 23948 35148 23950
rect 35204 23948 35228 23950
rect 34988 23928 35284 23948
rect 34988 22672 35284 22692
rect 35044 22670 35068 22672
rect 35124 22670 35148 22672
rect 35204 22670 35228 22672
rect 35066 22618 35068 22670
rect 35130 22618 35142 22670
rect 35204 22618 35206 22670
rect 35044 22616 35068 22618
rect 35124 22616 35148 22618
rect 35204 22616 35228 22618
rect 34988 22596 35284 22616
rect 34988 21340 35284 21360
rect 35044 21338 35068 21340
rect 35124 21338 35148 21340
rect 35204 21338 35228 21340
rect 35066 21286 35068 21338
rect 35130 21286 35142 21338
rect 35204 21286 35206 21338
rect 35044 21284 35068 21286
rect 35124 21284 35148 21286
rect 35204 21284 35228 21286
rect 34988 21264 35284 21284
rect 34988 20008 35284 20028
rect 35044 20006 35068 20008
rect 35124 20006 35148 20008
rect 35204 20006 35228 20008
rect 35066 19954 35068 20006
rect 35130 19954 35142 20006
rect 35204 19954 35206 20006
rect 35044 19952 35068 19954
rect 35124 19952 35148 19954
rect 35204 19952 35228 19954
rect 34988 19932 35284 19952
rect 34988 18676 35284 18696
rect 35044 18674 35068 18676
rect 35124 18674 35148 18676
rect 35204 18674 35228 18676
rect 35066 18622 35068 18674
rect 35130 18622 35142 18674
rect 35204 18622 35206 18674
rect 35044 18620 35068 18622
rect 35124 18620 35148 18622
rect 35204 18620 35228 18622
rect 34988 18600 35284 18620
rect 34988 17344 35284 17364
rect 35044 17342 35068 17344
rect 35124 17342 35148 17344
rect 35204 17342 35228 17344
rect 35066 17290 35068 17342
rect 35130 17290 35142 17342
rect 35204 17290 35206 17342
rect 35044 17288 35068 17290
rect 35124 17288 35148 17290
rect 35204 17288 35228 17290
rect 34988 17268 35284 17288
rect 34988 16012 35284 16032
rect 35044 16010 35068 16012
rect 35124 16010 35148 16012
rect 35204 16010 35228 16012
rect 35066 15958 35068 16010
rect 35130 15958 35142 16010
rect 35204 15958 35206 16010
rect 35044 15956 35068 15958
rect 35124 15956 35148 15958
rect 35204 15956 35228 15958
rect 34988 15936 35284 15956
rect 34870 15677 34922 15683
rect 34870 15619 34922 15625
rect 34988 14680 35284 14700
rect 35044 14678 35068 14680
rect 35124 14678 35148 14680
rect 35204 14678 35228 14680
rect 35066 14626 35068 14678
rect 35130 14626 35142 14678
rect 35204 14626 35206 14678
rect 35044 14624 35068 14626
rect 35124 14624 35148 14626
rect 35204 14624 35228 14626
rect 34988 14604 35284 14624
rect 34988 13348 35284 13368
rect 35044 13346 35068 13348
rect 35124 13346 35148 13348
rect 35204 13346 35228 13348
rect 35066 13294 35068 13346
rect 35130 13294 35142 13346
rect 35204 13294 35206 13346
rect 35044 13292 35068 13294
rect 35124 13292 35148 13294
rect 35204 13292 35228 13294
rect 34988 13272 35284 13292
rect 34988 12016 35284 12036
rect 35044 12014 35068 12016
rect 35124 12014 35148 12016
rect 35204 12014 35228 12016
rect 35066 11962 35068 12014
rect 35130 11962 35142 12014
rect 35204 11962 35206 12014
rect 35044 11960 35068 11962
rect 35124 11960 35148 11962
rect 35204 11960 35228 11962
rect 34988 11940 35284 11960
rect 34988 10684 35284 10704
rect 35044 10682 35068 10684
rect 35124 10682 35148 10684
rect 35204 10682 35228 10684
rect 35066 10630 35068 10682
rect 35130 10630 35142 10682
rect 35204 10630 35206 10682
rect 35044 10628 35068 10630
rect 35124 10628 35148 10630
rect 35204 10628 35228 10630
rect 34988 10608 35284 10628
rect 35350 10423 35402 10429
rect 35350 10365 35402 10371
rect 34988 9352 35284 9372
rect 35044 9350 35068 9352
rect 35124 9350 35148 9352
rect 35204 9350 35228 9352
rect 35066 9298 35068 9350
rect 35130 9298 35142 9350
rect 35204 9298 35206 9350
rect 35044 9296 35068 9298
rect 35124 9296 35148 9298
rect 35204 9296 35228 9298
rect 34988 9276 35284 9296
rect 34988 8020 35284 8040
rect 35044 8018 35068 8020
rect 35124 8018 35148 8020
rect 35204 8018 35228 8020
rect 35066 7966 35068 8018
rect 35130 7966 35142 8018
rect 35204 7966 35206 8018
rect 35044 7964 35068 7966
rect 35124 7964 35148 7966
rect 35204 7964 35228 7966
rect 34988 7944 35284 7964
rect 35362 7765 35390 10365
rect 35938 7913 35966 35451
rect 36322 25229 36350 54025
rect 36310 25223 36362 25229
rect 36310 25165 36362 25171
rect 36310 22781 36362 22787
rect 36310 22723 36362 22729
rect 36322 12974 36350 22723
rect 36610 13537 36638 56171
rect 36694 34251 36746 34257
rect 36694 34193 36746 34199
rect 36598 13531 36650 13537
rect 36598 13473 36650 13479
rect 36226 12946 36350 12974
rect 35926 7907 35978 7913
rect 35926 7849 35978 7855
rect 35350 7759 35402 7765
rect 35350 7701 35402 7707
rect 34774 7463 34826 7469
rect 34774 7405 34826 7411
rect 36022 7463 36074 7469
rect 36022 7405 36074 7411
rect 34678 6797 34730 6803
rect 34678 6739 34730 6745
rect 34678 5687 34730 5693
rect 34678 5629 34730 5635
rect 34582 4355 34634 4361
rect 34582 4297 34634 4303
rect 34486 3911 34538 3917
rect 34486 3853 34538 3859
rect 34498 800 34526 3853
rect 34594 800 34622 4297
rect 34690 4139 34718 5629
rect 34678 4133 34730 4139
rect 34678 4075 34730 4081
rect 34786 800 34814 7405
rect 35446 7167 35498 7173
rect 35446 7109 35498 7115
rect 35350 6945 35402 6951
rect 35350 6887 35402 6893
rect 34988 6688 35284 6708
rect 35044 6686 35068 6688
rect 35124 6686 35148 6688
rect 35204 6686 35228 6688
rect 35066 6634 35068 6686
rect 35130 6634 35142 6686
rect 35204 6634 35206 6686
rect 35044 6632 35068 6634
rect 35124 6632 35148 6634
rect 35204 6632 35228 6634
rect 34988 6612 35284 6632
rect 34988 5356 35284 5376
rect 35044 5354 35068 5356
rect 35124 5354 35148 5356
rect 35204 5354 35228 5356
rect 35066 5302 35068 5354
rect 35130 5302 35142 5354
rect 35204 5302 35206 5354
rect 35044 5300 35068 5302
rect 35124 5300 35148 5302
rect 35204 5300 35228 5302
rect 34988 5280 35284 5300
rect 34870 5021 34922 5027
rect 34870 4963 34922 4969
rect 34882 3473 34910 4963
rect 34988 4024 35284 4044
rect 35044 4022 35068 4024
rect 35124 4022 35148 4024
rect 35204 4022 35228 4024
rect 35066 3970 35068 4022
rect 35130 3970 35142 4022
rect 35204 3970 35206 4022
rect 35044 3968 35068 3970
rect 35124 3968 35148 3970
rect 35204 3968 35228 3970
rect 34988 3948 35284 3968
rect 35362 3788 35390 6887
rect 35458 3843 35486 7109
rect 35542 6945 35594 6951
rect 35542 6887 35594 6893
rect 35266 3760 35390 3788
rect 35446 3837 35498 3843
rect 35446 3779 35498 3785
rect 34966 3689 35018 3695
rect 34966 3631 35018 3637
rect 34870 3467 34922 3473
rect 34870 3409 34922 3415
rect 34978 2894 35006 3631
rect 34882 2866 35006 2894
rect 34882 1864 34910 2866
rect 35266 2807 35294 3760
rect 35350 3615 35402 3621
rect 35350 3557 35402 3563
rect 35254 2801 35306 2807
rect 35254 2743 35306 2749
rect 34988 2692 35284 2712
rect 35044 2690 35068 2692
rect 35124 2690 35148 2692
rect 35204 2690 35228 2692
rect 35066 2638 35068 2690
rect 35130 2638 35142 2690
rect 35204 2638 35206 2690
rect 35044 2636 35068 2638
rect 35124 2636 35148 2638
rect 35204 2636 35228 2638
rect 34988 2616 35284 2636
rect 35158 2579 35210 2585
rect 35158 2521 35210 2527
rect 34882 1836 35006 1864
rect 34870 1765 34922 1771
rect 34870 1707 34922 1713
rect 34882 800 34910 1707
rect 34978 800 35006 1836
rect 35170 800 35198 2521
rect 35362 2456 35390 3557
rect 35446 3023 35498 3029
rect 35446 2965 35498 2971
rect 35266 2428 35390 2456
rect 35266 800 35294 2428
rect 35458 1568 35486 2965
rect 35554 2585 35582 6887
rect 35734 6279 35786 6285
rect 35734 6221 35786 6227
rect 35638 5021 35690 5027
rect 35638 4963 35690 4969
rect 35650 3917 35678 4963
rect 35638 3911 35690 3917
rect 35638 3853 35690 3859
rect 35746 3751 35774 6221
rect 36034 4232 36062 7405
rect 36226 5915 36254 12946
rect 36706 10947 36734 34193
rect 36898 30409 36926 56689
rect 37090 56161 37118 57586
rect 37570 56531 37598 59200
rect 38050 56975 38078 59200
rect 38038 56969 38090 56975
rect 38038 56911 38090 56917
rect 38626 56531 38654 59200
rect 37558 56525 37610 56531
rect 37558 56467 37610 56473
rect 38614 56525 38666 56531
rect 38614 56467 38666 56473
rect 38902 56451 38954 56457
rect 38902 56393 38954 56399
rect 37750 56229 37802 56235
rect 37750 56171 37802 56177
rect 38710 56229 38762 56235
rect 38710 56171 38762 56177
rect 38806 56229 38858 56235
rect 38806 56171 38858 56177
rect 37078 56155 37130 56161
rect 37078 56097 37130 56103
rect 36886 30403 36938 30409
rect 36886 30345 36938 30351
rect 37762 28559 37790 56171
rect 38134 42835 38186 42841
rect 38134 42777 38186 42783
rect 37750 28553 37802 28559
rect 37750 28495 37802 28501
rect 36982 25445 37034 25451
rect 36982 25387 37034 25393
rect 36886 23743 36938 23749
rect 36886 23685 36938 23691
rect 36790 19525 36842 19531
rect 36790 19467 36842 19473
rect 36694 10941 36746 10947
rect 36694 10883 36746 10889
rect 36694 8869 36746 8875
rect 36694 8811 36746 8817
rect 36598 7463 36650 7469
rect 36598 7405 36650 7411
rect 36502 6945 36554 6951
rect 36502 6887 36554 6893
rect 36310 6353 36362 6359
rect 36310 6295 36362 6301
rect 36214 5909 36266 5915
rect 36214 5851 36266 5857
rect 36214 5687 36266 5693
rect 36214 5629 36266 5635
rect 36118 5021 36170 5027
rect 36118 4963 36170 4969
rect 35650 3723 35774 3751
rect 35842 4204 36062 4232
rect 35650 3071 35678 3723
rect 35734 3689 35786 3695
rect 35734 3631 35786 3637
rect 35636 3062 35692 3071
rect 35636 2997 35692 3006
rect 35638 2875 35690 2881
rect 35638 2817 35690 2823
rect 35542 2579 35594 2585
rect 35542 2521 35594 2527
rect 35540 2470 35596 2479
rect 35540 2405 35596 2414
rect 35362 1540 35486 1568
rect 35362 800 35390 1540
rect 35554 1420 35582 2405
rect 35458 1392 35582 1420
rect 35458 800 35486 1392
rect 35650 800 35678 2817
rect 35746 800 35774 3631
rect 35842 800 35870 4204
rect 36130 3936 36158 4963
rect 35938 3908 36158 3936
rect 35938 1771 35966 3908
rect 36022 3837 36074 3843
rect 36022 3779 36074 3785
rect 35926 1765 35978 1771
rect 35926 1707 35978 1713
rect 36034 800 36062 3779
rect 36226 3621 36254 5629
rect 36214 3615 36266 3621
rect 36214 3557 36266 3563
rect 36214 2949 36266 2955
rect 36214 2891 36266 2897
rect 36226 1568 36254 2891
rect 36130 1540 36254 1568
rect 36322 1549 36350 6295
rect 36406 5687 36458 5693
rect 36406 5629 36458 5635
rect 36418 3843 36446 5629
rect 36406 3837 36458 3843
rect 36406 3779 36458 3785
rect 36514 3751 36542 6887
rect 36418 3723 36542 3751
rect 36310 1543 36362 1549
rect 36130 800 36158 1540
rect 36310 1485 36362 1491
rect 36418 1420 36446 3723
rect 36502 3689 36554 3695
rect 36502 3631 36554 3637
rect 36226 1392 36446 1420
rect 36226 800 36254 1392
rect 36310 1173 36362 1179
rect 36310 1115 36362 1121
rect 36322 800 36350 1115
rect 36514 800 36542 3631
rect 36610 800 36638 7405
rect 36706 6581 36734 8811
rect 36802 7765 36830 19467
rect 36790 7759 36842 7765
rect 36790 7701 36842 7707
rect 36898 7099 36926 23685
rect 36994 10429 37022 25387
rect 38146 21603 38174 42777
rect 38518 36101 38570 36107
rect 38518 36043 38570 36049
rect 38230 30551 38282 30557
rect 38230 30493 38282 30499
rect 38134 21597 38186 21603
rect 38134 21539 38186 21545
rect 37654 18785 37706 18791
rect 37654 18727 37706 18733
rect 37462 17527 37514 17533
rect 37462 17469 37514 17475
rect 37474 11095 37502 17469
rect 37462 11089 37514 11095
rect 37462 11031 37514 11037
rect 36982 10423 37034 10429
rect 36982 10365 37034 10371
rect 37666 7099 37694 18727
rect 38242 10873 38270 30493
rect 38326 30329 38378 30335
rect 38326 30271 38378 30277
rect 38338 11021 38366 30271
rect 38422 21449 38474 21455
rect 38422 21391 38474 21397
rect 38434 13833 38462 21391
rect 38422 13827 38474 13833
rect 38422 13769 38474 13775
rect 38530 11021 38558 36043
rect 38722 24785 38750 56171
rect 38818 50167 38846 56171
rect 38914 55791 38942 56393
rect 38902 55785 38954 55791
rect 38902 55727 38954 55733
rect 39106 55199 39134 59200
rect 39682 56901 39710 59200
rect 39670 56895 39722 56901
rect 39670 56837 39722 56843
rect 39862 56821 39914 56827
rect 39778 56769 39862 56772
rect 39778 56763 39914 56769
rect 39670 56747 39722 56753
rect 39670 56689 39722 56695
rect 39778 56744 39902 56763
rect 39094 55193 39146 55199
rect 39094 55135 39146 55141
rect 39286 54897 39338 54903
rect 39286 54839 39338 54845
rect 38806 50161 38858 50167
rect 38806 50103 38858 50109
rect 38902 45425 38954 45431
rect 38902 45367 38954 45373
rect 38914 45209 38942 45367
rect 38902 45203 38954 45209
rect 38902 45145 38954 45151
rect 39190 38543 39242 38549
rect 39190 38485 39242 38491
rect 38710 24779 38762 24785
rect 38710 24721 38762 24727
rect 38806 23003 38858 23009
rect 38806 22945 38858 22951
rect 38326 11015 38378 11021
rect 38326 10957 38378 10963
rect 38518 11015 38570 11021
rect 38518 10957 38570 10963
rect 38230 10867 38282 10873
rect 38230 10809 38282 10815
rect 38818 7765 38846 22945
rect 38902 16787 38954 16793
rect 38902 16729 38954 16735
rect 38806 7759 38858 7765
rect 38806 7701 38858 7707
rect 38038 7463 38090 7469
rect 38038 7405 38090 7411
rect 38806 7463 38858 7469
rect 38806 7405 38858 7411
rect 36886 7093 36938 7099
rect 36886 7035 36938 7041
rect 37654 7093 37706 7099
rect 37654 7035 37706 7041
rect 37078 6945 37130 6951
rect 37078 6887 37130 6893
rect 36694 6575 36746 6581
rect 36694 6517 36746 6523
rect 36706 6285 36734 6517
rect 36694 6279 36746 6285
rect 36694 6221 36746 6227
rect 36886 5021 36938 5027
rect 37090 4972 37118 6887
rect 37270 6871 37322 6877
rect 37270 6813 37322 6819
rect 37366 6871 37418 6877
rect 37366 6813 37418 6819
rect 37282 6507 37310 6813
rect 37270 6501 37322 6507
rect 37270 6443 37322 6449
rect 36886 4963 36938 4969
rect 36790 4355 36842 4361
rect 36790 4297 36842 4303
rect 36694 4133 36746 4139
rect 36694 4075 36746 4081
rect 36706 800 36734 4075
rect 36802 800 36830 4297
rect 36898 2881 36926 4963
rect 36994 4944 37118 4972
rect 36886 2875 36938 2881
rect 36886 2817 36938 2823
rect 36994 800 37022 4944
rect 37174 4281 37226 4287
rect 37174 4223 37226 4229
rect 37078 3837 37130 3843
rect 37078 3779 37130 3785
rect 37090 800 37118 3779
rect 37186 800 37214 4223
rect 37270 2875 37322 2881
rect 37270 2817 37322 2823
rect 37282 2437 37310 2817
rect 37270 2431 37322 2437
rect 37270 2373 37322 2379
rect 37378 800 37406 6813
rect 37654 6797 37706 6803
rect 37654 6739 37706 6745
rect 37558 5687 37610 5693
rect 37558 5629 37610 5635
rect 37462 5613 37514 5619
rect 37462 5555 37514 5561
rect 37474 800 37502 5555
rect 37570 4139 37598 5629
rect 37558 4133 37610 4139
rect 37558 4075 37610 4081
rect 37558 3023 37610 3029
rect 37558 2965 37610 2971
rect 37570 800 37598 2965
rect 37666 800 37694 6739
rect 37846 5465 37898 5471
rect 37846 5407 37898 5413
rect 37858 4805 37886 5407
rect 37846 4799 37898 4805
rect 37846 4741 37898 4747
rect 37942 3689 37994 3695
rect 37942 3631 37994 3637
rect 37846 3541 37898 3547
rect 37846 3483 37898 3489
rect 37858 800 37886 3483
rect 37954 800 37982 3631
rect 38050 800 38078 7405
rect 38422 6575 38474 6581
rect 38422 6517 38474 6523
rect 38134 3911 38186 3917
rect 38134 3853 38186 3859
rect 38146 800 38174 3853
rect 38326 2949 38378 2955
rect 38326 2891 38378 2897
rect 38338 800 38366 2891
rect 38434 800 38462 6517
rect 38614 5021 38666 5027
rect 38614 4963 38666 4969
rect 38518 4133 38570 4139
rect 38518 4075 38570 4081
rect 38530 800 38558 4075
rect 38626 3843 38654 4963
rect 38614 3837 38666 3843
rect 38614 3779 38666 3785
rect 38710 3689 38762 3695
rect 38710 3631 38762 3637
rect 38722 800 38750 3631
rect 38818 800 38846 7405
rect 38914 7173 38942 16729
rect 39202 8579 39230 38485
rect 39298 30483 39326 54839
rect 39286 30477 39338 30483
rect 39286 30419 39338 30425
rect 39478 21597 39530 21603
rect 39478 21539 39530 21545
rect 39190 8573 39242 8579
rect 39190 8515 39242 8521
rect 39190 8277 39242 8283
rect 39190 8219 39242 8225
rect 38902 7167 38954 7173
rect 38902 7109 38954 7115
rect 38902 6353 38954 6359
rect 38902 6295 38954 6301
rect 38914 800 38942 6295
rect 39094 5687 39146 5693
rect 39094 5629 39146 5635
rect 38998 4355 39050 4361
rect 38998 4297 39050 4303
rect 39010 800 39038 4297
rect 39106 3917 39134 5629
rect 39094 3911 39146 3917
rect 39094 3853 39146 3859
rect 39202 800 39230 8219
rect 39490 7765 39518 21539
rect 39682 9689 39710 56689
rect 39778 55421 39806 56744
rect 40162 56531 40190 59200
rect 40342 56747 40394 56753
rect 40342 56689 40394 56695
rect 40150 56525 40202 56531
rect 40150 56467 40202 56473
rect 40354 56161 40382 56689
rect 40738 56161 40766 59200
rect 41218 56975 41246 59200
rect 41206 56969 41258 56975
rect 41206 56911 41258 56917
rect 40822 56895 40874 56901
rect 40822 56837 40874 56843
rect 40342 56155 40394 56161
rect 40342 56097 40394 56103
rect 40726 56155 40778 56161
rect 40726 56097 40778 56103
rect 39766 55415 39818 55421
rect 39766 55357 39818 55363
rect 39862 54749 39914 54755
rect 39862 54691 39914 54697
rect 39874 16571 39902 54691
rect 40834 42101 40862 56837
rect 41794 56531 41822 59200
rect 41782 56525 41834 56531
rect 41782 56467 41834 56473
rect 41782 56303 41834 56309
rect 41782 56245 41834 56251
rect 41590 56229 41642 56235
rect 41590 56171 41642 56177
rect 41014 46165 41066 46171
rect 41014 46107 41066 46113
rect 40822 42095 40874 42101
rect 40822 42037 40874 42043
rect 39958 35583 40010 35589
rect 39958 35525 40010 35531
rect 39862 16565 39914 16571
rect 39862 16507 39914 16513
rect 39670 9683 39722 9689
rect 39670 9625 39722 9631
rect 39970 7913 39998 35525
rect 40918 30847 40970 30853
rect 40918 30789 40970 30795
rect 40930 30483 40958 30789
rect 40918 30477 40970 30483
rect 40918 30419 40970 30425
rect 40150 26259 40202 26265
rect 40150 26201 40202 26207
rect 40162 25229 40190 26201
rect 40150 25223 40202 25229
rect 40150 25165 40202 25171
rect 40054 22411 40106 22417
rect 40054 22353 40106 22359
rect 39958 7907 40010 7913
rect 39958 7849 40010 7855
rect 39478 7759 39530 7765
rect 39478 7701 39530 7707
rect 39958 7537 40010 7543
rect 39958 7479 40010 7485
rect 39670 7463 39722 7469
rect 39670 7405 39722 7411
rect 39286 6945 39338 6951
rect 39286 6887 39338 6893
rect 39298 6581 39326 6887
rect 39286 6575 39338 6581
rect 39286 6517 39338 6523
rect 39286 5687 39338 5693
rect 39286 5629 39338 5635
rect 39298 800 39326 5629
rect 39382 5021 39434 5027
rect 39382 4963 39434 4969
rect 39394 3547 39422 4963
rect 39682 4084 39710 7405
rect 39862 6871 39914 6877
rect 39862 6813 39914 6819
rect 39766 4355 39818 4361
rect 39766 4297 39818 4303
rect 39586 4056 39710 4084
rect 39478 3689 39530 3695
rect 39478 3631 39530 3637
rect 39382 3541 39434 3547
rect 39382 3483 39434 3489
rect 39490 3233 39518 3631
rect 39394 3205 39518 3233
rect 39394 800 39422 3205
rect 39586 2894 39614 4056
rect 39670 3911 39722 3917
rect 39670 3853 39722 3859
rect 39490 2866 39614 2894
rect 39490 800 39518 2866
rect 39682 800 39710 3853
rect 39778 800 39806 4297
rect 39874 800 39902 6813
rect 39970 1771 39998 7479
rect 40066 7099 40094 22353
rect 41026 13019 41054 46107
rect 41110 42539 41162 42545
rect 41110 42481 41162 42487
rect 41122 14203 41150 42481
rect 41206 40763 41258 40769
rect 41206 40705 41258 40711
rect 41218 14573 41246 40705
rect 41302 38765 41354 38771
rect 41302 38707 41354 38713
rect 41314 15535 41342 38707
rect 41398 33511 41450 33517
rect 41398 33453 41450 33459
rect 41302 15529 41354 15535
rect 41302 15471 41354 15477
rect 41206 14567 41258 14573
rect 41206 14509 41258 14515
rect 41110 14197 41162 14203
rect 41110 14139 41162 14145
rect 41410 13907 41438 33453
rect 41602 29447 41630 56171
rect 41794 55865 41822 56245
rect 41782 55859 41834 55865
rect 41782 55801 41834 55807
rect 42274 55717 42302 59200
rect 42850 56975 42878 59200
rect 42838 56969 42890 56975
rect 42838 56911 42890 56917
rect 43030 56895 43082 56901
rect 43030 56837 43082 56843
rect 42838 56821 42890 56827
rect 42838 56763 42890 56769
rect 42262 55711 42314 55717
rect 42262 55653 42314 55659
rect 42550 55563 42602 55569
rect 42550 55505 42602 55511
rect 42070 41429 42122 41435
rect 42070 41371 42122 41377
rect 41782 37433 41834 37439
rect 41782 37375 41834 37381
rect 41794 37217 41822 37375
rect 41782 37211 41834 37217
rect 41782 37153 41834 37159
rect 41590 29441 41642 29447
rect 41590 29383 41642 29389
rect 41494 17453 41546 17459
rect 41494 17395 41546 17401
rect 41398 13901 41450 13907
rect 41398 13843 41450 13849
rect 41014 13013 41066 13019
rect 41014 12955 41066 12961
rect 41110 10793 41162 10799
rect 41110 10735 41162 10741
rect 41122 7765 41150 10735
rect 41110 7759 41162 7765
rect 41110 7701 41162 7707
rect 41110 7463 41162 7469
rect 41110 7405 41162 7411
rect 40630 7167 40682 7173
rect 40630 7109 40682 7115
rect 40054 7093 40106 7099
rect 40054 7035 40106 7041
rect 40342 6353 40394 6359
rect 40342 6295 40394 6301
rect 40150 5021 40202 5027
rect 40150 4963 40202 4969
rect 40162 4139 40190 4963
rect 40150 4133 40202 4139
rect 40150 4075 40202 4081
rect 40246 3689 40298 3695
rect 40246 3631 40298 3637
rect 40054 3615 40106 3621
rect 40054 3557 40106 3563
rect 39958 1765 40010 1771
rect 39958 1707 40010 1713
rect 40066 800 40094 3557
rect 40258 1864 40286 3631
rect 40162 1836 40286 1864
rect 40162 800 40190 1836
rect 40246 1765 40298 1771
rect 40246 1707 40298 1713
rect 40258 800 40286 1707
rect 40354 800 40382 6295
rect 40534 3023 40586 3029
rect 40534 2965 40586 2971
rect 40546 800 40574 2965
rect 40642 800 40670 7109
rect 40726 5687 40778 5693
rect 40726 5629 40778 5635
rect 40738 800 40766 5629
rect 40918 5021 40970 5027
rect 40918 4963 40970 4969
rect 40930 3917 40958 4963
rect 40918 3911 40970 3917
rect 40918 3853 40970 3859
rect 41014 3689 41066 3695
rect 41014 3631 41066 3637
rect 41026 3233 41054 3631
rect 40930 3205 41054 3233
rect 40930 800 40958 3205
rect 41122 3048 41150 7405
rect 41506 7099 41534 17395
rect 41878 13087 41930 13093
rect 41878 13029 41930 13035
rect 41890 7765 41918 13029
rect 41878 7759 41930 7765
rect 41878 7701 41930 7707
rect 41686 7537 41738 7543
rect 41686 7479 41738 7485
rect 41494 7093 41546 7099
rect 41494 7035 41546 7041
rect 41590 6945 41642 6951
rect 41590 6887 41642 6893
rect 41494 6353 41546 6359
rect 41494 6295 41546 6301
rect 41302 5021 41354 5027
rect 41302 4963 41354 4969
rect 41206 3911 41258 3917
rect 41206 3853 41258 3859
rect 41218 3251 41246 3853
rect 41314 3621 41342 4963
rect 41398 4281 41450 4287
rect 41398 4223 41450 4229
rect 41302 3615 41354 3621
rect 41302 3557 41354 3563
rect 41206 3245 41258 3251
rect 41206 3187 41258 3193
rect 41026 3020 41150 3048
rect 41026 800 41054 3020
rect 41110 2949 41162 2955
rect 41110 2891 41162 2897
rect 41206 2949 41258 2955
rect 41206 2891 41258 2897
rect 41122 800 41150 2891
rect 41218 800 41246 2891
rect 41410 800 41438 4223
rect 41506 800 41534 6295
rect 41602 4287 41630 6887
rect 41590 4281 41642 4287
rect 41590 4223 41642 4229
rect 41590 3615 41642 3621
rect 41590 3557 41642 3563
rect 41602 800 41630 3557
rect 41698 800 41726 7479
rect 42082 6507 42110 41371
rect 42262 14567 42314 14573
rect 42262 14509 42314 14515
rect 42274 8579 42302 14509
rect 42562 9615 42590 55505
rect 42850 32185 42878 56763
rect 42934 37507 42986 37513
rect 42934 37449 42986 37455
rect 42946 36773 42974 37449
rect 42934 36767 42986 36773
rect 42934 36709 42986 36715
rect 42838 32179 42890 32185
rect 42838 32121 42890 32127
rect 42934 13013 42986 13019
rect 42934 12955 42986 12961
rect 42646 12199 42698 12205
rect 42646 12141 42698 12147
rect 42550 9609 42602 9615
rect 42550 9551 42602 9557
rect 42262 8573 42314 8579
rect 42262 8515 42314 8521
rect 42358 8277 42410 8283
rect 42358 8219 42410 8225
rect 42070 6501 42122 6507
rect 42070 6443 42122 6449
rect 41878 6353 41930 6359
rect 41878 6295 41930 6301
rect 41890 800 41918 6295
rect 41974 4355 42026 4361
rect 41974 4297 42026 4303
rect 42262 4355 42314 4361
rect 42262 4297 42314 4303
rect 41986 800 42014 4297
rect 42070 4281 42122 4287
rect 42070 4223 42122 4229
rect 42082 800 42110 4223
rect 42166 3245 42218 3251
rect 42166 3187 42218 3193
rect 42178 2012 42206 3187
rect 42274 2160 42302 4297
rect 42370 2456 42398 8219
rect 42658 7765 42686 12141
rect 42646 7759 42698 7765
rect 42646 7701 42698 7707
rect 42946 7099 42974 12955
rect 43042 11761 43070 56837
rect 43330 56531 43358 59200
rect 43906 56531 43934 59200
rect 44386 56975 44414 59200
rect 44374 56969 44426 56975
rect 44374 56911 44426 56917
rect 44962 56531 44990 59200
rect 43318 56525 43370 56531
rect 43318 56467 43370 56473
rect 43894 56525 43946 56531
rect 43894 56467 43946 56473
rect 44950 56525 45002 56531
rect 44950 56467 45002 56473
rect 43414 56229 43466 56235
rect 43414 56171 43466 56177
rect 43894 56229 43946 56235
rect 43894 56171 43946 56177
rect 44758 56229 44810 56235
rect 44758 56171 44810 56177
rect 43030 11755 43082 11761
rect 43030 11697 43082 11703
rect 43426 11243 43454 56171
rect 43702 42243 43754 42249
rect 43702 42185 43754 42191
rect 43414 11237 43466 11243
rect 43414 11179 43466 11185
rect 43714 7913 43742 42185
rect 43906 27079 43934 56171
rect 44470 44759 44522 44765
rect 44470 44701 44522 44707
rect 44374 35435 44426 35441
rect 44374 35377 44426 35383
rect 44386 29891 44414 35377
rect 44374 29885 44426 29891
rect 44374 29827 44426 29833
rect 43894 27073 43946 27079
rect 43894 27015 43946 27021
rect 44086 13161 44138 13167
rect 44086 13103 44138 13109
rect 44098 8579 44126 13103
rect 44086 8573 44138 8579
rect 44086 8515 44138 8521
rect 44278 8277 44330 8283
rect 44278 8219 44330 8225
rect 43702 7907 43754 7913
rect 43702 7849 43754 7855
rect 43222 7463 43274 7469
rect 43222 7405 43274 7411
rect 42934 7093 42986 7099
rect 42934 7035 42986 7041
rect 43126 7093 43178 7099
rect 43126 7035 43178 7041
rect 42742 6871 42794 6877
rect 42742 6813 42794 6819
rect 42598 5650 42650 5656
rect 42598 5592 42650 5598
rect 42610 5471 42638 5592
rect 42598 5465 42650 5471
rect 42598 5407 42650 5413
rect 42454 5021 42506 5027
rect 42454 4963 42506 4969
rect 42466 3103 42494 4963
rect 42754 4824 42782 6813
rect 43030 5835 43082 5841
rect 43030 5777 43082 5783
rect 42886 5650 42938 5656
rect 42886 5592 42938 5598
rect 42898 5416 42926 5592
rect 42898 5388 42974 5416
rect 42754 4796 42878 4824
rect 42550 3837 42602 3843
rect 42550 3779 42602 3785
rect 42454 3097 42506 3103
rect 42454 3039 42506 3045
rect 42454 2801 42506 2807
rect 42454 2743 42506 2749
rect 42466 2585 42494 2743
rect 42454 2579 42506 2585
rect 42454 2521 42506 2527
rect 42370 2428 42494 2456
rect 42274 2132 42398 2160
rect 42178 1984 42302 2012
rect 42274 800 42302 1984
rect 42370 800 42398 2132
rect 42466 800 42494 2428
rect 42562 800 42590 3779
rect 42742 3689 42794 3695
rect 42742 3631 42794 3637
rect 42754 800 42782 3631
rect 42850 800 42878 4796
rect 42946 4509 42974 5388
rect 42934 4503 42986 4509
rect 42934 4445 42986 4451
rect 43042 4435 43070 5777
rect 43030 4429 43082 4435
rect 43030 4371 43082 4377
rect 43138 4287 43166 7035
rect 43126 4281 43178 4287
rect 43126 4223 43178 4229
rect 42934 3097 42986 3103
rect 42934 3039 42986 3045
rect 42946 800 42974 3039
rect 43030 3023 43082 3029
rect 43030 2965 43082 2971
rect 43042 800 43070 2965
rect 43234 800 43262 7405
rect 43798 6945 43850 6951
rect 43798 6887 43850 6893
rect 43606 6797 43658 6803
rect 43606 6739 43658 6745
rect 43318 6353 43370 6359
rect 43318 6295 43370 6301
rect 43330 800 43358 6295
rect 43510 5687 43562 5693
rect 43510 5629 43562 5635
rect 43414 4355 43466 4361
rect 43414 4297 43466 4303
rect 43426 800 43454 4297
rect 43522 3843 43550 5629
rect 43510 3837 43562 3843
rect 43510 3779 43562 3785
rect 43618 800 43646 6739
rect 43810 5249 43838 6887
rect 43798 5243 43850 5249
rect 43798 5185 43850 5191
rect 43894 5021 43946 5027
rect 43894 4963 43946 4969
rect 43990 5021 44042 5027
rect 43990 4963 44042 4969
rect 43798 4133 43850 4139
rect 43798 4075 43850 4081
rect 43702 3911 43754 3917
rect 43702 3853 43754 3859
rect 43714 800 43742 3853
rect 43810 3843 43838 4075
rect 43798 3837 43850 3843
rect 43798 3779 43850 3785
rect 43798 3615 43850 3621
rect 43798 3557 43850 3563
rect 43810 800 43838 3557
rect 43906 3251 43934 4963
rect 43894 3245 43946 3251
rect 43894 3187 43946 3193
rect 44002 3103 44030 4963
rect 44086 4281 44138 4287
rect 44086 4223 44138 4229
rect 43990 3097 44042 3103
rect 43990 3039 44042 3045
rect 43894 2949 43946 2955
rect 43894 2891 43946 2897
rect 43906 800 43934 2891
rect 44098 800 44126 4223
rect 44290 3219 44318 8219
rect 44482 7913 44510 44701
rect 44770 43214 44798 56171
rect 45442 55717 45470 59200
rect 45922 56901 45950 59200
rect 45910 56895 45962 56901
rect 45910 56837 45962 56843
rect 46102 56747 46154 56753
rect 46102 56689 46154 56695
rect 45430 55711 45482 55717
rect 45430 55653 45482 55659
rect 45526 55563 45578 55569
rect 45526 55505 45578 55511
rect 45538 43214 45566 55505
rect 44770 43186 44894 43214
rect 45538 43186 45662 43214
rect 44866 30280 44894 43186
rect 45334 39431 45386 39437
rect 45334 39373 45386 39379
rect 45190 30551 45242 30557
rect 45190 30493 45242 30499
rect 45202 30372 45230 30493
rect 45190 30366 45242 30372
rect 45190 30308 45242 30314
rect 44770 30252 44894 30280
rect 44614 30181 44666 30187
rect 44614 30123 44666 30129
rect 44626 29984 44654 30123
rect 44626 29956 44702 29984
rect 44566 29885 44618 29891
rect 44566 29827 44618 29833
rect 44470 7907 44522 7913
rect 44470 7849 44522 7855
rect 44374 7463 44426 7469
rect 44374 7405 44426 7411
rect 44276 3210 44332 3219
rect 44276 3145 44332 3154
rect 44386 3103 44414 7405
rect 44578 7099 44606 29827
rect 44674 15609 44702 29956
rect 44662 15603 44714 15609
rect 44662 15545 44714 15551
rect 44770 14573 44798 30252
rect 44902 30181 44954 30187
rect 44902 30123 44954 30129
rect 44914 29984 44942 30123
rect 44914 29956 44990 29984
rect 44962 15461 44990 29956
rect 45238 25149 45290 25155
rect 45238 25091 45290 25097
rect 44950 15455 45002 15461
rect 44950 15397 45002 15403
rect 44758 14567 44810 14573
rect 44758 14509 44810 14515
rect 45250 7913 45278 25091
rect 45346 10133 45374 39373
rect 45634 29984 45662 43186
rect 45718 33437 45770 33443
rect 45718 33379 45770 33385
rect 45538 29956 45662 29984
rect 45538 12945 45566 29956
rect 45730 27374 45758 33379
rect 45634 27346 45758 27374
rect 45634 13093 45662 27346
rect 45622 13087 45674 13093
rect 45622 13029 45674 13035
rect 45526 12939 45578 12945
rect 45526 12881 45578 12887
rect 45334 10127 45386 10133
rect 45334 10069 45386 10075
rect 45622 9461 45674 9467
rect 45622 9403 45674 9409
rect 45238 7907 45290 7913
rect 45238 7849 45290 7855
rect 45430 7537 45482 7543
rect 45430 7479 45482 7485
rect 45046 7463 45098 7469
rect 45046 7405 45098 7411
rect 44566 7093 44618 7099
rect 44566 7035 44618 7041
rect 44758 6353 44810 6359
rect 44758 6295 44810 6301
rect 44662 5687 44714 5693
rect 44662 5629 44714 5635
rect 44674 4287 44702 5629
rect 44662 4281 44714 4287
rect 44662 4223 44714 4229
rect 44470 3837 44522 3843
rect 44470 3779 44522 3785
rect 44374 3097 44426 3103
rect 44374 3039 44426 3045
rect 44182 2949 44234 2955
rect 44182 2891 44234 2897
rect 44276 2914 44332 2923
rect 44194 800 44222 2891
rect 44276 2849 44332 2858
rect 44290 800 44318 2849
rect 44482 800 44510 3779
rect 44566 3541 44618 3547
rect 44566 3483 44618 3489
rect 44578 800 44606 3483
rect 44662 2801 44714 2807
rect 44662 2743 44714 2749
rect 44674 800 44702 2743
rect 44770 800 44798 6295
rect 44854 5021 44906 5027
rect 44854 4963 44906 4969
rect 44866 3917 44894 4963
rect 44950 4355 45002 4361
rect 44950 4297 45002 4303
rect 44854 3911 44906 3917
rect 44854 3853 44906 3859
rect 44962 800 44990 4297
rect 45058 2807 45086 7405
rect 45334 6205 45386 6211
rect 45334 6147 45386 6153
rect 45238 3763 45290 3769
rect 45238 3705 45290 3711
rect 45142 3245 45194 3251
rect 45142 3187 45194 3193
rect 45046 2801 45098 2807
rect 45046 2743 45098 2749
rect 45046 2431 45098 2437
rect 45046 2373 45098 2379
rect 45058 800 45086 2373
rect 45154 800 45182 3187
rect 45250 800 45278 3705
rect 45346 3103 45374 6147
rect 45334 3097 45386 3103
rect 45334 3039 45386 3045
rect 45442 800 45470 7479
rect 45634 7025 45662 9403
rect 46114 9171 46142 56689
rect 46498 56531 46526 59200
rect 46486 56525 46538 56531
rect 46486 56467 46538 56473
rect 46198 56451 46250 56457
rect 46198 56393 46250 56399
rect 46210 50093 46238 56393
rect 46294 56303 46346 56309
rect 46294 56245 46346 56251
rect 46198 50087 46250 50093
rect 46198 50029 46250 50035
rect 46306 48761 46334 56245
rect 46774 56229 46826 56235
rect 46774 56171 46826 56177
rect 46786 49575 46814 56171
rect 46978 55717 47006 59200
rect 47554 56975 47582 59200
rect 47542 56969 47594 56975
rect 47542 56911 47594 56917
rect 48034 56531 48062 59200
rect 48610 56531 48638 59200
rect 49090 56975 49118 59200
rect 49078 56969 49130 56975
rect 49078 56911 49130 56917
rect 48886 56895 48938 56901
rect 48886 56837 48938 56843
rect 48022 56525 48074 56531
rect 48022 56467 48074 56473
rect 48598 56525 48650 56531
rect 48598 56467 48650 56473
rect 48310 56377 48362 56383
rect 48310 56319 48362 56325
rect 47830 56229 47882 56235
rect 47830 56171 47882 56177
rect 46966 55711 47018 55717
rect 46966 55653 47018 55659
rect 46966 55415 47018 55421
rect 46966 55357 47018 55363
rect 46774 49569 46826 49575
rect 46774 49511 46826 49517
rect 46294 48755 46346 48761
rect 46294 48697 46346 48703
rect 46678 39579 46730 39585
rect 46678 39521 46730 39527
rect 46690 39308 46718 39521
rect 46690 39280 46862 39308
rect 46834 39141 46862 39280
rect 46822 39135 46874 39141
rect 46822 39077 46874 39083
rect 46870 38765 46922 38771
rect 46870 38707 46922 38713
rect 46390 26925 46442 26931
rect 46390 26867 46442 26873
rect 46102 9165 46154 9171
rect 46102 9107 46154 9113
rect 46402 7765 46430 26867
rect 46774 21005 46826 21011
rect 46774 20947 46826 20953
rect 46582 18119 46634 18125
rect 46582 18061 46634 18067
rect 46390 7759 46442 7765
rect 46390 7701 46442 7707
rect 46390 7463 46442 7469
rect 46390 7405 46442 7411
rect 45622 7019 45674 7025
rect 45622 6961 45674 6967
rect 45814 6945 45866 6951
rect 45814 6887 45866 6893
rect 45718 6871 45770 6877
rect 45718 6813 45770 6819
rect 45526 6353 45578 6359
rect 45526 6295 45578 6301
rect 45538 800 45566 6295
rect 45622 5021 45674 5027
rect 45622 4963 45674 4969
rect 45634 3843 45662 4963
rect 45622 3837 45674 3843
rect 45622 3779 45674 3785
rect 45622 3023 45674 3029
rect 45622 2965 45674 2971
rect 45634 800 45662 2965
rect 45730 2308 45758 6813
rect 45826 2437 45854 6887
rect 46102 5687 46154 5693
rect 46102 5629 46154 5635
rect 46114 4269 46142 5629
rect 46402 4269 46430 7405
rect 46594 7099 46622 18061
rect 46786 9560 46814 20947
rect 46882 12974 46910 38707
rect 46978 33134 47006 55357
rect 47254 50457 47306 50463
rect 47254 50399 47306 50405
rect 47266 50093 47294 50399
rect 47254 50087 47306 50093
rect 47254 50029 47306 50035
rect 47266 33134 47294 50029
rect 47542 39505 47594 39511
rect 47542 39447 47594 39453
rect 47554 39215 47582 39447
rect 47542 39209 47594 39215
rect 47542 39151 47594 39157
rect 46978 33106 47102 33134
rect 47266 33106 47390 33134
rect 47074 17294 47102 33106
rect 47074 17266 47198 17294
rect 47170 12974 47198 17266
rect 46882 12946 47006 12974
rect 46786 9532 46910 9560
rect 46774 9461 46826 9467
rect 46774 9403 46826 9409
rect 46786 9245 46814 9403
rect 46774 9239 46826 9245
rect 46774 9181 46826 9187
rect 46882 7913 46910 9532
rect 46870 7907 46922 7913
rect 46870 7849 46922 7855
rect 46870 7537 46922 7543
rect 46870 7479 46922 7485
rect 46582 7093 46634 7099
rect 46582 7035 46634 7041
rect 46486 7019 46538 7025
rect 46486 6961 46538 6967
rect 46498 5120 46526 6961
rect 46678 5687 46730 5693
rect 46678 5629 46730 5635
rect 46498 5092 46622 5120
rect 46486 5021 46538 5027
rect 46486 4963 46538 4969
rect 45922 4241 46142 4269
rect 46210 4241 46430 4269
rect 45814 2431 45866 2437
rect 45814 2373 45866 2379
rect 45730 2280 45854 2308
rect 45826 800 45854 2280
rect 45922 800 45950 4241
rect 46006 3615 46058 3621
rect 46006 3557 46058 3563
rect 46018 800 46046 3557
rect 46210 2894 46238 4241
rect 46294 3911 46346 3917
rect 46294 3853 46346 3859
rect 46114 2866 46238 2894
rect 46114 800 46142 2866
rect 46306 800 46334 3853
rect 46498 3251 46526 4963
rect 46486 3245 46538 3251
rect 46486 3187 46538 3193
rect 46594 3085 46622 5092
rect 46498 3057 46622 3085
rect 46390 2949 46442 2955
rect 46390 2891 46442 2897
rect 46402 800 46430 2891
rect 46498 800 46526 3057
rect 46690 2894 46718 5629
rect 46774 4355 46826 4361
rect 46774 4297 46826 4303
rect 46594 2866 46718 2894
rect 46594 800 46622 2866
rect 46786 800 46814 4297
rect 46882 800 46910 7479
rect 46978 6507 47006 12946
rect 47074 12946 47198 12974
rect 46966 6501 47018 6507
rect 46966 6443 47018 6449
rect 46966 6353 47018 6359
rect 46966 6295 47018 6301
rect 46978 800 47006 6295
rect 47074 5101 47102 12946
rect 47158 10127 47210 10133
rect 47158 10069 47210 10075
rect 47170 7099 47198 10069
rect 47158 7093 47210 7099
rect 47158 7035 47210 7041
rect 47254 6871 47306 6877
rect 47254 6813 47306 6819
rect 47158 6501 47210 6507
rect 47158 6443 47210 6449
rect 47062 5095 47114 5101
rect 47062 5037 47114 5043
rect 47170 4139 47198 6443
rect 47158 4133 47210 4139
rect 47158 4075 47210 4081
rect 47158 3689 47210 3695
rect 47158 3631 47210 3637
rect 47170 800 47198 3631
rect 47266 800 47294 6813
rect 47362 6433 47390 33106
rect 47734 26259 47786 26265
rect 47734 26201 47786 26207
rect 47746 19013 47774 26201
rect 47734 19007 47786 19013
rect 47734 18949 47786 18955
rect 47842 13611 47870 56171
rect 48322 45727 48350 56319
rect 48598 56229 48650 56235
rect 48598 56171 48650 56177
rect 48310 45721 48362 45727
rect 48310 45663 48362 45669
rect 47926 35435 47978 35441
rect 47926 35377 47978 35383
rect 47830 13605 47882 13611
rect 47830 13547 47882 13553
rect 47830 10275 47882 10281
rect 47830 10217 47882 10223
rect 47638 8277 47690 8283
rect 47638 8219 47690 8225
rect 47350 6427 47402 6433
rect 47350 6369 47402 6375
rect 47542 5687 47594 5693
rect 47542 5629 47594 5635
rect 47554 4380 47582 5629
rect 47362 4352 47582 4380
rect 47362 800 47390 4352
rect 47446 4281 47498 4287
rect 47446 4223 47498 4229
rect 47458 800 47486 4223
rect 47650 800 47678 8219
rect 47842 7765 47870 10217
rect 47938 8431 47966 35377
rect 48214 26851 48266 26857
rect 48214 26793 48266 26799
rect 48118 11681 48170 11687
rect 48118 11623 48170 11629
rect 47926 8425 47978 8431
rect 47926 8367 47978 8373
rect 48022 8277 48074 8283
rect 48022 8219 48074 8225
rect 47830 7759 47882 7765
rect 47830 7701 47882 7707
rect 47734 6353 47786 6359
rect 47734 6295 47786 6301
rect 47746 800 47774 6295
rect 47926 5021 47978 5027
rect 47926 4963 47978 4969
rect 47830 4355 47882 4361
rect 47830 4297 47882 4303
rect 47842 800 47870 4297
rect 47938 3917 47966 4963
rect 47926 3911 47978 3917
rect 47926 3853 47978 3859
rect 48034 800 48062 8219
rect 48130 7099 48158 11623
rect 48226 8579 48254 26793
rect 48610 9911 48638 56171
rect 48898 31815 48926 56837
rect 49666 56531 49694 59200
rect 50146 56531 50174 59200
rect 50722 56975 50750 59200
rect 50710 56969 50762 56975
rect 50710 56911 50762 56917
rect 50902 56895 50954 56901
rect 50902 56837 50954 56843
rect 50348 56638 50644 56658
rect 50404 56636 50428 56638
rect 50484 56636 50508 56638
rect 50564 56636 50588 56638
rect 50426 56584 50428 56636
rect 50490 56584 50502 56636
rect 50564 56584 50566 56636
rect 50404 56582 50428 56584
rect 50484 56582 50508 56584
rect 50564 56582 50588 56584
rect 50348 56562 50644 56582
rect 49654 56525 49706 56531
rect 49654 56467 49706 56473
rect 50134 56525 50186 56531
rect 50134 56467 50186 56473
rect 50038 56303 50090 56309
rect 50038 56245 50090 56251
rect 49654 53417 49706 53423
rect 49654 53359 49706 53365
rect 48982 45129 49034 45135
rect 48982 45071 49034 45077
rect 48886 31809 48938 31815
rect 48886 31751 48938 31757
rect 48598 9905 48650 9911
rect 48598 9847 48650 9853
rect 48214 8573 48266 8579
rect 48214 8515 48266 8521
rect 48694 8277 48746 8283
rect 48694 8219 48746 8225
rect 48310 7463 48362 7469
rect 48310 7405 48362 7411
rect 48118 7093 48170 7099
rect 48118 7035 48170 7041
rect 48118 4207 48170 4213
rect 48118 4149 48170 4155
rect 48130 800 48158 4149
rect 48214 3689 48266 3695
rect 48214 3631 48266 3637
rect 48226 800 48254 3631
rect 48322 800 48350 7405
rect 48598 4281 48650 4287
rect 48598 4223 48650 4229
rect 48502 4133 48554 4139
rect 48502 4075 48554 4081
rect 48514 800 48542 4075
rect 48610 800 48638 4223
rect 48706 800 48734 8219
rect 48994 7913 49022 45071
rect 49366 22781 49418 22787
rect 49366 22723 49418 22729
rect 49078 19451 49130 19457
rect 49078 19393 49130 19399
rect 48982 7907 49034 7913
rect 48982 7849 49034 7855
rect 49090 7099 49118 19393
rect 49174 8943 49226 8949
rect 49174 8885 49226 8891
rect 49078 7093 49130 7099
rect 49078 7035 49130 7041
rect 49186 6803 49214 8885
rect 49378 8431 49406 22723
rect 49666 10133 49694 53359
rect 50050 46097 50078 56245
rect 50230 56229 50282 56235
rect 50230 56171 50282 56177
rect 50038 46091 50090 46097
rect 50038 46033 50090 46039
rect 49750 43723 49802 43729
rect 49750 43665 49802 43671
rect 49654 10127 49706 10133
rect 49654 10069 49706 10075
rect 49366 8425 49418 8431
rect 49366 8367 49418 8373
rect 49462 8277 49514 8283
rect 49462 8219 49514 8225
rect 49174 6797 49226 6803
rect 49174 6739 49226 6745
rect 48790 6353 48842 6359
rect 48790 6295 48842 6301
rect 48802 800 48830 6295
rect 48982 5687 49034 5693
rect 48982 5629 49034 5635
rect 48994 4213 49022 5629
rect 49366 5021 49418 5027
rect 49366 4963 49418 4969
rect 49174 4355 49226 4361
rect 49174 4297 49226 4303
rect 48982 4207 49034 4213
rect 48982 4149 49034 4155
rect 49186 3640 49214 4297
rect 49270 3911 49322 3917
rect 49270 3853 49322 3859
rect 48994 3612 49214 3640
rect 48994 800 49022 3612
rect 49078 3541 49130 3547
rect 49078 3483 49130 3489
rect 49090 800 49118 3483
rect 49282 2894 49310 3853
rect 49186 2866 49310 2894
rect 49186 800 49214 2866
rect 49378 800 49406 4963
rect 49474 800 49502 8219
rect 49762 7913 49790 43665
rect 49942 19007 49994 19013
rect 49942 18949 49994 18955
rect 49750 7907 49802 7913
rect 49750 7849 49802 7855
rect 49954 7099 49982 18949
rect 50134 13013 50186 13019
rect 50134 12955 50186 12961
rect 50146 8431 50174 12955
rect 50242 12131 50270 56171
rect 50348 55306 50644 55326
rect 50404 55304 50428 55306
rect 50484 55304 50508 55306
rect 50564 55304 50588 55306
rect 50426 55252 50428 55304
rect 50490 55252 50502 55304
rect 50564 55252 50566 55304
rect 50404 55250 50428 55252
rect 50484 55250 50508 55252
rect 50564 55250 50588 55252
rect 50348 55230 50644 55250
rect 50348 53974 50644 53994
rect 50404 53972 50428 53974
rect 50484 53972 50508 53974
rect 50564 53972 50588 53974
rect 50426 53920 50428 53972
rect 50490 53920 50502 53972
rect 50564 53920 50566 53972
rect 50404 53918 50428 53920
rect 50484 53918 50508 53920
rect 50564 53918 50588 53920
rect 50348 53898 50644 53918
rect 50348 52642 50644 52662
rect 50404 52640 50428 52642
rect 50484 52640 50508 52642
rect 50564 52640 50588 52642
rect 50426 52588 50428 52640
rect 50490 52588 50502 52640
rect 50564 52588 50566 52640
rect 50404 52586 50428 52588
rect 50484 52586 50508 52588
rect 50564 52586 50588 52588
rect 50348 52566 50644 52586
rect 50348 51310 50644 51330
rect 50404 51308 50428 51310
rect 50484 51308 50508 51310
rect 50564 51308 50588 51310
rect 50426 51256 50428 51308
rect 50490 51256 50502 51308
rect 50564 51256 50566 51308
rect 50404 51254 50428 51256
rect 50484 51254 50508 51256
rect 50564 51254 50588 51256
rect 50348 51234 50644 51254
rect 50348 49978 50644 49998
rect 50404 49976 50428 49978
rect 50484 49976 50508 49978
rect 50564 49976 50588 49978
rect 50426 49924 50428 49976
rect 50490 49924 50502 49976
rect 50564 49924 50566 49976
rect 50404 49922 50428 49924
rect 50484 49922 50508 49924
rect 50564 49922 50588 49924
rect 50348 49902 50644 49922
rect 50348 48646 50644 48666
rect 50404 48644 50428 48646
rect 50484 48644 50508 48646
rect 50564 48644 50588 48646
rect 50426 48592 50428 48644
rect 50490 48592 50502 48644
rect 50564 48592 50566 48644
rect 50404 48590 50428 48592
rect 50484 48590 50508 48592
rect 50564 48590 50588 48592
rect 50348 48570 50644 48590
rect 50348 47314 50644 47334
rect 50404 47312 50428 47314
rect 50484 47312 50508 47314
rect 50564 47312 50588 47314
rect 50426 47260 50428 47312
rect 50490 47260 50502 47312
rect 50564 47260 50566 47312
rect 50404 47258 50428 47260
rect 50484 47258 50508 47260
rect 50564 47258 50588 47260
rect 50348 47238 50644 47258
rect 50348 45982 50644 46002
rect 50404 45980 50428 45982
rect 50484 45980 50508 45982
rect 50564 45980 50588 45982
rect 50426 45928 50428 45980
rect 50490 45928 50502 45980
rect 50564 45928 50566 45980
rect 50404 45926 50428 45928
rect 50484 45926 50508 45928
rect 50564 45926 50588 45928
rect 50348 45906 50644 45926
rect 50348 44650 50644 44670
rect 50404 44648 50428 44650
rect 50484 44648 50508 44650
rect 50564 44648 50588 44650
rect 50426 44596 50428 44648
rect 50490 44596 50502 44648
rect 50564 44596 50566 44648
rect 50404 44594 50428 44596
rect 50484 44594 50508 44596
rect 50564 44594 50588 44596
rect 50348 44574 50644 44594
rect 50348 43318 50644 43338
rect 50404 43316 50428 43318
rect 50484 43316 50508 43318
rect 50564 43316 50588 43318
rect 50426 43264 50428 43316
rect 50490 43264 50502 43316
rect 50564 43264 50566 43316
rect 50404 43262 50428 43264
rect 50484 43262 50508 43264
rect 50564 43262 50588 43264
rect 50348 43242 50644 43262
rect 50348 41986 50644 42006
rect 50404 41984 50428 41986
rect 50484 41984 50508 41986
rect 50564 41984 50588 41986
rect 50426 41932 50428 41984
rect 50490 41932 50502 41984
rect 50564 41932 50566 41984
rect 50404 41930 50428 41932
rect 50484 41930 50508 41932
rect 50564 41930 50588 41932
rect 50348 41910 50644 41930
rect 50348 40654 50644 40674
rect 50404 40652 50428 40654
rect 50484 40652 50508 40654
rect 50564 40652 50588 40654
rect 50426 40600 50428 40652
rect 50490 40600 50502 40652
rect 50564 40600 50566 40652
rect 50404 40598 50428 40600
rect 50484 40598 50508 40600
rect 50564 40598 50588 40600
rect 50348 40578 50644 40598
rect 50348 39322 50644 39342
rect 50404 39320 50428 39322
rect 50484 39320 50508 39322
rect 50564 39320 50588 39322
rect 50426 39268 50428 39320
rect 50490 39268 50502 39320
rect 50564 39268 50566 39320
rect 50404 39266 50428 39268
rect 50484 39266 50508 39268
rect 50564 39266 50588 39268
rect 50348 39246 50644 39266
rect 50348 37990 50644 38010
rect 50404 37988 50428 37990
rect 50484 37988 50508 37990
rect 50564 37988 50588 37990
rect 50426 37936 50428 37988
rect 50490 37936 50502 37988
rect 50564 37936 50566 37988
rect 50404 37934 50428 37936
rect 50484 37934 50508 37936
rect 50564 37934 50588 37936
rect 50348 37914 50644 37934
rect 50348 36658 50644 36678
rect 50404 36656 50428 36658
rect 50484 36656 50508 36658
rect 50564 36656 50588 36658
rect 50426 36604 50428 36656
rect 50490 36604 50502 36656
rect 50564 36604 50566 36656
rect 50404 36602 50428 36604
rect 50484 36602 50508 36604
rect 50564 36602 50588 36604
rect 50348 36582 50644 36602
rect 50348 35326 50644 35346
rect 50404 35324 50428 35326
rect 50484 35324 50508 35326
rect 50564 35324 50588 35326
rect 50426 35272 50428 35324
rect 50490 35272 50502 35324
rect 50564 35272 50566 35324
rect 50404 35270 50428 35272
rect 50484 35270 50508 35272
rect 50564 35270 50588 35272
rect 50348 35250 50644 35270
rect 50348 33994 50644 34014
rect 50404 33992 50428 33994
rect 50484 33992 50508 33994
rect 50564 33992 50588 33994
rect 50426 33940 50428 33992
rect 50490 33940 50502 33992
rect 50564 33940 50566 33992
rect 50404 33938 50428 33940
rect 50484 33938 50508 33940
rect 50564 33938 50588 33940
rect 50348 33918 50644 33938
rect 50348 32662 50644 32682
rect 50404 32660 50428 32662
rect 50484 32660 50508 32662
rect 50564 32660 50588 32662
rect 50426 32608 50428 32660
rect 50490 32608 50502 32660
rect 50564 32608 50566 32660
rect 50404 32606 50428 32608
rect 50484 32606 50508 32608
rect 50564 32606 50588 32608
rect 50348 32586 50644 32606
rect 50914 32259 50942 56837
rect 51202 56161 51230 59200
rect 51670 56229 51722 56235
rect 51670 56171 51722 56177
rect 51190 56155 51242 56161
rect 51190 56097 51242 56103
rect 51574 46757 51626 46763
rect 51574 46699 51626 46705
rect 51190 35435 51242 35441
rect 51190 35377 51242 35383
rect 51202 35219 51230 35377
rect 51190 35213 51242 35219
rect 51190 35155 51242 35161
rect 50902 32253 50954 32259
rect 50902 32195 50954 32201
rect 50348 31330 50644 31350
rect 50404 31328 50428 31330
rect 50484 31328 50508 31330
rect 50564 31328 50588 31330
rect 50426 31276 50428 31328
rect 50490 31276 50502 31328
rect 50564 31276 50566 31328
rect 50404 31274 50428 31276
rect 50484 31274 50508 31276
rect 50564 31274 50588 31276
rect 50348 31254 50644 31274
rect 51094 30329 51146 30335
rect 51094 30271 51146 30277
rect 50348 29998 50644 30018
rect 50404 29996 50428 29998
rect 50484 29996 50508 29998
rect 50564 29996 50588 29998
rect 50426 29944 50428 29996
rect 50490 29944 50502 29996
rect 50564 29944 50566 29996
rect 50404 29942 50428 29944
rect 50484 29942 50508 29944
rect 50564 29942 50588 29944
rect 50348 29922 50644 29942
rect 50348 28666 50644 28686
rect 50404 28664 50428 28666
rect 50484 28664 50508 28666
rect 50564 28664 50588 28666
rect 50426 28612 50428 28664
rect 50490 28612 50502 28664
rect 50564 28612 50566 28664
rect 50404 28610 50428 28612
rect 50484 28610 50508 28612
rect 50564 28610 50588 28612
rect 50348 28590 50644 28610
rect 50348 27334 50644 27354
rect 50404 27332 50428 27334
rect 50484 27332 50508 27334
rect 50564 27332 50588 27334
rect 50426 27280 50428 27332
rect 50490 27280 50502 27332
rect 50564 27280 50566 27332
rect 50404 27278 50428 27280
rect 50484 27278 50508 27280
rect 50564 27278 50588 27280
rect 50348 27258 50644 27278
rect 50348 26002 50644 26022
rect 50404 26000 50428 26002
rect 50484 26000 50508 26002
rect 50564 26000 50588 26002
rect 50426 25948 50428 26000
rect 50490 25948 50502 26000
rect 50564 25948 50566 26000
rect 50404 25946 50428 25948
rect 50484 25946 50508 25948
rect 50564 25946 50588 25948
rect 50348 25926 50644 25946
rect 50348 24670 50644 24690
rect 50404 24668 50428 24670
rect 50484 24668 50508 24670
rect 50564 24668 50588 24670
rect 50426 24616 50428 24668
rect 50490 24616 50502 24668
rect 50564 24616 50566 24668
rect 50404 24614 50428 24616
rect 50484 24614 50508 24616
rect 50564 24614 50588 24616
rect 50348 24594 50644 24614
rect 50348 23338 50644 23358
rect 50404 23336 50428 23338
rect 50484 23336 50508 23338
rect 50564 23336 50588 23338
rect 50426 23284 50428 23336
rect 50490 23284 50502 23336
rect 50564 23284 50566 23336
rect 50404 23282 50428 23284
rect 50484 23282 50508 23284
rect 50564 23282 50588 23284
rect 50348 23262 50644 23282
rect 50348 22006 50644 22026
rect 50404 22004 50428 22006
rect 50484 22004 50508 22006
rect 50564 22004 50588 22006
rect 50426 21952 50428 22004
rect 50490 21952 50502 22004
rect 50564 21952 50566 22004
rect 50404 21950 50428 21952
rect 50484 21950 50508 21952
rect 50564 21950 50588 21952
rect 50348 21930 50644 21950
rect 50348 20674 50644 20694
rect 50404 20672 50428 20674
rect 50484 20672 50508 20674
rect 50564 20672 50588 20674
rect 50426 20620 50428 20672
rect 50490 20620 50502 20672
rect 50564 20620 50566 20672
rect 50404 20618 50428 20620
rect 50484 20618 50508 20620
rect 50564 20618 50588 20620
rect 50348 20598 50644 20618
rect 50348 19342 50644 19362
rect 50404 19340 50428 19342
rect 50484 19340 50508 19342
rect 50564 19340 50588 19342
rect 50426 19288 50428 19340
rect 50490 19288 50502 19340
rect 50564 19288 50566 19340
rect 50404 19286 50428 19288
rect 50484 19286 50508 19288
rect 50564 19286 50588 19288
rect 50348 19266 50644 19286
rect 50348 18010 50644 18030
rect 50404 18008 50428 18010
rect 50484 18008 50508 18010
rect 50564 18008 50588 18010
rect 50426 17956 50428 18008
rect 50490 17956 50502 18008
rect 50564 17956 50566 18008
rect 50404 17954 50428 17956
rect 50484 17954 50508 17956
rect 50564 17954 50588 17956
rect 50348 17934 50644 17954
rect 51106 17294 51134 30271
rect 51478 25223 51530 25229
rect 51478 25165 51530 25171
rect 51106 17266 51230 17294
rect 50348 16678 50644 16698
rect 50404 16676 50428 16678
rect 50484 16676 50508 16678
rect 50564 16676 50588 16678
rect 50426 16624 50428 16676
rect 50490 16624 50502 16676
rect 50564 16624 50566 16676
rect 50404 16622 50428 16624
rect 50484 16622 50508 16624
rect 50564 16622 50588 16624
rect 50348 16602 50644 16622
rect 50348 15346 50644 15366
rect 50404 15344 50428 15346
rect 50484 15344 50508 15346
rect 50564 15344 50588 15346
rect 50426 15292 50428 15344
rect 50490 15292 50502 15344
rect 50564 15292 50566 15344
rect 50404 15290 50428 15292
rect 50484 15290 50508 15292
rect 50564 15290 50588 15292
rect 50348 15270 50644 15290
rect 50348 14014 50644 14034
rect 50404 14012 50428 14014
rect 50484 14012 50508 14014
rect 50564 14012 50588 14014
rect 50426 13960 50428 14012
rect 50490 13960 50502 14012
rect 50564 13960 50566 14012
rect 50404 13958 50428 13960
rect 50484 13958 50508 13960
rect 50564 13958 50588 13960
rect 50348 13938 50644 13958
rect 50348 12682 50644 12702
rect 50404 12680 50428 12682
rect 50484 12680 50508 12682
rect 50564 12680 50588 12682
rect 50426 12628 50428 12680
rect 50490 12628 50502 12680
rect 50564 12628 50566 12680
rect 50404 12626 50428 12628
rect 50484 12626 50508 12628
rect 50564 12626 50588 12628
rect 50348 12606 50644 12626
rect 50230 12125 50282 12131
rect 50230 12067 50282 12073
rect 50348 11350 50644 11370
rect 50404 11348 50428 11350
rect 50484 11348 50508 11350
rect 50564 11348 50588 11350
rect 50426 11296 50428 11348
rect 50490 11296 50502 11348
rect 50564 11296 50566 11348
rect 50404 11294 50428 11296
rect 50484 11294 50508 11296
rect 50564 11294 50588 11296
rect 50348 11274 50644 11294
rect 50710 10127 50762 10133
rect 50710 10069 50762 10075
rect 50348 10018 50644 10038
rect 50404 10016 50428 10018
rect 50484 10016 50508 10018
rect 50564 10016 50588 10018
rect 50426 9964 50428 10016
rect 50490 9964 50502 10016
rect 50564 9964 50566 10016
rect 50404 9962 50428 9964
rect 50484 9962 50508 9964
rect 50564 9962 50588 9964
rect 50348 9942 50644 9962
rect 50348 8686 50644 8706
rect 50404 8684 50428 8686
rect 50484 8684 50508 8686
rect 50564 8684 50588 8686
rect 50426 8632 50428 8684
rect 50490 8632 50502 8684
rect 50564 8632 50566 8684
rect 50404 8630 50428 8632
rect 50484 8630 50508 8632
rect 50564 8630 50588 8632
rect 50348 8610 50644 8630
rect 50134 8425 50186 8431
rect 50134 8367 50186 8373
rect 50038 7463 50090 7469
rect 50038 7405 50090 7411
rect 49942 7093 49994 7099
rect 49942 7035 49994 7041
rect 49558 6353 49610 6359
rect 49558 6295 49610 6301
rect 49570 800 49598 6295
rect 49750 6131 49802 6137
rect 49750 6073 49802 6079
rect 49654 5687 49706 5693
rect 49654 5629 49706 5635
rect 49666 4139 49694 5629
rect 49654 4133 49706 4139
rect 49654 4075 49706 4081
rect 49654 3023 49706 3029
rect 49654 2965 49706 2971
rect 49666 800 49694 2965
rect 49762 2012 49790 6073
rect 49846 4207 49898 4213
rect 49846 4149 49898 4155
rect 49858 2160 49886 4149
rect 50050 3547 50078 7405
rect 50348 7354 50644 7374
rect 50404 7352 50428 7354
rect 50484 7352 50508 7354
rect 50564 7352 50588 7354
rect 50426 7300 50428 7352
rect 50490 7300 50502 7352
rect 50564 7300 50566 7352
rect 50404 7298 50428 7300
rect 50484 7298 50508 7300
rect 50564 7298 50588 7300
rect 50348 7278 50644 7298
rect 50134 6945 50186 6951
rect 50134 6887 50186 6893
rect 50038 3541 50090 3547
rect 50038 3483 50090 3489
rect 49942 2949 49994 2955
rect 49942 2894 49994 2897
rect 49942 2891 50078 2894
rect 49954 2866 50078 2891
rect 49858 2132 49982 2160
rect 49762 1984 49886 2012
rect 49858 800 49886 1984
rect 49954 800 49982 2132
rect 50050 800 50078 2866
rect 50146 800 50174 6887
rect 50722 6581 50750 10069
rect 51094 8129 51146 8135
rect 51094 8071 51146 8077
rect 51106 7765 51134 8071
rect 51094 7759 51146 7765
rect 51094 7701 51146 7707
rect 50710 6575 50762 6581
rect 50710 6517 50762 6523
rect 51202 6285 51230 17266
rect 51286 6945 51338 6951
rect 51286 6887 51338 6893
rect 51190 6279 51242 6285
rect 51190 6221 51242 6227
rect 51094 6131 51146 6137
rect 51094 6073 51146 6079
rect 50348 6022 50644 6042
rect 50404 6020 50428 6022
rect 50484 6020 50508 6022
rect 50564 6020 50588 6022
rect 50426 5968 50428 6020
rect 50490 5968 50502 6020
rect 50564 5968 50566 6020
rect 50404 5966 50428 5968
rect 50484 5966 50508 5968
rect 50564 5966 50588 5968
rect 50348 5946 50644 5966
rect 50710 5687 50762 5693
rect 50710 5629 50762 5635
rect 50422 5021 50474 5027
rect 50422 4963 50474 4969
rect 50434 4824 50462 4963
rect 50242 4796 50462 4824
rect 50242 2604 50270 4796
rect 50348 4690 50644 4710
rect 50404 4688 50428 4690
rect 50484 4688 50508 4690
rect 50564 4688 50588 4690
rect 50426 4636 50428 4688
rect 50490 4636 50502 4688
rect 50564 4636 50566 4688
rect 50404 4634 50428 4636
rect 50484 4634 50508 4636
rect 50564 4634 50588 4636
rect 50348 4614 50644 4634
rect 50722 3917 50750 5629
rect 50902 5021 50954 5027
rect 50902 4963 50954 4969
rect 50710 3911 50762 3917
rect 50710 3853 50762 3859
rect 50710 3689 50762 3695
rect 50710 3631 50762 3637
rect 50806 3689 50858 3695
rect 50806 3631 50858 3637
rect 50348 3358 50644 3378
rect 50404 3356 50428 3358
rect 50484 3356 50508 3358
rect 50564 3356 50588 3358
rect 50426 3304 50428 3356
rect 50490 3304 50502 3356
rect 50564 3304 50566 3356
rect 50404 3302 50428 3304
rect 50484 3302 50508 3304
rect 50564 3302 50588 3304
rect 50348 3282 50644 3302
rect 50242 2576 50366 2604
rect 50338 800 50366 2576
rect 50722 1864 50750 3631
rect 50434 1836 50750 1864
rect 50434 800 50462 1836
rect 50710 1765 50762 1771
rect 50710 1707 50762 1713
rect 50518 1691 50570 1697
rect 50518 1633 50570 1639
rect 50530 800 50558 1633
rect 50722 800 50750 1707
rect 50818 800 50846 3631
rect 50914 1771 50942 4963
rect 50998 4281 51050 4287
rect 50998 4223 51050 4229
rect 50902 1765 50954 1771
rect 50902 1707 50954 1713
rect 50902 1617 50954 1623
rect 50902 1559 50954 1565
rect 50914 800 50942 1559
rect 51010 800 51038 4223
rect 51106 1697 51134 6073
rect 51190 3541 51242 3547
rect 51190 3483 51242 3489
rect 51094 1691 51146 1697
rect 51094 1633 51146 1639
rect 51202 800 51230 3483
rect 51298 800 51326 6887
rect 51490 6433 51518 25165
rect 51586 12205 51614 46699
rect 51574 12199 51626 12205
rect 51574 12141 51626 12147
rect 51682 8801 51710 56171
rect 51778 55717 51806 59200
rect 52258 56901 52286 59200
rect 52834 57614 52862 59200
rect 52834 57586 52958 57614
rect 52246 56895 52298 56901
rect 52246 56837 52298 56843
rect 52822 56747 52874 56753
rect 52822 56689 52874 56695
rect 51766 55711 51818 55717
rect 51766 55653 51818 55659
rect 52054 55563 52106 55569
rect 52054 55505 52106 55511
rect 52066 40325 52094 55505
rect 52438 50235 52490 50241
rect 52438 50177 52490 50183
rect 52054 40319 52106 40325
rect 52054 40261 52106 40267
rect 52342 28849 52394 28855
rect 52342 28791 52394 28797
rect 52054 13827 52106 13833
rect 52054 13769 52106 13775
rect 51670 8795 51722 8801
rect 51670 8737 51722 8743
rect 51670 7463 51722 7469
rect 51670 7405 51722 7411
rect 51478 6427 51530 6433
rect 51478 6369 51530 6375
rect 51574 6353 51626 6359
rect 51574 6295 51626 6301
rect 51382 3911 51434 3917
rect 51382 3853 51434 3859
rect 51394 800 51422 3853
rect 51478 3023 51530 3029
rect 51478 2965 51530 2971
rect 51490 800 51518 2965
rect 51586 1623 51614 6295
rect 51574 1617 51626 1623
rect 51574 1559 51626 1565
rect 51682 800 51710 7405
rect 52066 7099 52094 13769
rect 52354 8579 52382 28791
rect 52342 8573 52394 8579
rect 52342 8515 52394 8521
rect 52342 7463 52394 7469
rect 52342 7405 52394 7411
rect 52054 7093 52106 7099
rect 52054 7035 52106 7041
rect 52150 5687 52202 5693
rect 52150 5629 52202 5635
rect 51862 5021 51914 5027
rect 51862 4963 51914 4969
rect 51958 5021 52010 5027
rect 51958 4963 52010 4969
rect 51874 3917 51902 4963
rect 51862 3911 51914 3917
rect 51862 3853 51914 3859
rect 51970 3788 51998 4963
rect 51778 3760 51998 3788
rect 51778 800 51806 3760
rect 52054 3689 52106 3695
rect 51970 3649 52054 3677
rect 51970 1864 51998 3649
rect 52054 3631 52106 3637
rect 52054 3541 52106 3547
rect 52054 3483 52106 3489
rect 51874 1836 51998 1864
rect 51874 800 51902 1836
rect 52066 800 52094 3483
rect 52162 800 52190 5629
rect 52246 2949 52298 2955
rect 52246 2891 52298 2897
rect 52258 800 52286 2891
rect 52354 800 52382 7405
rect 52450 7099 52478 50177
rect 52534 42761 52586 42767
rect 52534 42703 52586 42709
rect 52546 42545 52574 42703
rect 52534 42539 52586 42545
rect 52534 42481 52586 42487
rect 52834 31889 52862 56689
rect 52930 56531 52958 57586
rect 53314 56531 53342 59200
rect 53890 56975 53918 59200
rect 53878 56969 53930 56975
rect 53878 56911 53930 56917
rect 54370 56531 54398 59200
rect 54838 56821 54890 56827
rect 54838 56763 54890 56769
rect 52918 56525 52970 56531
rect 52918 56467 52970 56473
rect 53302 56525 53354 56531
rect 53302 56467 53354 56473
rect 54358 56525 54410 56531
rect 54358 56467 54410 56473
rect 54850 56383 54878 56763
rect 54946 56531 54974 59200
rect 55426 56975 55454 59200
rect 55414 56969 55466 56975
rect 55414 56911 55466 56917
rect 55702 56747 55754 56753
rect 55702 56689 55754 56695
rect 54934 56525 54986 56531
rect 54934 56467 54986 56473
rect 54838 56377 54890 56383
rect 54838 56319 54890 56325
rect 53398 56229 53450 56235
rect 53398 56171 53450 56177
rect 53410 51573 53438 56171
rect 55606 55415 55658 55421
rect 55606 55357 55658 55363
rect 55618 55051 55646 55357
rect 55606 55045 55658 55051
rect 55606 54987 55658 54993
rect 53974 54823 54026 54829
rect 53974 54765 54026 54771
rect 53878 54749 53930 54755
rect 53878 54691 53930 54697
rect 53398 51567 53450 51573
rect 53398 51509 53450 51515
rect 53206 51419 53258 51425
rect 53206 51361 53258 51367
rect 53110 37211 53162 37217
rect 53110 37153 53162 37159
rect 52822 31883 52874 31889
rect 52822 31825 52874 31831
rect 52630 15159 52682 15165
rect 52630 15101 52682 15107
rect 52642 7765 52670 15101
rect 52918 10349 52970 10355
rect 52918 10291 52970 10297
rect 52930 8579 52958 10291
rect 53122 9097 53150 37153
rect 53110 9091 53162 9097
rect 53110 9033 53162 9039
rect 52918 8573 52970 8579
rect 52918 8515 52970 8521
rect 53110 8351 53162 8357
rect 53110 8293 53162 8299
rect 52630 7759 52682 7765
rect 52630 7701 52682 7707
rect 52726 7759 52778 7765
rect 52726 7701 52778 7707
rect 52438 7093 52490 7099
rect 52438 7035 52490 7041
rect 52534 5687 52586 5693
rect 52534 5629 52586 5635
rect 52546 800 52574 5629
rect 52630 4355 52682 4361
rect 52630 4297 52682 4303
rect 52642 800 52670 4297
rect 52738 800 52766 7701
rect 52918 7611 52970 7617
rect 52918 7553 52970 7559
rect 52822 6945 52874 6951
rect 52822 6887 52874 6893
rect 52834 3547 52862 6887
rect 52822 3541 52874 3547
rect 52822 3483 52874 3489
rect 52930 3344 52958 7553
rect 53014 4281 53066 4287
rect 53014 4223 53066 4229
rect 52834 3316 52958 3344
rect 52834 2511 52862 3316
rect 52918 2949 52970 2955
rect 52918 2891 52970 2897
rect 52822 2505 52874 2511
rect 52822 2447 52874 2453
rect 52930 800 52958 2891
rect 53026 800 53054 4223
rect 53122 800 53150 8293
rect 53218 7691 53246 51361
rect 53782 37433 53834 37439
rect 53782 37375 53834 37381
rect 53794 37143 53822 37375
rect 53782 37137 53834 37143
rect 53782 37079 53834 37085
rect 53890 28337 53918 54691
rect 53878 28331 53930 28337
rect 53878 28273 53930 28279
rect 53986 15239 54014 54765
rect 55030 50753 55082 50759
rect 55030 50695 55082 50701
rect 54454 50087 54506 50093
rect 54454 50029 54506 50035
rect 54262 26259 54314 26265
rect 54262 26201 54314 26207
rect 53974 15233 54026 15239
rect 53974 15175 54026 15181
rect 54274 12224 54302 26201
rect 54466 16793 54494 50029
rect 54742 36101 54794 36107
rect 54742 36043 54794 36049
rect 54754 29521 54782 36043
rect 54742 29515 54794 29521
rect 54742 29457 54794 29463
rect 54934 22337 54986 22343
rect 54934 22279 54986 22285
rect 54646 16935 54698 16941
rect 54646 16877 54698 16883
rect 54454 16787 54506 16793
rect 54454 16729 54506 16735
rect 54658 13759 54686 16877
rect 54646 13753 54698 13759
rect 54646 13695 54698 13701
rect 54274 12196 54494 12224
rect 54358 10793 54410 10799
rect 54358 10735 54410 10741
rect 54166 9831 54218 9837
rect 54166 9773 54218 9779
rect 54178 9245 54206 9773
rect 54262 9609 54314 9615
rect 54262 9551 54314 9557
rect 54166 9239 54218 9245
rect 54166 9181 54218 9187
rect 53878 9091 53930 9097
rect 53878 9033 53930 9039
rect 53494 8277 53546 8283
rect 53494 8219 53546 8225
rect 53206 7685 53258 7691
rect 53206 7627 53258 7633
rect 53302 5021 53354 5027
rect 53302 4963 53354 4969
rect 53314 2900 53342 4963
rect 53398 3689 53450 3695
rect 53398 3631 53450 3637
rect 53218 2872 53342 2900
rect 53218 800 53246 2872
rect 53410 800 53438 3631
rect 53506 800 53534 8219
rect 53686 5687 53738 5693
rect 53686 5629 53738 5635
rect 53590 5613 53642 5619
rect 53590 5555 53642 5561
rect 53602 800 53630 5555
rect 53698 2955 53726 5629
rect 53782 3023 53834 3029
rect 53782 2965 53834 2971
rect 53686 2949 53738 2955
rect 53686 2891 53738 2897
rect 53794 1568 53822 2965
rect 53698 1540 53822 1568
rect 53698 800 53726 1540
rect 53890 800 53918 9033
rect 54178 8949 54206 9181
rect 54166 8943 54218 8949
rect 54166 8885 54218 8891
rect 53974 6353 54026 6359
rect 53974 6295 54026 6301
rect 53986 800 54014 6295
rect 54070 4355 54122 4361
rect 54070 4297 54122 4303
rect 54082 800 54110 4297
rect 54274 800 54302 9551
rect 54370 8431 54398 10735
rect 54358 8425 54410 8431
rect 54358 8367 54410 8373
rect 54466 7214 54494 12196
rect 54838 9609 54890 9615
rect 54838 9551 54890 9557
rect 54550 8795 54602 8801
rect 54550 8737 54602 8743
rect 54370 7186 54494 7214
rect 54370 7099 54398 7186
rect 54358 7093 54410 7099
rect 54358 7035 54410 7041
rect 54358 3615 54410 3621
rect 54358 3557 54410 3563
rect 54370 1864 54398 3557
rect 54454 2801 54506 2807
rect 54454 2743 54506 2749
rect 54466 2585 54494 2743
rect 54454 2579 54506 2585
rect 54454 2521 54506 2527
rect 54370 1836 54494 1864
rect 54358 1765 54410 1771
rect 54358 1707 54410 1713
rect 54370 800 54398 1707
rect 54466 800 54494 1836
rect 54562 800 54590 8737
rect 54742 7019 54794 7025
rect 54742 6961 54794 6967
rect 54646 6353 54698 6359
rect 54646 6295 54698 6301
rect 54658 1771 54686 6295
rect 54646 1765 54698 1771
rect 54646 1707 54698 1713
rect 54754 800 54782 6961
rect 54850 4287 54878 9551
rect 54946 5915 54974 22279
rect 55042 10429 55070 50695
rect 55714 50315 55742 56689
rect 56002 56531 56030 59200
rect 55990 56525 56042 56531
rect 55990 56467 56042 56473
rect 56482 55717 56510 59200
rect 57058 57049 57086 59200
rect 57046 57043 57098 57049
rect 57046 56985 57098 56991
rect 56950 56747 57002 56753
rect 56950 56689 57002 56695
rect 56470 55711 56522 55717
rect 56470 55653 56522 55659
rect 55894 55563 55946 55569
rect 55894 55505 55946 55511
rect 55702 50309 55754 50315
rect 55702 50251 55754 50257
rect 55906 49205 55934 55505
rect 56962 49723 56990 56689
rect 57538 55717 57566 59200
rect 57526 55711 57578 55717
rect 57526 55653 57578 55659
rect 57334 55415 57386 55421
rect 57334 55357 57386 55363
rect 56950 49717 57002 49723
rect 56950 49659 57002 49665
rect 55894 49199 55946 49205
rect 55894 49141 55946 49147
rect 56278 48977 56330 48983
rect 56278 48919 56330 48925
rect 55318 44093 55370 44099
rect 55318 44035 55370 44041
rect 55330 11687 55358 44035
rect 55894 43871 55946 43877
rect 55894 43813 55946 43819
rect 55318 11681 55370 11687
rect 55318 11623 55370 11629
rect 55030 10423 55082 10429
rect 55030 10365 55082 10371
rect 55702 10127 55754 10133
rect 55702 10069 55754 10075
rect 55030 9535 55082 9541
rect 55030 9477 55082 9483
rect 55318 9535 55370 9541
rect 55318 9477 55370 9483
rect 54934 5909 54986 5915
rect 54934 5851 54986 5857
rect 54838 4281 54890 4287
rect 54838 4223 54890 4229
rect 55042 3640 55070 9477
rect 55126 6279 55178 6285
rect 55126 6221 55178 6227
rect 54946 3612 55070 3640
rect 54838 2949 54890 2955
rect 54838 2891 54890 2897
rect 54850 800 54878 2891
rect 54946 800 54974 3612
rect 55138 3196 55166 6221
rect 55222 3541 55274 3547
rect 55222 3483 55274 3489
rect 55042 3168 55166 3196
rect 55042 800 55070 3168
rect 55234 800 55262 3483
rect 55330 800 55358 9477
rect 55414 7019 55466 7025
rect 55414 6961 55466 6967
rect 55426 800 55454 6961
rect 55606 4355 55658 4361
rect 55606 4297 55658 4303
rect 55618 800 55646 4297
rect 55714 800 55742 10069
rect 55906 9763 55934 43813
rect 55990 28109 56042 28115
rect 55990 28051 56042 28057
rect 56002 10429 56030 28051
rect 56182 12347 56234 12353
rect 56182 12289 56234 12295
rect 56194 11909 56222 12289
rect 56182 11903 56234 11909
rect 56182 11845 56234 11851
rect 56290 10577 56318 48919
rect 57142 43575 57194 43581
rect 57142 43517 57194 43523
rect 57154 12575 57182 43517
rect 57238 41429 57290 41435
rect 57238 41371 57290 41377
rect 57250 33887 57278 41371
rect 57238 33881 57290 33887
rect 57238 33823 57290 33829
rect 57346 23083 57374 55357
rect 57910 54897 57962 54903
rect 57910 54839 57962 54845
rect 57814 54231 57866 54237
rect 57814 54173 57866 54179
rect 57826 43063 57854 54173
rect 57814 43057 57866 43063
rect 57814 42999 57866 43005
rect 57922 33221 57950 54839
rect 58114 54385 58142 59200
rect 58594 56309 58622 59200
rect 58582 56303 58634 56309
rect 58582 56245 58634 56251
rect 58198 56229 58250 56235
rect 58198 56171 58250 56177
rect 58102 54379 58154 54385
rect 58102 54321 58154 54327
rect 57910 33215 57962 33221
rect 57910 33157 57962 33163
rect 57430 31735 57482 31741
rect 57430 31677 57482 31683
rect 57334 23077 57386 23083
rect 57334 23019 57386 23025
rect 57142 12569 57194 12575
rect 57142 12511 57194 12517
rect 56854 11607 56906 11613
rect 56854 11549 56906 11555
rect 56374 10941 56426 10947
rect 56374 10883 56426 10889
rect 56278 10571 56330 10577
rect 56278 10513 56330 10519
rect 55990 10423 56042 10429
rect 55990 10365 56042 10371
rect 56086 10127 56138 10133
rect 56086 10069 56138 10075
rect 55894 9757 55946 9763
rect 55894 9699 55946 9705
rect 55990 9165 56042 9171
rect 55990 9107 56042 9113
rect 55798 7685 55850 7691
rect 55798 7627 55850 7633
rect 55810 800 55838 7627
rect 56002 3917 56030 9107
rect 55990 3911 56042 3917
rect 55990 3853 56042 3859
rect 55894 3763 55946 3769
rect 55894 3705 55946 3711
rect 55906 800 55934 3705
rect 56098 800 56126 10069
rect 56386 9116 56414 10883
rect 56758 10127 56810 10133
rect 56758 10069 56810 10075
rect 56770 9116 56798 10069
rect 56290 9088 56414 9116
rect 56482 9088 56798 9116
rect 56182 7685 56234 7691
rect 56182 7627 56234 7633
rect 56194 800 56222 7627
rect 56290 7044 56318 9088
rect 56374 8943 56426 8949
rect 56374 8885 56426 8891
rect 56386 7173 56414 8885
rect 56374 7167 56426 7173
rect 56374 7109 56426 7115
rect 56290 7016 56414 7044
rect 56278 6945 56330 6951
rect 56278 6887 56330 6893
rect 56290 5841 56318 6887
rect 56278 5835 56330 5841
rect 56278 5777 56330 5783
rect 56278 3615 56330 3621
rect 56278 3557 56330 3563
rect 56290 800 56318 3557
rect 56386 3547 56414 7016
rect 56374 3541 56426 3547
rect 56374 3483 56426 3489
rect 56482 800 56510 9088
rect 56566 9017 56618 9023
rect 56566 8959 56618 8965
rect 56578 4139 56606 8959
rect 56866 8949 56894 11549
rect 57142 10867 57194 10873
rect 57142 10809 57194 10815
rect 56854 8943 56906 8949
rect 56854 8885 56906 8891
rect 56950 8351 57002 8357
rect 56950 8293 57002 8299
rect 56758 7167 56810 7173
rect 56758 7109 56810 7115
rect 56662 4355 56714 4361
rect 56662 4297 56714 4303
rect 56566 4133 56618 4139
rect 56566 4075 56618 4081
rect 56566 3467 56618 3473
rect 56566 3409 56618 3415
rect 56578 800 56606 3409
rect 56674 800 56702 4297
rect 56770 3843 56798 7109
rect 56854 6427 56906 6433
rect 56854 6369 56906 6375
rect 56758 3837 56810 3843
rect 56758 3779 56810 3785
rect 56758 3541 56810 3547
rect 56758 3483 56810 3489
rect 56770 800 56798 3483
rect 56866 3251 56894 6369
rect 56854 3245 56906 3251
rect 56854 3187 56906 3193
rect 56962 800 56990 8293
rect 57046 5021 57098 5027
rect 57046 4963 57098 4969
rect 57058 800 57086 4963
rect 57154 4213 57182 10809
rect 57442 10429 57470 31677
rect 58006 28109 58058 28115
rect 58006 28051 58058 28057
rect 58018 27893 58046 28051
rect 58006 27887 58058 27893
rect 58006 27829 58058 27835
rect 58210 13241 58238 56171
rect 59170 55199 59198 59200
rect 59158 55193 59210 55199
rect 59158 55135 59210 55141
rect 59650 53867 59678 59200
rect 59638 53861 59690 53867
rect 59638 53803 59690 53809
rect 58198 13235 58250 13241
rect 58198 13177 58250 13183
rect 57526 12199 57578 12205
rect 57526 12141 57578 12147
rect 57430 10423 57482 10429
rect 57430 10365 57482 10371
rect 57238 9017 57290 9023
rect 57238 8959 57290 8965
rect 57142 4207 57194 4213
rect 57142 4149 57194 4155
rect 57142 3837 57194 3843
rect 57142 3779 57194 3785
rect 57154 800 57182 3779
rect 57250 800 57278 8959
rect 57334 7685 57386 7691
rect 57334 7627 57386 7633
rect 57346 3473 57374 7627
rect 57430 5687 57482 5693
rect 57430 5629 57482 5635
rect 57334 3467 57386 3473
rect 57334 3409 57386 3415
rect 57442 800 57470 5629
rect 57538 800 57566 12141
rect 58198 11829 58250 11835
rect 58198 11771 58250 11777
rect 57622 9683 57674 9689
rect 57622 9625 57674 9631
rect 57634 800 57662 9625
rect 58102 6353 58154 6359
rect 58102 6295 58154 6301
rect 57718 5835 57770 5841
rect 57718 5777 57770 5783
rect 57730 2955 57758 5777
rect 57814 5095 57866 5101
rect 57814 5037 57866 5043
rect 57718 2949 57770 2955
rect 57718 2891 57770 2897
rect 57826 800 57854 5037
rect 57910 3837 57962 3843
rect 57910 3779 57962 3785
rect 57922 800 57950 3779
rect 58006 3245 58058 3251
rect 58006 3187 58058 3193
rect 58018 800 58046 3187
rect 58114 800 58142 6295
rect 58210 3695 58238 11771
rect 58582 10201 58634 10207
rect 58582 10143 58634 10149
rect 58390 8277 58442 8283
rect 58390 8219 58442 8225
rect 58294 4281 58346 4287
rect 58294 4223 58346 4229
rect 58198 3689 58250 3695
rect 58198 3631 58250 3637
rect 58306 800 58334 4223
rect 58402 800 58430 8219
rect 58486 7019 58538 7025
rect 58486 6961 58538 6967
rect 58498 800 58526 6961
rect 58594 800 58622 10143
rect 59830 8203 59882 8209
rect 59830 8145 59882 8151
rect 58966 8129 59018 8135
rect 58966 8071 59018 8077
rect 58774 7611 58826 7617
rect 58774 7553 58826 7559
rect 58786 800 58814 7553
rect 58870 6279 58922 6285
rect 58870 6221 58922 6227
rect 58882 800 58910 6221
rect 58978 800 59006 8071
rect 59350 7537 59402 7543
rect 59350 7479 59402 7485
rect 59254 5169 59306 5175
rect 59254 5111 59306 5117
rect 59158 4133 59210 4139
rect 59158 4075 59210 4081
rect 59170 800 59198 4075
rect 59266 800 59294 5111
rect 59362 800 59390 7479
rect 59638 5613 59690 5619
rect 59638 5555 59690 5561
rect 59446 2949 59498 2955
rect 59446 2891 59498 2897
rect 59458 800 59486 2891
rect 59650 800 59678 5555
rect 59734 3689 59786 3695
rect 59734 3631 59786 3637
rect 59746 800 59774 3631
rect 59842 800 59870 8145
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< via2 >>
rect 4268 57302 4324 57304
rect 4348 57302 4404 57304
rect 4428 57302 4484 57304
rect 4508 57302 4564 57304
rect 4268 57250 4294 57302
rect 4294 57250 4324 57302
rect 4348 57250 4358 57302
rect 4358 57250 4404 57302
rect 4428 57250 4474 57302
rect 4474 57250 4484 57302
rect 4508 57250 4538 57302
rect 4538 57250 4564 57302
rect 4268 57248 4324 57250
rect 4348 57248 4404 57250
rect 4428 57248 4484 57250
rect 4508 57248 4564 57250
rect 4268 55970 4324 55972
rect 4348 55970 4404 55972
rect 4428 55970 4484 55972
rect 4508 55970 4564 55972
rect 4268 55918 4294 55970
rect 4294 55918 4324 55970
rect 4348 55918 4358 55970
rect 4358 55918 4404 55970
rect 4428 55918 4474 55970
rect 4474 55918 4484 55970
rect 4508 55918 4538 55970
rect 4538 55918 4564 55970
rect 4268 55916 4324 55918
rect 4348 55916 4404 55918
rect 4428 55916 4484 55918
rect 4508 55916 4564 55918
rect 4268 54638 4324 54640
rect 4348 54638 4404 54640
rect 4428 54638 4484 54640
rect 4508 54638 4564 54640
rect 4268 54586 4294 54638
rect 4294 54586 4324 54638
rect 4348 54586 4358 54638
rect 4358 54586 4404 54638
rect 4428 54586 4474 54638
rect 4474 54586 4484 54638
rect 4508 54586 4538 54638
rect 4538 54586 4564 54638
rect 4268 54584 4324 54586
rect 4348 54584 4404 54586
rect 4428 54584 4484 54586
rect 4508 54584 4564 54586
rect 4268 53306 4324 53308
rect 4348 53306 4404 53308
rect 4428 53306 4484 53308
rect 4508 53306 4564 53308
rect 4268 53254 4294 53306
rect 4294 53254 4324 53306
rect 4348 53254 4358 53306
rect 4358 53254 4404 53306
rect 4428 53254 4474 53306
rect 4474 53254 4484 53306
rect 4508 53254 4538 53306
rect 4538 53254 4564 53306
rect 4268 53252 4324 53254
rect 4348 53252 4404 53254
rect 4428 53252 4484 53254
rect 4508 53252 4564 53254
rect 4268 51974 4324 51976
rect 4348 51974 4404 51976
rect 4428 51974 4484 51976
rect 4508 51974 4564 51976
rect 4268 51922 4294 51974
rect 4294 51922 4324 51974
rect 4348 51922 4358 51974
rect 4358 51922 4404 51974
rect 4428 51922 4474 51974
rect 4474 51922 4484 51974
rect 4508 51922 4538 51974
rect 4538 51922 4564 51974
rect 4268 51920 4324 51922
rect 4348 51920 4404 51922
rect 4428 51920 4484 51922
rect 4508 51920 4564 51922
rect 4268 50642 4324 50644
rect 4348 50642 4404 50644
rect 4428 50642 4484 50644
rect 4508 50642 4564 50644
rect 4268 50590 4294 50642
rect 4294 50590 4324 50642
rect 4348 50590 4358 50642
rect 4358 50590 4404 50642
rect 4428 50590 4474 50642
rect 4474 50590 4484 50642
rect 4508 50590 4538 50642
rect 4538 50590 4564 50642
rect 4268 50588 4324 50590
rect 4348 50588 4404 50590
rect 4428 50588 4484 50590
rect 4508 50588 4564 50590
rect 4268 49310 4324 49312
rect 4348 49310 4404 49312
rect 4428 49310 4484 49312
rect 4508 49310 4564 49312
rect 4268 49258 4294 49310
rect 4294 49258 4324 49310
rect 4348 49258 4358 49310
rect 4358 49258 4404 49310
rect 4428 49258 4474 49310
rect 4474 49258 4484 49310
rect 4508 49258 4538 49310
rect 4538 49258 4564 49310
rect 4268 49256 4324 49258
rect 4348 49256 4404 49258
rect 4428 49256 4484 49258
rect 4508 49256 4564 49258
rect 4268 47978 4324 47980
rect 4348 47978 4404 47980
rect 4428 47978 4484 47980
rect 4508 47978 4564 47980
rect 4268 47926 4294 47978
rect 4294 47926 4324 47978
rect 4348 47926 4358 47978
rect 4358 47926 4404 47978
rect 4428 47926 4474 47978
rect 4474 47926 4484 47978
rect 4508 47926 4538 47978
rect 4538 47926 4564 47978
rect 4268 47924 4324 47926
rect 4348 47924 4404 47926
rect 4428 47924 4484 47926
rect 4508 47924 4564 47926
rect 4268 46646 4324 46648
rect 4348 46646 4404 46648
rect 4428 46646 4484 46648
rect 4508 46646 4564 46648
rect 4268 46594 4294 46646
rect 4294 46594 4324 46646
rect 4348 46594 4358 46646
rect 4358 46594 4404 46646
rect 4428 46594 4474 46646
rect 4474 46594 4484 46646
rect 4508 46594 4538 46646
rect 4538 46594 4564 46646
rect 4268 46592 4324 46594
rect 4348 46592 4404 46594
rect 4428 46592 4484 46594
rect 4508 46592 4564 46594
rect 4268 45314 4324 45316
rect 4348 45314 4404 45316
rect 4428 45314 4484 45316
rect 4508 45314 4564 45316
rect 4268 45262 4294 45314
rect 4294 45262 4324 45314
rect 4348 45262 4358 45314
rect 4358 45262 4404 45314
rect 4428 45262 4474 45314
rect 4474 45262 4484 45314
rect 4508 45262 4538 45314
rect 4538 45262 4564 45314
rect 4268 45260 4324 45262
rect 4348 45260 4404 45262
rect 4428 45260 4484 45262
rect 4508 45260 4564 45262
rect 4268 43982 4324 43984
rect 4348 43982 4404 43984
rect 4428 43982 4484 43984
rect 4508 43982 4564 43984
rect 4268 43930 4294 43982
rect 4294 43930 4324 43982
rect 4348 43930 4358 43982
rect 4358 43930 4404 43982
rect 4428 43930 4474 43982
rect 4474 43930 4484 43982
rect 4508 43930 4538 43982
rect 4538 43930 4564 43982
rect 4268 43928 4324 43930
rect 4348 43928 4404 43930
rect 4428 43928 4484 43930
rect 4508 43928 4564 43930
rect 4268 42650 4324 42652
rect 4348 42650 4404 42652
rect 4428 42650 4484 42652
rect 4508 42650 4564 42652
rect 4268 42598 4294 42650
rect 4294 42598 4324 42650
rect 4348 42598 4358 42650
rect 4358 42598 4404 42650
rect 4428 42598 4474 42650
rect 4474 42598 4484 42650
rect 4508 42598 4538 42650
rect 4538 42598 4564 42650
rect 4268 42596 4324 42598
rect 4348 42596 4404 42598
rect 4428 42596 4484 42598
rect 4508 42596 4564 42598
rect 4268 41318 4324 41320
rect 4348 41318 4404 41320
rect 4428 41318 4484 41320
rect 4508 41318 4564 41320
rect 4268 41266 4294 41318
rect 4294 41266 4324 41318
rect 4348 41266 4358 41318
rect 4358 41266 4404 41318
rect 4428 41266 4474 41318
rect 4474 41266 4484 41318
rect 4508 41266 4538 41318
rect 4538 41266 4564 41318
rect 4268 41264 4324 41266
rect 4348 41264 4404 41266
rect 4428 41264 4484 41266
rect 4508 41264 4564 41266
rect 4268 39986 4324 39988
rect 4348 39986 4404 39988
rect 4428 39986 4484 39988
rect 4508 39986 4564 39988
rect 4268 39934 4294 39986
rect 4294 39934 4324 39986
rect 4348 39934 4358 39986
rect 4358 39934 4404 39986
rect 4428 39934 4474 39986
rect 4474 39934 4484 39986
rect 4508 39934 4538 39986
rect 4538 39934 4564 39986
rect 4268 39932 4324 39934
rect 4348 39932 4404 39934
rect 4428 39932 4484 39934
rect 4508 39932 4564 39934
rect 4268 38654 4324 38656
rect 4348 38654 4404 38656
rect 4428 38654 4484 38656
rect 4508 38654 4564 38656
rect 4268 38602 4294 38654
rect 4294 38602 4324 38654
rect 4348 38602 4358 38654
rect 4358 38602 4404 38654
rect 4428 38602 4474 38654
rect 4474 38602 4484 38654
rect 4508 38602 4538 38654
rect 4538 38602 4564 38654
rect 4268 38600 4324 38602
rect 4348 38600 4404 38602
rect 4428 38600 4484 38602
rect 4508 38600 4564 38602
rect 4268 37322 4324 37324
rect 4348 37322 4404 37324
rect 4428 37322 4484 37324
rect 4508 37322 4564 37324
rect 4268 37270 4294 37322
rect 4294 37270 4324 37322
rect 4348 37270 4358 37322
rect 4358 37270 4404 37322
rect 4428 37270 4474 37322
rect 4474 37270 4484 37322
rect 4508 37270 4538 37322
rect 4538 37270 4564 37322
rect 4268 37268 4324 37270
rect 4348 37268 4404 37270
rect 4428 37268 4484 37270
rect 4508 37268 4564 37270
rect 4268 35990 4324 35992
rect 4348 35990 4404 35992
rect 4428 35990 4484 35992
rect 4508 35990 4564 35992
rect 4268 35938 4294 35990
rect 4294 35938 4324 35990
rect 4348 35938 4358 35990
rect 4358 35938 4404 35990
rect 4428 35938 4474 35990
rect 4474 35938 4484 35990
rect 4508 35938 4538 35990
rect 4538 35938 4564 35990
rect 4268 35936 4324 35938
rect 4348 35936 4404 35938
rect 4428 35936 4484 35938
rect 4508 35936 4564 35938
rect 4268 34658 4324 34660
rect 4348 34658 4404 34660
rect 4428 34658 4484 34660
rect 4508 34658 4564 34660
rect 4268 34606 4294 34658
rect 4294 34606 4324 34658
rect 4348 34606 4358 34658
rect 4358 34606 4404 34658
rect 4428 34606 4474 34658
rect 4474 34606 4484 34658
rect 4508 34606 4538 34658
rect 4538 34606 4564 34658
rect 4268 34604 4324 34606
rect 4348 34604 4404 34606
rect 4428 34604 4484 34606
rect 4508 34604 4564 34606
rect 4268 33326 4324 33328
rect 4348 33326 4404 33328
rect 4428 33326 4484 33328
rect 4508 33326 4564 33328
rect 4268 33274 4294 33326
rect 4294 33274 4324 33326
rect 4348 33274 4358 33326
rect 4358 33274 4404 33326
rect 4428 33274 4474 33326
rect 4474 33274 4484 33326
rect 4508 33274 4538 33326
rect 4538 33274 4564 33326
rect 4268 33272 4324 33274
rect 4348 33272 4404 33274
rect 4428 33272 4484 33274
rect 4508 33272 4564 33274
rect 4268 31994 4324 31996
rect 4348 31994 4404 31996
rect 4428 31994 4484 31996
rect 4508 31994 4564 31996
rect 4268 31942 4294 31994
rect 4294 31942 4324 31994
rect 4348 31942 4358 31994
rect 4358 31942 4404 31994
rect 4428 31942 4474 31994
rect 4474 31942 4484 31994
rect 4508 31942 4538 31994
rect 4538 31942 4564 31994
rect 4268 31940 4324 31942
rect 4348 31940 4404 31942
rect 4428 31940 4484 31942
rect 4508 31940 4564 31942
rect 4268 30662 4324 30664
rect 4348 30662 4404 30664
rect 4428 30662 4484 30664
rect 4508 30662 4564 30664
rect 4268 30610 4294 30662
rect 4294 30610 4324 30662
rect 4348 30610 4358 30662
rect 4358 30610 4404 30662
rect 4428 30610 4474 30662
rect 4474 30610 4484 30662
rect 4508 30610 4538 30662
rect 4538 30610 4564 30662
rect 4268 30608 4324 30610
rect 4348 30608 4404 30610
rect 4428 30608 4484 30610
rect 4508 30608 4564 30610
rect 4268 29330 4324 29332
rect 4348 29330 4404 29332
rect 4428 29330 4484 29332
rect 4508 29330 4564 29332
rect 4268 29278 4294 29330
rect 4294 29278 4324 29330
rect 4348 29278 4358 29330
rect 4358 29278 4404 29330
rect 4428 29278 4474 29330
rect 4474 29278 4484 29330
rect 4508 29278 4538 29330
rect 4538 29278 4564 29330
rect 4268 29276 4324 29278
rect 4348 29276 4404 29278
rect 4428 29276 4484 29278
rect 4508 29276 4564 29278
rect 4268 27998 4324 28000
rect 4348 27998 4404 28000
rect 4428 27998 4484 28000
rect 4508 27998 4564 28000
rect 4268 27946 4294 27998
rect 4294 27946 4324 27998
rect 4348 27946 4358 27998
rect 4358 27946 4404 27998
rect 4428 27946 4474 27998
rect 4474 27946 4484 27998
rect 4508 27946 4538 27998
rect 4538 27946 4564 27998
rect 4268 27944 4324 27946
rect 4348 27944 4404 27946
rect 4428 27944 4484 27946
rect 4508 27944 4564 27946
rect 4268 26666 4324 26668
rect 4348 26666 4404 26668
rect 4428 26666 4484 26668
rect 4508 26666 4564 26668
rect 4268 26614 4294 26666
rect 4294 26614 4324 26666
rect 4348 26614 4358 26666
rect 4358 26614 4404 26666
rect 4428 26614 4474 26666
rect 4474 26614 4484 26666
rect 4508 26614 4538 26666
rect 4538 26614 4564 26666
rect 4268 26612 4324 26614
rect 4348 26612 4404 26614
rect 4428 26612 4484 26614
rect 4508 26612 4564 26614
rect 4268 25334 4324 25336
rect 4348 25334 4404 25336
rect 4428 25334 4484 25336
rect 4508 25334 4564 25336
rect 4268 25282 4294 25334
rect 4294 25282 4324 25334
rect 4348 25282 4358 25334
rect 4358 25282 4404 25334
rect 4428 25282 4474 25334
rect 4474 25282 4484 25334
rect 4508 25282 4538 25334
rect 4538 25282 4564 25334
rect 4268 25280 4324 25282
rect 4348 25280 4404 25282
rect 4428 25280 4484 25282
rect 4508 25280 4564 25282
rect 4268 24002 4324 24004
rect 4348 24002 4404 24004
rect 4428 24002 4484 24004
rect 4508 24002 4564 24004
rect 4268 23950 4294 24002
rect 4294 23950 4324 24002
rect 4348 23950 4358 24002
rect 4358 23950 4404 24002
rect 4428 23950 4474 24002
rect 4474 23950 4484 24002
rect 4508 23950 4538 24002
rect 4538 23950 4564 24002
rect 4268 23948 4324 23950
rect 4348 23948 4404 23950
rect 4428 23948 4484 23950
rect 4508 23948 4564 23950
rect 4268 22670 4324 22672
rect 4348 22670 4404 22672
rect 4428 22670 4484 22672
rect 4508 22670 4564 22672
rect 4268 22618 4294 22670
rect 4294 22618 4324 22670
rect 4348 22618 4358 22670
rect 4358 22618 4404 22670
rect 4428 22618 4474 22670
rect 4474 22618 4484 22670
rect 4508 22618 4538 22670
rect 4538 22618 4564 22670
rect 4268 22616 4324 22618
rect 4348 22616 4404 22618
rect 4428 22616 4484 22618
rect 4508 22616 4564 22618
rect 4268 21338 4324 21340
rect 4348 21338 4404 21340
rect 4428 21338 4484 21340
rect 4508 21338 4564 21340
rect 4268 21286 4294 21338
rect 4294 21286 4324 21338
rect 4348 21286 4358 21338
rect 4358 21286 4404 21338
rect 4428 21286 4474 21338
rect 4474 21286 4484 21338
rect 4508 21286 4538 21338
rect 4538 21286 4564 21338
rect 4268 21284 4324 21286
rect 4348 21284 4404 21286
rect 4428 21284 4484 21286
rect 4508 21284 4564 21286
rect 4268 20006 4324 20008
rect 4348 20006 4404 20008
rect 4428 20006 4484 20008
rect 4508 20006 4564 20008
rect 4268 19954 4294 20006
rect 4294 19954 4324 20006
rect 4348 19954 4358 20006
rect 4358 19954 4404 20006
rect 4428 19954 4474 20006
rect 4474 19954 4484 20006
rect 4508 19954 4538 20006
rect 4538 19954 4564 20006
rect 4268 19952 4324 19954
rect 4348 19952 4404 19954
rect 4428 19952 4484 19954
rect 4508 19952 4564 19954
rect 4268 18674 4324 18676
rect 4348 18674 4404 18676
rect 4428 18674 4484 18676
rect 4508 18674 4564 18676
rect 4268 18622 4294 18674
rect 4294 18622 4324 18674
rect 4348 18622 4358 18674
rect 4358 18622 4404 18674
rect 4428 18622 4474 18674
rect 4474 18622 4484 18674
rect 4508 18622 4538 18674
rect 4538 18622 4564 18674
rect 4268 18620 4324 18622
rect 4348 18620 4404 18622
rect 4428 18620 4484 18622
rect 4508 18620 4564 18622
rect 4268 17342 4324 17344
rect 4348 17342 4404 17344
rect 4428 17342 4484 17344
rect 4508 17342 4564 17344
rect 4268 17290 4294 17342
rect 4294 17290 4324 17342
rect 4348 17290 4358 17342
rect 4358 17290 4404 17342
rect 4428 17290 4474 17342
rect 4474 17290 4484 17342
rect 4508 17290 4538 17342
rect 4538 17290 4564 17342
rect 4268 17288 4324 17290
rect 4348 17288 4404 17290
rect 4428 17288 4484 17290
rect 4508 17288 4564 17290
rect 4268 16010 4324 16012
rect 4348 16010 4404 16012
rect 4428 16010 4484 16012
rect 4508 16010 4564 16012
rect 4268 15958 4294 16010
rect 4294 15958 4324 16010
rect 4348 15958 4358 16010
rect 4358 15958 4404 16010
rect 4428 15958 4474 16010
rect 4474 15958 4484 16010
rect 4508 15958 4538 16010
rect 4538 15958 4564 16010
rect 4268 15956 4324 15958
rect 4348 15956 4404 15958
rect 4428 15956 4484 15958
rect 4508 15956 4564 15958
rect 4268 14678 4324 14680
rect 4348 14678 4404 14680
rect 4428 14678 4484 14680
rect 4508 14678 4564 14680
rect 4268 14626 4294 14678
rect 4294 14626 4324 14678
rect 4348 14626 4358 14678
rect 4358 14626 4404 14678
rect 4428 14626 4474 14678
rect 4474 14626 4484 14678
rect 4508 14626 4538 14678
rect 4538 14626 4564 14678
rect 4268 14624 4324 14626
rect 4348 14624 4404 14626
rect 4428 14624 4484 14626
rect 4508 14624 4564 14626
rect 4268 13346 4324 13348
rect 4348 13346 4404 13348
rect 4428 13346 4484 13348
rect 4508 13346 4564 13348
rect 4268 13294 4294 13346
rect 4294 13294 4324 13346
rect 4348 13294 4358 13346
rect 4358 13294 4404 13346
rect 4428 13294 4474 13346
rect 4474 13294 4484 13346
rect 4508 13294 4538 13346
rect 4538 13294 4564 13346
rect 4268 13292 4324 13294
rect 4348 13292 4404 13294
rect 4428 13292 4484 13294
rect 4508 13292 4564 13294
rect 4268 12014 4324 12016
rect 4348 12014 4404 12016
rect 4428 12014 4484 12016
rect 4508 12014 4564 12016
rect 4268 11962 4294 12014
rect 4294 11962 4324 12014
rect 4348 11962 4358 12014
rect 4358 11962 4404 12014
rect 4428 11962 4474 12014
rect 4474 11962 4484 12014
rect 4508 11962 4538 12014
rect 4538 11962 4564 12014
rect 4268 11960 4324 11962
rect 4348 11960 4404 11962
rect 4428 11960 4484 11962
rect 4508 11960 4564 11962
rect 4268 10682 4324 10684
rect 4348 10682 4404 10684
rect 4428 10682 4484 10684
rect 4508 10682 4564 10684
rect 4268 10630 4294 10682
rect 4294 10630 4324 10682
rect 4348 10630 4358 10682
rect 4358 10630 4404 10682
rect 4428 10630 4474 10682
rect 4474 10630 4484 10682
rect 4508 10630 4538 10682
rect 4538 10630 4564 10682
rect 4268 10628 4324 10630
rect 4348 10628 4404 10630
rect 4428 10628 4484 10630
rect 4508 10628 4564 10630
rect 4268 9350 4324 9352
rect 4348 9350 4404 9352
rect 4428 9350 4484 9352
rect 4508 9350 4564 9352
rect 4268 9298 4294 9350
rect 4294 9298 4324 9350
rect 4348 9298 4358 9350
rect 4358 9298 4404 9350
rect 4428 9298 4474 9350
rect 4474 9298 4484 9350
rect 4508 9298 4538 9350
rect 4538 9298 4564 9350
rect 4268 9296 4324 9298
rect 4348 9296 4404 9298
rect 4428 9296 4484 9298
rect 4508 9296 4564 9298
rect 4268 8018 4324 8020
rect 4348 8018 4404 8020
rect 4428 8018 4484 8020
rect 4508 8018 4564 8020
rect 4268 7966 4294 8018
rect 4294 7966 4324 8018
rect 4348 7966 4358 8018
rect 4358 7966 4404 8018
rect 4428 7966 4474 8018
rect 4474 7966 4484 8018
rect 4508 7966 4538 8018
rect 4538 7966 4564 8018
rect 4268 7964 4324 7966
rect 4348 7964 4404 7966
rect 4428 7964 4484 7966
rect 4508 7964 4564 7966
rect 4268 6686 4324 6688
rect 4348 6686 4404 6688
rect 4428 6686 4484 6688
rect 4508 6686 4564 6688
rect 4268 6634 4294 6686
rect 4294 6634 4324 6686
rect 4348 6634 4358 6686
rect 4358 6634 4404 6686
rect 4428 6634 4474 6686
rect 4474 6634 4484 6686
rect 4508 6634 4538 6686
rect 4538 6634 4564 6686
rect 4268 6632 4324 6634
rect 4348 6632 4404 6634
rect 4428 6632 4484 6634
rect 4508 6632 4564 6634
rect 4268 5354 4324 5356
rect 4348 5354 4404 5356
rect 4428 5354 4484 5356
rect 4508 5354 4564 5356
rect 4268 5302 4294 5354
rect 4294 5302 4324 5354
rect 4348 5302 4358 5354
rect 4358 5302 4404 5354
rect 4428 5302 4474 5354
rect 4474 5302 4484 5354
rect 4508 5302 4538 5354
rect 4538 5302 4564 5354
rect 4268 5300 4324 5302
rect 4348 5300 4404 5302
rect 4428 5300 4484 5302
rect 4508 5300 4564 5302
rect 4268 4022 4324 4024
rect 4348 4022 4404 4024
rect 4428 4022 4484 4024
rect 4508 4022 4564 4024
rect 4268 3970 4294 4022
rect 4294 3970 4324 4022
rect 4348 3970 4358 4022
rect 4358 3970 4404 4022
rect 4428 3970 4474 4022
rect 4474 3970 4484 4022
rect 4508 3970 4538 4022
rect 4538 3970 4564 4022
rect 4268 3968 4324 3970
rect 4348 3968 4404 3970
rect 4428 3968 4484 3970
rect 4508 3968 4564 3970
rect 4268 2690 4324 2692
rect 4348 2690 4404 2692
rect 4428 2690 4484 2692
rect 4508 2690 4564 2692
rect 4268 2638 4294 2690
rect 4294 2638 4324 2690
rect 4348 2638 4358 2690
rect 4358 2638 4404 2690
rect 4428 2638 4474 2690
rect 4474 2638 4484 2690
rect 4508 2638 4538 2690
rect 4538 2638 4564 2690
rect 4268 2636 4324 2638
rect 4348 2636 4404 2638
rect 4428 2636 4484 2638
rect 4508 2636 4564 2638
rect 19628 56636 19684 56638
rect 19708 56636 19764 56638
rect 19788 56636 19844 56638
rect 19868 56636 19924 56638
rect 19628 56584 19654 56636
rect 19654 56584 19684 56636
rect 19708 56584 19718 56636
rect 19718 56584 19764 56636
rect 19788 56584 19834 56636
rect 19834 56584 19844 56636
rect 19868 56584 19898 56636
rect 19898 56584 19924 56636
rect 19628 56582 19684 56584
rect 19708 56582 19764 56584
rect 19788 56582 19844 56584
rect 19868 56582 19924 56584
rect 19628 55304 19684 55306
rect 19708 55304 19764 55306
rect 19788 55304 19844 55306
rect 19868 55304 19924 55306
rect 19628 55252 19654 55304
rect 19654 55252 19684 55304
rect 19708 55252 19718 55304
rect 19718 55252 19764 55304
rect 19788 55252 19834 55304
rect 19834 55252 19844 55304
rect 19868 55252 19898 55304
rect 19898 55252 19924 55304
rect 19628 55250 19684 55252
rect 19708 55250 19764 55252
rect 19788 55250 19844 55252
rect 19868 55250 19924 55252
rect 19628 53972 19684 53974
rect 19708 53972 19764 53974
rect 19788 53972 19844 53974
rect 19868 53972 19924 53974
rect 19628 53920 19654 53972
rect 19654 53920 19684 53972
rect 19708 53920 19718 53972
rect 19718 53920 19764 53972
rect 19788 53920 19834 53972
rect 19834 53920 19844 53972
rect 19868 53920 19898 53972
rect 19898 53920 19924 53972
rect 19628 53918 19684 53920
rect 19708 53918 19764 53920
rect 19788 53918 19844 53920
rect 19868 53918 19924 53920
rect 19628 52640 19684 52642
rect 19708 52640 19764 52642
rect 19788 52640 19844 52642
rect 19868 52640 19924 52642
rect 19628 52588 19654 52640
rect 19654 52588 19684 52640
rect 19708 52588 19718 52640
rect 19718 52588 19764 52640
rect 19788 52588 19834 52640
rect 19834 52588 19844 52640
rect 19868 52588 19898 52640
rect 19898 52588 19924 52640
rect 19628 52586 19684 52588
rect 19708 52586 19764 52588
rect 19788 52586 19844 52588
rect 19868 52586 19924 52588
rect 19628 51308 19684 51310
rect 19708 51308 19764 51310
rect 19788 51308 19844 51310
rect 19868 51308 19924 51310
rect 19628 51256 19654 51308
rect 19654 51256 19684 51308
rect 19708 51256 19718 51308
rect 19718 51256 19764 51308
rect 19788 51256 19834 51308
rect 19834 51256 19844 51308
rect 19868 51256 19898 51308
rect 19898 51256 19924 51308
rect 19628 51254 19684 51256
rect 19708 51254 19764 51256
rect 19788 51254 19844 51256
rect 19868 51254 19924 51256
rect 19628 49976 19684 49978
rect 19708 49976 19764 49978
rect 19788 49976 19844 49978
rect 19868 49976 19924 49978
rect 19628 49924 19654 49976
rect 19654 49924 19684 49976
rect 19708 49924 19718 49976
rect 19718 49924 19764 49976
rect 19788 49924 19834 49976
rect 19834 49924 19844 49976
rect 19868 49924 19898 49976
rect 19898 49924 19924 49976
rect 19628 49922 19684 49924
rect 19708 49922 19764 49924
rect 19788 49922 19844 49924
rect 19868 49922 19924 49924
rect 19628 48644 19684 48646
rect 19708 48644 19764 48646
rect 19788 48644 19844 48646
rect 19868 48644 19924 48646
rect 19628 48592 19654 48644
rect 19654 48592 19684 48644
rect 19708 48592 19718 48644
rect 19718 48592 19764 48644
rect 19788 48592 19834 48644
rect 19834 48592 19844 48644
rect 19868 48592 19898 48644
rect 19898 48592 19924 48644
rect 19628 48590 19684 48592
rect 19708 48590 19764 48592
rect 19788 48590 19844 48592
rect 19868 48590 19924 48592
rect 19628 47312 19684 47314
rect 19708 47312 19764 47314
rect 19788 47312 19844 47314
rect 19868 47312 19924 47314
rect 19628 47260 19654 47312
rect 19654 47260 19684 47312
rect 19708 47260 19718 47312
rect 19718 47260 19764 47312
rect 19788 47260 19834 47312
rect 19834 47260 19844 47312
rect 19868 47260 19898 47312
rect 19898 47260 19924 47312
rect 19628 47258 19684 47260
rect 19708 47258 19764 47260
rect 19788 47258 19844 47260
rect 19868 47258 19924 47260
rect 19628 45980 19684 45982
rect 19708 45980 19764 45982
rect 19788 45980 19844 45982
rect 19868 45980 19924 45982
rect 19628 45928 19654 45980
rect 19654 45928 19684 45980
rect 19708 45928 19718 45980
rect 19718 45928 19764 45980
rect 19788 45928 19834 45980
rect 19834 45928 19844 45980
rect 19868 45928 19898 45980
rect 19898 45928 19924 45980
rect 19628 45926 19684 45928
rect 19708 45926 19764 45928
rect 19788 45926 19844 45928
rect 19868 45926 19924 45928
rect 19628 44648 19684 44650
rect 19708 44648 19764 44650
rect 19788 44648 19844 44650
rect 19868 44648 19924 44650
rect 19628 44596 19654 44648
rect 19654 44596 19684 44648
rect 19708 44596 19718 44648
rect 19718 44596 19764 44648
rect 19788 44596 19834 44648
rect 19834 44596 19844 44648
rect 19868 44596 19898 44648
rect 19898 44596 19924 44648
rect 19628 44594 19684 44596
rect 19708 44594 19764 44596
rect 19788 44594 19844 44596
rect 19868 44594 19924 44596
rect 19628 43316 19684 43318
rect 19708 43316 19764 43318
rect 19788 43316 19844 43318
rect 19868 43316 19924 43318
rect 19628 43264 19654 43316
rect 19654 43264 19684 43316
rect 19708 43264 19718 43316
rect 19718 43264 19764 43316
rect 19788 43264 19834 43316
rect 19834 43264 19844 43316
rect 19868 43264 19898 43316
rect 19898 43264 19924 43316
rect 19628 43262 19684 43264
rect 19708 43262 19764 43264
rect 19788 43262 19844 43264
rect 19868 43262 19924 43264
rect 19628 41984 19684 41986
rect 19708 41984 19764 41986
rect 19788 41984 19844 41986
rect 19868 41984 19924 41986
rect 19628 41932 19654 41984
rect 19654 41932 19684 41984
rect 19708 41932 19718 41984
rect 19718 41932 19764 41984
rect 19788 41932 19834 41984
rect 19834 41932 19844 41984
rect 19868 41932 19898 41984
rect 19898 41932 19924 41984
rect 19628 41930 19684 41932
rect 19708 41930 19764 41932
rect 19788 41930 19844 41932
rect 19868 41930 19924 41932
rect 19628 40652 19684 40654
rect 19708 40652 19764 40654
rect 19788 40652 19844 40654
rect 19868 40652 19924 40654
rect 19628 40600 19654 40652
rect 19654 40600 19684 40652
rect 19708 40600 19718 40652
rect 19718 40600 19764 40652
rect 19788 40600 19834 40652
rect 19834 40600 19844 40652
rect 19868 40600 19898 40652
rect 19898 40600 19924 40652
rect 19628 40598 19684 40600
rect 19708 40598 19764 40600
rect 19788 40598 19844 40600
rect 19868 40598 19924 40600
rect 19628 39320 19684 39322
rect 19708 39320 19764 39322
rect 19788 39320 19844 39322
rect 19868 39320 19924 39322
rect 19628 39268 19654 39320
rect 19654 39268 19684 39320
rect 19708 39268 19718 39320
rect 19718 39268 19764 39320
rect 19788 39268 19834 39320
rect 19834 39268 19844 39320
rect 19868 39268 19898 39320
rect 19898 39268 19924 39320
rect 19628 39266 19684 39268
rect 19708 39266 19764 39268
rect 19788 39266 19844 39268
rect 19868 39266 19924 39268
rect 19628 37988 19684 37990
rect 19708 37988 19764 37990
rect 19788 37988 19844 37990
rect 19868 37988 19924 37990
rect 19628 37936 19654 37988
rect 19654 37936 19684 37988
rect 19708 37936 19718 37988
rect 19718 37936 19764 37988
rect 19788 37936 19834 37988
rect 19834 37936 19844 37988
rect 19868 37936 19898 37988
rect 19898 37936 19924 37988
rect 19628 37934 19684 37936
rect 19708 37934 19764 37936
rect 19788 37934 19844 37936
rect 19868 37934 19924 37936
rect 19628 36656 19684 36658
rect 19708 36656 19764 36658
rect 19788 36656 19844 36658
rect 19868 36656 19924 36658
rect 19628 36604 19654 36656
rect 19654 36604 19684 36656
rect 19708 36604 19718 36656
rect 19718 36604 19764 36656
rect 19788 36604 19834 36656
rect 19834 36604 19844 36656
rect 19868 36604 19898 36656
rect 19898 36604 19924 36656
rect 19628 36602 19684 36604
rect 19708 36602 19764 36604
rect 19788 36602 19844 36604
rect 19868 36602 19924 36604
rect 19628 35324 19684 35326
rect 19708 35324 19764 35326
rect 19788 35324 19844 35326
rect 19868 35324 19924 35326
rect 19628 35272 19654 35324
rect 19654 35272 19684 35324
rect 19708 35272 19718 35324
rect 19718 35272 19764 35324
rect 19788 35272 19834 35324
rect 19834 35272 19844 35324
rect 19868 35272 19898 35324
rect 19898 35272 19924 35324
rect 19628 35270 19684 35272
rect 19708 35270 19764 35272
rect 19788 35270 19844 35272
rect 19868 35270 19924 35272
rect 19628 33992 19684 33994
rect 19708 33992 19764 33994
rect 19788 33992 19844 33994
rect 19868 33992 19924 33994
rect 19628 33940 19654 33992
rect 19654 33940 19684 33992
rect 19708 33940 19718 33992
rect 19718 33940 19764 33992
rect 19788 33940 19834 33992
rect 19834 33940 19844 33992
rect 19868 33940 19898 33992
rect 19898 33940 19924 33992
rect 19628 33938 19684 33940
rect 19708 33938 19764 33940
rect 19788 33938 19844 33940
rect 19868 33938 19924 33940
rect 19628 32660 19684 32662
rect 19708 32660 19764 32662
rect 19788 32660 19844 32662
rect 19868 32660 19924 32662
rect 19628 32608 19654 32660
rect 19654 32608 19684 32660
rect 19708 32608 19718 32660
rect 19718 32608 19764 32660
rect 19788 32608 19834 32660
rect 19834 32608 19844 32660
rect 19868 32608 19898 32660
rect 19898 32608 19924 32660
rect 19628 32606 19684 32608
rect 19708 32606 19764 32608
rect 19788 32606 19844 32608
rect 19868 32606 19924 32608
rect 19628 31328 19684 31330
rect 19708 31328 19764 31330
rect 19788 31328 19844 31330
rect 19868 31328 19924 31330
rect 19628 31276 19654 31328
rect 19654 31276 19684 31328
rect 19708 31276 19718 31328
rect 19718 31276 19764 31328
rect 19788 31276 19834 31328
rect 19834 31276 19844 31328
rect 19868 31276 19898 31328
rect 19898 31276 19924 31328
rect 19628 31274 19684 31276
rect 19708 31274 19764 31276
rect 19788 31274 19844 31276
rect 19868 31274 19924 31276
rect 19628 29996 19684 29998
rect 19708 29996 19764 29998
rect 19788 29996 19844 29998
rect 19868 29996 19924 29998
rect 19628 29944 19654 29996
rect 19654 29944 19684 29996
rect 19708 29944 19718 29996
rect 19718 29944 19764 29996
rect 19788 29944 19834 29996
rect 19834 29944 19844 29996
rect 19868 29944 19898 29996
rect 19898 29944 19924 29996
rect 19628 29942 19684 29944
rect 19708 29942 19764 29944
rect 19788 29942 19844 29944
rect 19868 29942 19924 29944
rect 19628 28664 19684 28666
rect 19708 28664 19764 28666
rect 19788 28664 19844 28666
rect 19868 28664 19924 28666
rect 19628 28612 19654 28664
rect 19654 28612 19684 28664
rect 19708 28612 19718 28664
rect 19718 28612 19764 28664
rect 19788 28612 19834 28664
rect 19834 28612 19844 28664
rect 19868 28612 19898 28664
rect 19898 28612 19924 28664
rect 19628 28610 19684 28612
rect 19708 28610 19764 28612
rect 19788 28610 19844 28612
rect 19868 28610 19924 28612
rect 19628 27332 19684 27334
rect 19708 27332 19764 27334
rect 19788 27332 19844 27334
rect 19868 27332 19924 27334
rect 19628 27280 19654 27332
rect 19654 27280 19684 27332
rect 19708 27280 19718 27332
rect 19718 27280 19764 27332
rect 19788 27280 19834 27332
rect 19834 27280 19844 27332
rect 19868 27280 19898 27332
rect 19898 27280 19924 27332
rect 19628 27278 19684 27280
rect 19708 27278 19764 27280
rect 19788 27278 19844 27280
rect 19868 27278 19924 27280
rect 19628 26000 19684 26002
rect 19708 26000 19764 26002
rect 19788 26000 19844 26002
rect 19868 26000 19924 26002
rect 19628 25948 19654 26000
rect 19654 25948 19684 26000
rect 19708 25948 19718 26000
rect 19718 25948 19764 26000
rect 19788 25948 19834 26000
rect 19834 25948 19844 26000
rect 19868 25948 19898 26000
rect 19898 25948 19924 26000
rect 19628 25946 19684 25948
rect 19708 25946 19764 25948
rect 19788 25946 19844 25948
rect 19868 25946 19924 25948
rect 19628 24668 19684 24670
rect 19708 24668 19764 24670
rect 19788 24668 19844 24670
rect 19868 24668 19924 24670
rect 19628 24616 19654 24668
rect 19654 24616 19684 24668
rect 19708 24616 19718 24668
rect 19718 24616 19764 24668
rect 19788 24616 19834 24668
rect 19834 24616 19844 24668
rect 19868 24616 19898 24668
rect 19898 24616 19924 24668
rect 19628 24614 19684 24616
rect 19708 24614 19764 24616
rect 19788 24614 19844 24616
rect 19868 24614 19924 24616
rect 19628 23336 19684 23338
rect 19708 23336 19764 23338
rect 19788 23336 19844 23338
rect 19868 23336 19924 23338
rect 19628 23284 19654 23336
rect 19654 23284 19684 23336
rect 19708 23284 19718 23336
rect 19718 23284 19764 23336
rect 19788 23284 19834 23336
rect 19834 23284 19844 23336
rect 19868 23284 19898 23336
rect 19898 23284 19924 23336
rect 19628 23282 19684 23284
rect 19708 23282 19764 23284
rect 19788 23282 19844 23284
rect 19868 23282 19924 23284
rect 19628 22004 19684 22006
rect 19708 22004 19764 22006
rect 19788 22004 19844 22006
rect 19868 22004 19924 22006
rect 19628 21952 19654 22004
rect 19654 21952 19684 22004
rect 19708 21952 19718 22004
rect 19718 21952 19764 22004
rect 19788 21952 19834 22004
rect 19834 21952 19844 22004
rect 19868 21952 19898 22004
rect 19898 21952 19924 22004
rect 19628 21950 19684 21952
rect 19708 21950 19764 21952
rect 19788 21950 19844 21952
rect 19868 21950 19924 21952
rect 19628 20672 19684 20674
rect 19708 20672 19764 20674
rect 19788 20672 19844 20674
rect 19868 20672 19924 20674
rect 19628 20620 19654 20672
rect 19654 20620 19684 20672
rect 19708 20620 19718 20672
rect 19718 20620 19764 20672
rect 19788 20620 19834 20672
rect 19834 20620 19844 20672
rect 19868 20620 19898 20672
rect 19898 20620 19924 20672
rect 19628 20618 19684 20620
rect 19708 20618 19764 20620
rect 19788 20618 19844 20620
rect 19868 20618 19924 20620
rect 19628 19340 19684 19342
rect 19708 19340 19764 19342
rect 19788 19340 19844 19342
rect 19868 19340 19924 19342
rect 19628 19288 19654 19340
rect 19654 19288 19684 19340
rect 19708 19288 19718 19340
rect 19718 19288 19764 19340
rect 19788 19288 19834 19340
rect 19834 19288 19844 19340
rect 19868 19288 19898 19340
rect 19898 19288 19924 19340
rect 19628 19286 19684 19288
rect 19708 19286 19764 19288
rect 19788 19286 19844 19288
rect 19868 19286 19924 19288
rect 19628 18008 19684 18010
rect 19708 18008 19764 18010
rect 19788 18008 19844 18010
rect 19868 18008 19924 18010
rect 19628 17956 19654 18008
rect 19654 17956 19684 18008
rect 19708 17956 19718 18008
rect 19718 17956 19764 18008
rect 19788 17956 19834 18008
rect 19834 17956 19844 18008
rect 19868 17956 19898 18008
rect 19898 17956 19924 18008
rect 19628 17954 19684 17956
rect 19708 17954 19764 17956
rect 19788 17954 19844 17956
rect 19868 17954 19924 17956
rect 19628 16676 19684 16678
rect 19708 16676 19764 16678
rect 19788 16676 19844 16678
rect 19868 16676 19924 16678
rect 19628 16624 19654 16676
rect 19654 16624 19684 16676
rect 19708 16624 19718 16676
rect 19718 16624 19764 16676
rect 19788 16624 19834 16676
rect 19834 16624 19844 16676
rect 19868 16624 19898 16676
rect 19898 16624 19924 16676
rect 19628 16622 19684 16624
rect 19708 16622 19764 16624
rect 19788 16622 19844 16624
rect 19868 16622 19924 16624
rect 19628 15344 19684 15346
rect 19708 15344 19764 15346
rect 19788 15344 19844 15346
rect 19868 15344 19924 15346
rect 19628 15292 19654 15344
rect 19654 15292 19684 15344
rect 19708 15292 19718 15344
rect 19718 15292 19764 15344
rect 19788 15292 19834 15344
rect 19834 15292 19844 15344
rect 19868 15292 19898 15344
rect 19898 15292 19924 15344
rect 19628 15290 19684 15292
rect 19708 15290 19764 15292
rect 19788 15290 19844 15292
rect 19868 15290 19924 15292
rect 19628 14012 19684 14014
rect 19708 14012 19764 14014
rect 19788 14012 19844 14014
rect 19868 14012 19924 14014
rect 19628 13960 19654 14012
rect 19654 13960 19684 14012
rect 19708 13960 19718 14012
rect 19718 13960 19764 14012
rect 19788 13960 19834 14012
rect 19834 13960 19844 14012
rect 19868 13960 19898 14012
rect 19898 13960 19924 14012
rect 19628 13958 19684 13960
rect 19708 13958 19764 13960
rect 19788 13958 19844 13960
rect 19868 13958 19924 13960
rect 19628 12680 19684 12682
rect 19708 12680 19764 12682
rect 19788 12680 19844 12682
rect 19868 12680 19924 12682
rect 19628 12628 19654 12680
rect 19654 12628 19684 12680
rect 19708 12628 19718 12680
rect 19718 12628 19764 12680
rect 19788 12628 19834 12680
rect 19834 12628 19844 12680
rect 19868 12628 19898 12680
rect 19898 12628 19924 12680
rect 19628 12626 19684 12628
rect 19708 12626 19764 12628
rect 19788 12626 19844 12628
rect 19868 12626 19924 12628
rect 19628 11348 19684 11350
rect 19708 11348 19764 11350
rect 19788 11348 19844 11350
rect 19868 11348 19924 11350
rect 19628 11296 19654 11348
rect 19654 11296 19684 11348
rect 19708 11296 19718 11348
rect 19718 11296 19764 11348
rect 19788 11296 19834 11348
rect 19834 11296 19844 11348
rect 19868 11296 19898 11348
rect 19898 11296 19924 11348
rect 19628 11294 19684 11296
rect 19708 11294 19764 11296
rect 19788 11294 19844 11296
rect 19868 11294 19924 11296
rect 19628 10016 19684 10018
rect 19708 10016 19764 10018
rect 19788 10016 19844 10018
rect 19868 10016 19924 10018
rect 19628 9964 19654 10016
rect 19654 9964 19684 10016
rect 19708 9964 19718 10016
rect 19718 9964 19764 10016
rect 19788 9964 19834 10016
rect 19834 9964 19844 10016
rect 19868 9964 19898 10016
rect 19898 9964 19924 10016
rect 19628 9962 19684 9964
rect 19708 9962 19764 9964
rect 19788 9962 19844 9964
rect 19868 9962 19924 9964
rect 19628 8684 19684 8686
rect 19708 8684 19764 8686
rect 19788 8684 19844 8686
rect 19868 8684 19924 8686
rect 19628 8632 19654 8684
rect 19654 8632 19684 8684
rect 19708 8632 19718 8684
rect 19718 8632 19764 8684
rect 19788 8632 19834 8684
rect 19834 8632 19844 8684
rect 19868 8632 19898 8684
rect 19898 8632 19924 8684
rect 19628 8630 19684 8632
rect 19708 8630 19764 8632
rect 19788 8630 19844 8632
rect 19868 8630 19924 8632
rect 19628 7352 19684 7354
rect 19708 7352 19764 7354
rect 19788 7352 19844 7354
rect 19868 7352 19924 7354
rect 19628 7300 19654 7352
rect 19654 7300 19684 7352
rect 19708 7300 19718 7352
rect 19718 7300 19764 7352
rect 19788 7300 19834 7352
rect 19834 7300 19844 7352
rect 19868 7300 19898 7352
rect 19898 7300 19924 7352
rect 19628 7298 19684 7300
rect 19708 7298 19764 7300
rect 19788 7298 19844 7300
rect 19868 7298 19924 7300
rect 19628 6020 19684 6022
rect 19708 6020 19764 6022
rect 19788 6020 19844 6022
rect 19868 6020 19924 6022
rect 19628 5968 19654 6020
rect 19654 5968 19684 6020
rect 19708 5968 19718 6020
rect 19718 5968 19764 6020
rect 19788 5968 19834 6020
rect 19834 5968 19844 6020
rect 19868 5968 19898 6020
rect 19898 5968 19924 6020
rect 19628 5966 19684 5968
rect 19708 5966 19764 5968
rect 19788 5966 19844 5968
rect 19868 5966 19924 5968
rect 19628 4688 19684 4690
rect 19708 4688 19764 4690
rect 19788 4688 19844 4690
rect 19868 4688 19924 4690
rect 19628 4636 19654 4688
rect 19654 4636 19684 4688
rect 19708 4636 19718 4688
rect 19718 4636 19764 4688
rect 19788 4636 19834 4688
rect 19834 4636 19844 4688
rect 19868 4636 19898 4688
rect 19898 4636 19924 4688
rect 19628 4634 19684 4636
rect 19708 4634 19764 4636
rect 19788 4634 19844 4636
rect 19868 4634 19924 4636
rect 19892 3467 19948 3506
rect 19892 3450 19894 3467
rect 19894 3450 19946 3467
rect 19946 3450 19948 3467
rect 19628 3356 19684 3358
rect 19708 3356 19764 3358
rect 19788 3356 19844 3358
rect 19868 3356 19924 3358
rect 19628 3304 19654 3356
rect 19654 3304 19684 3356
rect 19708 3304 19718 3356
rect 19718 3304 19764 3356
rect 19788 3304 19834 3356
rect 19834 3304 19844 3356
rect 19868 3304 19898 3356
rect 19898 3304 19924 3356
rect 19628 3302 19684 3304
rect 19708 3302 19764 3304
rect 19788 3302 19844 3304
rect 19868 3302 19924 3304
rect 19796 3154 19852 3210
rect 34988 57302 35044 57304
rect 35068 57302 35124 57304
rect 35148 57302 35204 57304
rect 35228 57302 35284 57304
rect 34988 57250 35014 57302
rect 35014 57250 35044 57302
rect 35068 57250 35078 57302
rect 35078 57250 35124 57302
rect 35148 57250 35194 57302
rect 35194 57250 35204 57302
rect 35228 57250 35258 57302
rect 35258 57250 35284 57302
rect 34988 57248 35044 57250
rect 35068 57248 35124 57250
rect 35148 57248 35204 57250
rect 35228 57248 35284 57250
rect 33524 3746 33580 3802
rect 33716 3302 33772 3358
rect 34988 55970 35044 55972
rect 35068 55970 35124 55972
rect 35148 55970 35204 55972
rect 35228 55970 35284 55972
rect 34988 55918 35014 55970
rect 35014 55918 35044 55970
rect 35068 55918 35078 55970
rect 35078 55918 35124 55970
rect 35148 55918 35194 55970
rect 35194 55918 35204 55970
rect 35228 55918 35258 55970
rect 35258 55918 35284 55970
rect 34988 55916 35044 55918
rect 35068 55916 35124 55918
rect 35148 55916 35204 55918
rect 35228 55916 35284 55918
rect 34988 54638 35044 54640
rect 35068 54638 35124 54640
rect 35148 54638 35204 54640
rect 35228 54638 35284 54640
rect 34988 54586 35014 54638
rect 35014 54586 35044 54638
rect 35068 54586 35078 54638
rect 35078 54586 35124 54638
rect 35148 54586 35194 54638
rect 35194 54586 35204 54638
rect 35228 54586 35258 54638
rect 35258 54586 35284 54638
rect 34988 54584 35044 54586
rect 35068 54584 35124 54586
rect 35148 54584 35204 54586
rect 35228 54584 35284 54586
rect 34988 53306 35044 53308
rect 35068 53306 35124 53308
rect 35148 53306 35204 53308
rect 35228 53306 35284 53308
rect 34988 53254 35014 53306
rect 35014 53254 35044 53306
rect 35068 53254 35078 53306
rect 35078 53254 35124 53306
rect 35148 53254 35194 53306
rect 35194 53254 35204 53306
rect 35228 53254 35258 53306
rect 35258 53254 35284 53306
rect 34988 53252 35044 53254
rect 35068 53252 35124 53254
rect 35148 53252 35204 53254
rect 35228 53252 35284 53254
rect 34988 51974 35044 51976
rect 35068 51974 35124 51976
rect 35148 51974 35204 51976
rect 35228 51974 35284 51976
rect 34988 51922 35014 51974
rect 35014 51922 35044 51974
rect 35068 51922 35078 51974
rect 35078 51922 35124 51974
rect 35148 51922 35194 51974
rect 35194 51922 35204 51974
rect 35228 51922 35258 51974
rect 35258 51922 35284 51974
rect 34988 51920 35044 51922
rect 35068 51920 35124 51922
rect 35148 51920 35204 51922
rect 35228 51920 35284 51922
rect 34988 50642 35044 50644
rect 35068 50642 35124 50644
rect 35148 50642 35204 50644
rect 35228 50642 35284 50644
rect 34988 50590 35014 50642
rect 35014 50590 35044 50642
rect 35068 50590 35078 50642
rect 35078 50590 35124 50642
rect 35148 50590 35194 50642
rect 35194 50590 35204 50642
rect 35228 50590 35258 50642
rect 35258 50590 35284 50642
rect 34988 50588 35044 50590
rect 35068 50588 35124 50590
rect 35148 50588 35204 50590
rect 35228 50588 35284 50590
rect 34988 49310 35044 49312
rect 35068 49310 35124 49312
rect 35148 49310 35204 49312
rect 35228 49310 35284 49312
rect 34988 49258 35014 49310
rect 35014 49258 35044 49310
rect 35068 49258 35078 49310
rect 35078 49258 35124 49310
rect 35148 49258 35194 49310
rect 35194 49258 35204 49310
rect 35228 49258 35258 49310
rect 35258 49258 35284 49310
rect 34988 49256 35044 49258
rect 35068 49256 35124 49258
rect 35148 49256 35204 49258
rect 35228 49256 35284 49258
rect 34988 47978 35044 47980
rect 35068 47978 35124 47980
rect 35148 47978 35204 47980
rect 35228 47978 35284 47980
rect 34988 47926 35014 47978
rect 35014 47926 35044 47978
rect 35068 47926 35078 47978
rect 35078 47926 35124 47978
rect 35148 47926 35194 47978
rect 35194 47926 35204 47978
rect 35228 47926 35258 47978
rect 35258 47926 35284 47978
rect 34988 47924 35044 47926
rect 35068 47924 35124 47926
rect 35148 47924 35204 47926
rect 35228 47924 35284 47926
rect 34988 46646 35044 46648
rect 35068 46646 35124 46648
rect 35148 46646 35204 46648
rect 35228 46646 35284 46648
rect 34988 46594 35014 46646
rect 35014 46594 35044 46646
rect 35068 46594 35078 46646
rect 35078 46594 35124 46646
rect 35148 46594 35194 46646
rect 35194 46594 35204 46646
rect 35228 46594 35258 46646
rect 35258 46594 35284 46646
rect 34988 46592 35044 46594
rect 35068 46592 35124 46594
rect 35148 46592 35204 46594
rect 35228 46592 35284 46594
rect 34988 45314 35044 45316
rect 35068 45314 35124 45316
rect 35148 45314 35204 45316
rect 35228 45314 35284 45316
rect 34988 45262 35014 45314
rect 35014 45262 35044 45314
rect 35068 45262 35078 45314
rect 35078 45262 35124 45314
rect 35148 45262 35194 45314
rect 35194 45262 35204 45314
rect 35228 45262 35258 45314
rect 35258 45262 35284 45314
rect 34988 45260 35044 45262
rect 35068 45260 35124 45262
rect 35148 45260 35204 45262
rect 35228 45260 35284 45262
rect 34988 43982 35044 43984
rect 35068 43982 35124 43984
rect 35148 43982 35204 43984
rect 35228 43982 35284 43984
rect 34988 43930 35014 43982
rect 35014 43930 35044 43982
rect 35068 43930 35078 43982
rect 35078 43930 35124 43982
rect 35148 43930 35194 43982
rect 35194 43930 35204 43982
rect 35228 43930 35258 43982
rect 35258 43930 35284 43982
rect 34988 43928 35044 43930
rect 35068 43928 35124 43930
rect 35148 43928 35204 43930
rect 35228 43928 35284 43930
rect 34988 42650 35044 42652
rect 35068 42650 35124 42652
rect 35148 42650 35204 42652
rect 35228 42650 35284 42652
rect 34988 42598 35014 42650
rect 35014 42598 35044 42650
rect 35068 42598 35078 42650
rect 35078 42598 35124 42650
rect 35148 42598 35194 42650
rect 35194 42598 35204 42650
rect 35228 42598 35258 42650
rect 35258 42598 35284 42650
rect 34988 42596 35044 42598
rect 35068 42596 35124 42598
rect 35148 42596 35204 42598
rect 35228 42596 35284 42598
rect 34988 41318 35044 41320
rect 35068 41318 35124 41320
rect 35148 41318 35204 41320
rect 35228 41318 35284 41320
rect 34988 41266 35014 41318
rect 35014 41266 35044 41318
rect 35068 41266 35078 41318
rect 35078 41266 35124 41318
rect 35148 41266 35194 41318
rect 35194 41266 35204 41318
rect 35228 41266 35258 41318
rect 35258 41266 35284 41318
rect 34988 41264 35044 41266
rect 35068 41264 35124 41266
rect 35148 41264 35204 41266
rect 35228 41264 35284 41266
rect 34988 39986 35044 39988
rect 35068 39986 35124 39988
rect 35148 39986 35204 39988
rect 35228 39986 35284 39988
rect 34988 39934 35014 39986
rect 35014 39934 35044 39986
rect 35068 39934 35078 39986
rect 35078 39934 35124 39986
rect 35148 39934 35194 39986
rect 35194 39934 35204 39986
rect 35228 39934 35258 39986
rect 35258 39934 35284 39986
rect 34988 39932 35044 39934
rect 35068 39932 35124 39934
rect 35148 39932 35204 39934
rect 35228 39932 35284 39934
rect 34988 38654 35044 38656
rect 35068 38654 35124 38656
rect 35148 38654 35204 38656
rect 35228 38654 35284 38656
rect 34988 38602 35014 38654
rect 35014 38602 35044 38654
rect 35068 38602 35078 38654
rect 35078 38602 35124 38654
rect 35148 38602 35194 38654
rect 35194 38602 35204 38654
rect 35228 38602 35258 38654
rect 35258 38602 35284 38654
rect 34988 38600 35044 38602
rect 35068 38600 35124 38602
rect 35148 38600 35204 38602
rect 35228 38600 35284 38602
rect 34988 37322 35044 37324
rect 35068 37322 35124 37324
rect 35148 37322 35204 37324
rect 35228 37322 35284 37324
rect 34988 37270 35014 37322
rect 35014 37270 35044 37322
rect 35068 37270 35078 37322
rect 35078 37270 35124 37322
rect 35148 37270 35194 37322
rect 35194 37270 35204 37322
rect 35228 37270 35258 37322
rect 35258 37270 35284 37322
rect 34988 37268 35044 37270
rect 35068 37268 35124 37270
rect 35148 37268 35204 37270
rect 35228 37268 35284 37270
rect 34988 35990 35044 35992
rect 35068 35990 35124 35992
rect 35148 35990 35204 35992
rect 35228 35990 35284 35992
rect 34988 35938 35014 35990
rect 35014 35938 35044 35990
rect 35068 35938 35078 35990
rect 35078 35938 35124 35990
rect 35148 35938 35194 35990
rect 35194 35938 35204 35990
rect 35228 35938 35258 35990
rect 35258 35938 35284 35990
rect 34988 35936 35044 35938
rect 35068 35936 35124 35938
rect 35148 35936 35204 35938
rect 35228 35936 35284 35938
rect 34988 34658 35044 34660
rect 35068 34658 35124 34660
rect 35148 34658 35204 34660
rect 35228 34658 35284 34660
rect 34988 34606 35014 34658
rect 35014 34606 35044 34658
rect 35068 34606 35078 34658
rect 35078 34606 35124 34658
rect 35148 34606 35194 34658
rect 35194 34606 35204 34658
rect 35228 34606 35258 34658
rect 35258 34606 35284 34658
rect 34988 34604 35044 34606
rect 35068 34604 35124 34606
rect 35148 34604 35204 34606
rect 35228 34604 35284 34606
rect 34988 33326 35044 33328
rect 35068 33326 35124 33328
rect 35148 33326 35204 33328
rect 35228 33326 35284 33328
rect 34988 33274 35014 33326
rect 35014 33274 35044 33326
rect 35068 33274 35078 33326
rect 35078 33274 35124 33326
rect 35148 33274 35194 33326
rect 35194 33274 35204 33326
rect 35228 33274 35258 33326
rect 35258 33274 35284 33326
rect 34988 33272 35044 33274
rect 35068 33272 35124 33274
rect 35148 33272 35204 33274
rect 35228 33272 35284 33274
rect 34988 31994 35044 31996
rect 35068 31994 35124 31996
rect 35148 31994 35204 31996
rect 35228 31994 35284 31996
rect 34988 31942 35014 31994
rect 35014 31942 35044 31994
rect 35068 31942 35078 31994
rect 35078 31942 35124 31994
rect 35148 31942 35194 31994
rect 35194 31942 35204 31994
rect 35228 31942 35258 31994
rect 35258 31942 35284 31994
rect 34988 31940 35044 31942
rect 35068 31940 35124 31942
rect 35148 31940 35204 31942
rect 35228 31940 35284 31942
rect 34988 30662 35044 30664
rect 35068 30662 35124 30664
rect 35148 30662 35204 30664
rect 35228 30662 35284 30664
rect 34988 30610 35014 30662
rect 35014 30610 35044 30662
rect 35068 30610 35078 30662
rect 35078 30610 35124 30662
rect 35148 30610 35194 30662
rect 35194 30610 35204 30662
rect 35228 30610 35258 30662
rect 35258 30610 35284 30662
rect 34988 30608 35044 30610
rect 35068 30608 35124 30610
rect 35148 30608 35204 30610
rect 35228 30608 35284 30610
rect 34988 29330 35044 29332
rect 35068 29330 35124 29332
rect 35148 29330 35204 29332
rect 35228 29330 35284 29332
rect 34988 29278 35014 29330
rect 35014 29278 35044 29330
rect 35068 29278 35078 29330
rect 35078 29278 35124 29330
rect 35148 29278 35194 29330
rect 35194 29278 35204 29330
rect 35228 29278 35258 29330
rect 35258 29278 35284 29330
rect 34988 29276 35044 29278
rect 35068 29276 35124 29278
rect 35148 29276 35204 29278
rect 35228 29276 35284 29278
rect 34988 27998 35044 28000
rect 35068 27998 35124 28000
rect 35148 27998 35204 28000
rect 35228 27998 35284 28000
rect 34988 27946 35014 27998
rect 35014 27946 35044 27998
rect 35068 27946 35078 27998
rect 35078 27946 35124 27998
rect 35148 27946 35194 27998
rect 35194 27946 35204 27998
rect 35228 27946 35258 27998
rect 35258 27946 35284 27998
rect 34988 27944 35044 27946
rect 35068 27944 35124 27946
rect 35148 27944 35204 27946
rect 35228 27944 35284 27946
rect 34988 26666 35044 26668
rect 35068 26666 35124 26668
rect 35148 26666 35204 26668
rect 35228 26666 35284 26668
rect 34988 26614 35014 26666
rect 35014 26614 35044 26666
rect 35068 26614 35078 26666
rect 35078 26614 35124 26666
rect 35148 26614 35194 26666
rect 35194 26614 35204 26666
rect 35228 26614 35258 26666
rect 35258 26614 35284 26666
rect 34988 26612 35044 26614
rect 35068 26612 35124 26614
rect 35148 26612 35204 26614
rect 35228 26612 35284 26614
rect 34988 25334 35044 25336
rect 35068 25334 35124 25336
rect 35148 25334 35204 25336
rect 35228 25334 35284 25336
rect 34988 25282 35014 25334
rect 35014 25282 35044 25334
rect 35068 25282 35078 25334
rect 35078 25282 35124 25334
rect 35148 25282 35194 25334
rect 35194 25282 35204 25334
rect 35228 25282 35258 25334
rect 35258 25282 35284 25334
rect 34988 25280 35044 25282
rect 35068 25280 35124 25282
rect 35148 25280 35204 25282
rect 35228 25280 35284 25282
rect 34988 24002 35044 24004
rect 35068 24002 35124 24004
rect 35148 24002 35204 24004
rect 35228 24002 35284 24004
rect 34988 23950 35014 24002
rect 35014 23950 35044 24002
rect 35068 23950 35078 24002
rect 35078 23950 35124 24002
rect 35148 23950 35194 24002
rect 35194 23950 35204 24002
rect 35228 23950 35258 24002
rect 35258 23950 35284 24002
rect 34988 23948 35044 23950
rect 35068 23948 35124 23950
rect 35148 23948 35204 23950
rect 35228 23948 35284 23950
rect 34988 22670 35044 22672
rect 35068 22670 35124 22672
rect 35148 22670 35204 22672
rect 35228 22670 35284 22672
rect 34988 22618 35014 22670
rect 35014 22618 35044 22670
rect 35068 22618 35078 22670
rect 35078 22618 35124 22670
rect 35148 22618 35194 22670
rect 35194 22618 35204 22670
rect 35228 22618 35258 22670
rect 35258 22618 35284 22670
rect 34988 22616 35044 22618
rect 35068 22616 35124 22618
rect 35148 22616 35204 22618
rect 35228 22616 35284 22618
rect 34988 21338 35044 21340
rect 35068 21338 35124 21340
rect 35148 21338 35204 21340
rect 35228 21338 35284 21340
rect 34988 21286 35014 21338
rect 35014 21286 35044 21338
rect 35068 21286 35078 21338
rect 35078 21286 35124 21338
rect 35148 21286 35194 21338
rect 35194 21286 35204 21338
rect 35228 21286 35258 21338
rect 35258 21286 35284 21338
rect 34988 21284 35044 21286
rect 35068 21284 35124 21286
rect 35148 21284 35204 21286
rect 35228 21284 35284 21286
rect 34988 20006 35044 20008
rect 35068 20006 35124 20008
rect 35148 20006 35204 20008
rect 35228 20006 35284 20008
rect 34988 19954 35014 20006
rect 35014 19954 35044 20006
rect 35068 19954 35078 20006
rect 35078 19954 35124 20006
rect 35148 19954 35194 20006
rect 35194 19954 35204 20006
rect 35228 19954 35258 20006
rect 35258 19954 35284 20006
rect 34988 19952 35044 19954
rect 35068 19952 35124 19954
rect 35148 19952 35204 19954
rect 35228 19952 35284 19954
rect 34988 18674 35044 18676
rect 35068 18674 35124 18676
rect 35148 18674 35204 18676
rect 35228 18674 35284 18676
rect 34988 18622 35014 18674
rect 35014 18622 35044 18674
rect 35068 18622 35078 18674
rect 35078 18622 35124 18674
rect 35148 18622 35194 18674
rect 35194 18622 35204 18674
rect 35228 18622 35258 18674
rect 35258 18622 35284 18674
rect 34988 18620 35044 18622
rect 35068 18620 35124 18622
rect 35148 18620 35204 18622
rect 35228 18620 35284 18622
rect 34988 17342 35044 17344
rect 35068 17342 35124 17344
rect 35148 17342 35204 17344
rect 35228 17342 35284 17344
rect 34988 17290 35014 17342
rect 35014 17290 35044 17342
rect 35068 17290 35078 17342
rect 35078 17290 35124 17342
rect 35148 17290 35194 17342
rect 35194 17290 35204 17342
rect 35228 17290 35258 17342
rect 35258 17290 35284 17342
rect 34988 17288 35044 17290
rect 35068 17288 35124 17290
rect 35148 17288 35204 17290
rect 35228 17288 35284 17290
rect 34988 16010 35044 16012
rect 35068 16010 35124 16012
rect 35148 16010 35204 16012
rect 35228 16010 35284 16012
rect 34988 15958 35014 16010
rect 35014 15958 35044 16010
rect 35068 15958 35078 16010
rect 35078 15958 35124 16010
rect 35148 15958 35194 16010
rect 35194 15958 35204 16010
rect 35228 15958 35258 16010
rect 35258 15958 35284 16010
rect 34988 15956 35044 15958
rect 35068 15956 35124 15958
rect 35148 15956 35204 15958
rect 35228 15956 35284 15958
rect 34988 14678 35044 14680
rect 35068 14678 35124 14680
rect 35148 14678 35204 14680
rect 35228 14678 35284 14680
rect 34988 14626 35014 14678
rect 35014 14626 35044 14678
rect 35068 14626 35078 14678
rect 35078 14626 35124 14678
rect 35148 14626 35194 14678
rect 35194 14626 35204 14678
rect 35228 14626 35258 14678
rect 35258 14626 35284 14678
rect 34988 14624 35044 14626
rect 35068 14624 35124 14626
rect 35148 14624 35204 14626
rect 35228 14624 35284 14626
rect 34988 13346 35044 13348
rect 35068 13346 35124 13348
rect 35148 13346 35204 13348
rect 35228 13346 35284 13348
rect 34988 13294 35014 13346
rect 35014 13294 35044 13346
rect 35068 13294 35078 13346
rect 35078 13294 35124 13346
rect 35148 13294 35194 13346
rect 35194 13294 35204 13346
rect 35228 13294 35258 13346
rect 35258 13294 35284 13346
rect 34988 13292 35044 13294
rect 35068 13292 35124 13294
rect 35148 13292 35204 13294
rect 35228 13292 35284 13294
rect 34988 12014 35044 12016
rect 35068 12014 35124 12016
rect 35148 12014 35204 12016
rect 35228 12014 35284 12016
rect 34988 11962 35014 12014
rect 35014 11962 35044 12014
rect 35068 11962 35078 12014
rect 35078 11962 35124 12014
rect 35148 11962 35194 12014
rect 35194 11962 35204 12014
rect 35228 11962 35258 12014
rect 35258 11962 35284 12014
rect 34988 11960 35044 11962
rect 35068 11960 35124 11962
rect 35148 11960 35204 11962
rect 35228 11960 35284 11962
rect 34988 10682 35044 10684
rect 35068 10682 35124 10684
rect 35148 10682 35204 10684
rect 35228 10682 35284 10684
rect 34988 10630 35014 10682
rect 35014 10630 35044 10682
rect 35068 10630 35078 10682
rect 35078 10630 35124 10682
rect 35148 10630 35194 10682
rect 35194 10630 35204 10682
rect 35228 10630 35258 10682
rect 35258 10630 35284 10682
rect 34988 10628 35044 10630
rect 35068 10628 35124 10630
rect 35148 10628 35204 10630
rect 35228 10628 35284 10630
rect 34988 9350 35044 9352
rect 35068 9350 35124 9352
rect 35148 9350 35204 9352
rect 35228 9350 35284 9352
rect 34988 9298 35014 9350
rect 35014 9298 35044 9350
rect 35068 9298 35078 9350
rect 35078 9298 35124 9350
rect 35148 9298 35194 9350
rect 35194 9298 35204 9350
rect 35228 9298 35258 9350
rect 35258 9298 35284 9350
rect 34988 9296 35044 9298
rect 35068 9296 35124 9298
rect 35148 9296 35204 9298
rect 35228 9296 35284 9298
rect 34988 8018 35044 8020
rect 35068 8018 35124 8020
rect 35148 8018 35204 8020
rect 35228 8018 35284 8020
rect 34988 7966 35014 8018
rect 35014 7966 35044 8018
rect 35068 7966 35078 8018
rect 35078 7966 35124 8018
rect 35148 7966 35194 8018
rect 35194 7966 35204 8018
rect 35228 7966 35258 8018
rect 35258 7966 35284 8018
rect 34988 7964 35044 7966
rect 35068 7964 35124 7966
rect 35148 7964 35204 7966
rect 35228 7964 35284 7966
rect 34988 6686 35044 6688
rect 35068 6686 35124 6688
rect 35148 6686 35204 6688
rect 35228 6686 35284 6688
rect 34988 6634 35014 6686
rect 35014 6634 35044 6686
rect 35068 6634 35078 6686
rect 35078 6634 35124 6686
rect 35148 6634 35194 6686
rect 35194 6634 35204 6686
rect 35228 6634 35258 6686
rect 35258 6634 35284 6686
rect 34988 6632 35044 6634
rect 35068 6632 35124 6634
rect 35148 6632 35204 6634
rect 35228 6632 35284 6634
rect 34988 5354 35044 5356
rect 35068 5354 35124 5356
rect 35148 5354 35204 5356
rect 35228 5354 35284 5356
rect 34988 5302 35014 5354
rect 35014 5302 35044 5354
rect 35068 5302 35078 5354
rect 35078 5302 35124 5354
rect 35148 5302 35194 5354
rect 35194 5302 35204 5354
rect 35228 5302 35258 5354
rect 35258 5302 35284 5354
rect 34988 5300 35044 5302
rect 35068 5300 35124 5302
rect 35148 5300 35204 5302
rect 35228 5300 35284 5302
rect 34988 4022 35044 4024
rect 35068 4022 35124 4024
rect 35148 4022 35204 4024
rect 35228 4022 35284 4024
rect 34988 3970 35014 4022
rect 35014 3970 35044 4022
rect 35068 3970 35078 4022
rect 35078 3970 35124 4022
rect 35148 3970 35194 4022
rect 35194 3970 35204 4022
rect 35228 3970 35258 4022
rect 35258 3970 35284 4022
rect 34988 3968 35044 3970
rect 35068 3968 35124 3970
rect 35148 3968 35204 3970
rect 35228 3968 35284 3970
rect 34988 2690 35044 2692
rect 35068 2690 35124 2692
rect 35148 2690 35204 2692
rect 35228 2690 35284 2692
rect 34988 2638 35014 2690
rect 35014 2638 35044 2690
rect 35068 2638 35078 2690
rect 35078 2638 35124 2690
rect 35148 2638 35194 2690
rect 35194 2638 35204 2690
rect 35228 2638 35258 2690
rect 35258 2638 35284 2690
rect 34988 2636 35044 2638
rect 35068 2636 35124 2638
rect 35148 2636 35204 2638
rect 35228 2636 35284 2638
rect 35636 3006 35692 3062
rect 35540 2414 35596 2470
rect 44276 3154 44332 3210
rect 44276 2858 44332 2914
rect 50348 56636 50404 56638
rect 50428 56636 50484 56638
rect 50508 56636 50564 56638
rect 50588 56636 50644 56638
rect 50348 56584 50374 56636
rect 50374 56584 50404 56636
rect 50428 56584 50438 56636
rect 50438 56584 50484 56636
rect 50508 56584 50554 56636
rect 50554 56584 50564 56636
rect 50588 56584 50618 56636
rect 50618 56584 50644 56636
rect 50348 56582 50404 56584
rect 50428 56582 50484 56584
rect 50508 56582 50564 56584
rect 50588 56582 50644 56584
rect 50348 55304 50404 55306
rect 50428 55304 50484 55306
rect 50508 55304 50564 55306
rect 50588 55304 50644 55306
rect 50348 55252 50374 55304
rect 50374 55252 50404 55304
rect 50428 55252 50438 55304
rect 50438 55252 50484 55304
rect 50508 55252 50554 55304
rect 50554 55252 50564 55304
rect 50588 55252 50618 55304
rect 50618 55252 50644 55304
rect 50348 55250 50404 55252
rect 50428 55250 50484 55252
rect 50508 55250 50564 55252
rect 50588 55250 50644 55252
rect 50348 53972 50404 53974
rect 50428 53972 50484 53974
rect 50508 53972 50564 53974
rect 50588 53972 50644 53974
rect 50348 53920 50374 53972
rect 50374 53920 50404 53972
rect 50428 53920 50438 53972
rect 50438 53920 50484 53972
rect 50508 53920 50554 53972
rect 50554 53920 50564 53972
rect 50588 53920 50618 53972
rect 50618 53920 50644 53972
rect 50348 53918 50404 53920
rect 50428 53918 50484 53920
rect 50508 53918 50564 53920
rect 50588 53918 50644 53920
rect 50348 52640 50404 52642
rect 50428 52640 50484 52642
rect 50508 52640 50564 52642
rect 50588 52640 50644 52642
rect 50348 52588 50374 52640
rect 50374 52588 50404 52640
rect 50428 52588 50438 52640
rect 50438 52588 50484 52640
rect 50508 52588 50554 52640
rect 50554 52588 50564 52640
rect 50588 52588 50618 52640
rect 50618 52588 50644 52640
rect 50348 52586 50404 52588
rect 50428 52586 50484 52588
rect 50508 52586 50564 52588
rect 50588 52586 50644 52588
rect 50348 51308 50404 51310
rect 50428 51308 50484 51310
rect 50508 51308 50564 51310
rect 50588 51308 50644 51310
rect 50348 51256 50374 51308
rect 50374 51256 50404 51308
rect 50428 51256 50438 51308
rect 50438 51256 50484 51308
rect 50508 51256 50554 51308
rect 50554 51256 50564 51308
rect 50588 51256 50618 51308
rect 50618 51256 50644 51308
rect 50348 51254 50404 51256
rect 50428 51254 50484 51256
rect 50508 51254 50564 51256
rect 50588 51254 50644 51256
rect 50348 49976 50404 49978
rect 50428 49976 50484 49978
rect 50508 49976 50564 49978
rect 50588 49976 50644 49978
rect 50348 49924 50374 49976
rect 50374 49924 50404 49976
rect 50428 49924 50438 49976
rect 50438 49924 50484 49976
rect 50508 49924 50554 49976
rect 50554 49924 50564 49976
rect 50588 49924 50618 49976
rect 50618 49924 50644 49976
rect 50348 49922 50404 49924
rect 50428 49922 50484 49924
rect 50508 49922 50564 49924
rect 50588 49922 50644 49924
rect 50348 48644 50404 48646
rect 50428 48644 50484 48646
rect 50508 48644 50564 48646
rect 50588 48644 50644 48646
rect 50348 48592 50374 48644
rect 50374 48592 50404 48644
rect 50428 48592 50438 48644
rect 50438 48592 50484 48644
rect 50508 48592 50554 48644
rect 50554 48592 50564 48644
rect 50588 48592 50618 48644
rect 50618 48592 50644 48644
rect 50348 48590 50404 48592
rect 50428 48590 50484 48592
rect 50508 48590 50564 48592
rect 50588 48590 50644 48592
rect 50348 47312 50404 47314
rect 50428 47312 50484 47314
rect 50508 47312 50564 47314
rect 50588 47312 50644 47314
rect 50348 47260 50374 47312
rect 50374 47260 50404 47312
rect 50428 47260 50438 47312
rect 50438 47260 50484 47312
rect 50508 47260 50554 47312
rect 50554 47260 50564 47312
rect 50588 47260 50618 47312
rect 50618 47260 50644 47312
rect 50348 47258 50404 47260
rect 50428 47258 50484 47260
rect 50508 47258 50564 47260
rect 50588 47258 50644 47260
rect 50348 45980 50404 45982
rect 50428 45980 50484 45982
rect 50508 45980 50564 45982
rect 50588 45980 50644 45982
rect 50348 45928 50374 45980
rect 50374 45928 50404 45980
rect 50428 45928 50438 45980
rect 50438 45928 50484 45980
rect 50508 45928 50554 45980
rect 50554 45928 50564 45980
rect 50588 45928 50618 45980
rect 50618 45928 50644 45980
rect 50348 45926 50404 45928
rect 50428 45926 50484 45928
rect 50508 45926 50564 45928
rect 50588 45926 50644 45928
rect 50348 44648 50404 44650
rect 50428 44648 50484 44650
rect 50508 44648 50564 44650
rect 50588 44648 50644 44650
rect 50348 44596 50374 44648
rect 50374 44596 50404 44648
rect 50428 44596 50438 44648
rect 50438 44596 50484 44648
rect 50508 44596 50554 44648
rect 50554 44596 50564 44648
rect 50588 44596 50618 44648
rect 50618 44596 50644 44648
rect 50348 44594 50404 44596
rect 50428 44594 50484 44596
rect 50508 44594 50564 44596
rect 50588 44594 50644 44596
rect 50348 43316 50404 43318
rect 50428 43316 50484 43318
rect 50508 43316 50564 43318
rect 50588 43316 50644 43318
rect 50348 43264 50374 43316
rect 50374 43264 50404 43316
rect 50428 43264 50438 43316
rect 50438 43264 50484 43316
rect 50508 43264 50554 43316
rect 50554 43264 50564 43316
rect 50588 43264 50618 43316
rect 50618 43264 50644 43316
rect 50348 43262 50404 43264
rect 50428 43262 50484 43264
rect 50508 43262 50564 43264
rect 50588 43262 50644 43264
rect 50348 41984 50404 41986
rect 50428 41984 50484 41986
rect 50508 41984 50564 41986
rect 50588 41984 50644 41986
rect 50348 41932 50374 41984
rect 50374 41932 50404 41984
rect 50428 41932 50438 41984
rect 50438 41932 50484 41984
rect 50508 41932 50554 41984
rect 50554 41932 50564 41984
rect 50588 41932 50618 41984
rect 50618 41932 50644 41984
rect 50348 41930 50404 41932
rect 50428 41930 50484 41932
rect 50508 41930 50564 41932
rect 50588 41930 50644 41932
rect 50348 40652 50404 40654
rect 50428 40652 50484 40654
rect 50508 40652 50564 40654
rect 50588 40652 50644 40654
rect 50348 40600 50374 40652
rect 50374 40600 50404 40652
rect 50428 40600 50438 40652
rect 50438 40600 50484 40652
rect 50508 40600 50554 40652
rect 50554 40600 50564 40652
rect 50588 40600 50618 40652
rect 50618 40600 50644 40652
rect 50348 40598 50404 40600
rect 50428 40598 50484 40600
rect 50508 40598 50564 40600
rect 50588 40598 50644 40600
rect 50348 39320 50404 39322
rect 50428 39320 50484 39322
rect 50508 39320 50564 39322
rect 50588 39320 50644 39322
rect 50348 39268 50374 39320
rect 50374 39268 50404 39320
rect 50428 39268 50438 39320
rect 50438 39268 50484 39320
rect 50508 39268 50554 39320
rect 50554 39268 50564 39320
rect 50588 39268 50618 39320
rect 50618 39268 50644 39320
rect 50348 39266 50404 39268
rect 50428 39266 50484 39268
rect 50508 39266 50564 39268
rect 50588 39266 50644 39268
rect 50348 37988 50404 37990
rect 50428 37988 50484 37990
rect 50508 37988 50564 37990
rect 50588 37988 50644 37990
rect 50348 37936 50374 37988
rect 50374 37936 50404 37988
rect 50428 37936 50438 37988
rect 50438 37936 50484 37988
rect 50508 37936 50554 37988
rect 50554 37936 50564 37988
rect 50588 37936 50618 37988
rect 50618 37936 50644 37988
rect 50348 37934 50404 37936
rect 50428 37934 50484 37936
rect 50508 37934 50564 37936
rect 50588 37934 50644 37936
rect 50348 36656 50404 36658
rect 50428 36656 50484 36658
rect 50508 36656 50564 36658
rect 50588 36656 50644 36658
rect 50348 36604 50374 36656
rect 50374 36604 50404 36656
rect 50428 36604 50438 36656
rect 50438 36604 50484 36656
rect 50508 36604 50554 36656
rect 50554 36604 50564 36656
rect 50588 36604 50618 36656
rect 50618 36604 50644 36656
rect 50348 36602 50404 36604
rect 50428 36602 50484 36604
rect 50508 36602 50564 36604
rect 50588 36602 50644 36604
rect 50348 35324 50404 35326
rect 50428 35324 50484 35326
rect 50508 35324 50564 35326
rect 50588 35324 50644 35326
rect 50348 35272 50374 35324
rect 50374 35272 50404 35324
rect 50428 35272 50438 35324
rect 50438 35272 50484 35324
rect 50508 35272 50554 35324
rect 50554 35272 50564 35324
rect 50588 35272 50618 35324
rect 50618 35272 50644 35324
rect 50348 35270 50404 35272
rect 50428 35270 50484 35272
rect 50508 35270 50564 35272
rect 50588 35270 50644 35272
rect 50348 33992 50404 33994
rect 50428 33992 50484 33994
rect 50508 33992 50564 33994
rect 50588 33992 50644 33994
rect 50348 33940 50374 33992
rect 50374 33940 50404 33992
rect 50428 33940 50438 33992
rect 50438 33940 50484 33992
rect 50508 33940 50554 33992
rect 50554 33940 50564 33992
rect 50588 33940 50618 33992
rect 50618 33940 50644 33992
rect 50348 33938 50404 33940
rect 50428 33938 50484 33940
rect 50508 33938 50564 33940
rect 50588 33938 50644 33940
rect 50348 32660 50404 32662
rect 50428 32660 50484 32662
rect 50508 32660 50564 32662
rect 50588 32660 50644 32662
rect 50348 32608 50374 32660
rect 50374 32608 50404 32660
rect 50428 32608 50438 32660
rect 50438 32608 50484 32660
rect 50508 32608 50554 32660
rect 50554 32608 50564 32660
rect 50588 32608 50618 32660
rect 50618 32608 50644 32660
rect 50348 32606 50404 32608
rect 50428 32606 50484 32608
rect 50508 32606 50564 32608
rect 50588 32606 50644 32608
rect 50348 31328 50404 31330
rect 50428 31328 50484 31330
rect 50508 31328 50564 31330
rect 50588 31328 50644 31330
rect 50348 31276 50374 31328
rect 50374 31276 50404 31328
rect 50428 31276 50438 31328
rect 50438 31276 50484 31328
rect 50508 31276 50554 31328
rect 50554 31276 50564 31328
rect 50588 31276 50618 31328
rect 50618 31276 50644 31328
rect 50348 31274 50404 31276
rect 50428 31274 50484 31276
rect 50508 31274 50564 31276
rect 50588 31274 50644 31276
rect 50348 29996 50404 29998
rect 50428 29996 50484 29998
rect 50508 29996 50564 29998
rect 50588 29996 50644 29998
rect 50348 29944 50374 29996
rect 50374 29944 50404 29996
rect 50428 29944 50438 29996
rect 50438 29944 50484 29996
rect 50508 29944 50554 29996
rect 50554 29944 50564 29996
rect 50588 29944 50618 29996
rect 50618 29944 50644 29996
rect 50348 29942 50404 29944
rect 50428 29942 50484 29944
rect 50508 29942 50564 29944
rect 50588 29942 50644 29944
rect 50348 28664 50404 28666
rect 50428 28664 50484 28666
rect 50508 28664 50564 28666
rect 50588 28664 50644 28666
rect 50348 28612 50374 28664
rect 50374 28612 50404 28664
rect 50428 28612 50438 28664
rect 50438 28612 50484 28664
rect 50508 28612 50554 28664
rect 50554 28612 50564 28664
rect 50588 28612 50618 28664
rect 50618 28612 50644 28664
rect 50348 28610 50404 28612
rect 50428 28610 50484 28612
rect 50508 28610 50564 28612
rect 50588 28610 50644 28612
rect 50348 27332 50404 27334
rect 50428 27332 50484 27334
rect 50508 27332 50564 27334
rect 50588 27332 50644 27334
rect 50348 27280 50374 27332
rect 50374 27280 50404 27332
rect 50428 27280 50438 27332
rect 50438 27280 50484 27332
rect 50508 27280 50554 27332
rect 50554 27280 50564 27332
rect 50588 27280 50618 27332
rect 50618 27280 50644 27332
rect 50348 27278 50404 27280
rect 50428 27278 50484 27280
rect 50508 27278 50564 27280
rect 50588 27278 50644 27280
rect 50348 26000 50404 26002
rect 50428 26000 50484 26002
rect 50508 26000 50564 26002
rect 50588 26000 50644 26002
rect 50348 25948 50374 26000
rect 50374 25948 50404 26000
rect 50428 25948 50438 26000
rect 50438 25948 50484 26000
rect 50508 25948 50554 26000
rect 50554 25948 50564 26000
rect 50588 25948 50618 26000
rect 50618 25948 50644 26000
rect 50348 25946 50404 25948
rect 50428 25946 50484 25948
rect 50508 25946 50564 25948
rect 50588 25946 50644 25948
rect 50348 24668 50404 24670
rect 50428 24668 50484 24670
rect 50508 24668 50564 24670
rect 50588 24668 50644 24670
rect 50348 24616 50374 24668
rect 50374 24616 50404 24668
rect 50428 24616 50438 24668
rect 50438 24616 50484 24668
rect 50508 24616 50554 24668
rect 50554 24616 50564 24668
rect 50588 24616 50618 24668
rect 50618 24616 50644 24668
rect 50348 24614 50404 24616
rect 50428 24614 50484 24616
rect 50508 24614 50564 24616
rect 50588 24614 50644 24616
rect 50348 23336 50404 23338
rect 50428 23336 50484 23338
rect 50508 23336 50564 23338
rect 50588 23336 50644 23338
rect 50348 23284 50374 23336
rect 50374 23284 50404 23336
rect 50428 23284 50438 23336
rect 50438 23284 50484 23336
rect 50508 23284 50554 23336
rect 50554 23284 50564 23336
rect 50588 23284 50618 23336
rect 50618 23284 50644 23336
rect 50348 23282 50404 23284
rect 50428 23282 50484 23284
rect 50508 23282 50564 23284
rect 50588 23282 50644 23284
rect 50348 22004 50404 22006
rect 50428 22004 50484 22006
rect 50508 22004 50564 22006
rect 50588 22004 50644 22006
rect 50348 21952 50374 22004
rect 50374 21952 50404 22004
rect 50428 21952 50438 22004
rect 50438 21952 50484 22004
rect 50508 21952 50554 22004
rect 50554 21952 50564 22004
rect 50588 21952 50618 22004
rect 50618 21952 50644 22004
rect 50348 21950 50404 21952
rect 50428 21950 50484 21952
rect 50508 21950 50564 21952
rect 50588 21950 50644 21952
rect 50348 20672 50404 20674
rect 50428 20672 50484 20674
rect 50508 20672 50564 20674
rect 50588 20672 50644 20674
rect 50348 20620 50374 20672
rect 50374 20620 50404 20672
rect 50428 20620 50438 20672
rect 50438 20620 50484 20672
rect 50508 20620 50554 20672
rect 50554 20620 50564 20672
rect 50588 20620 50618 20672
rect 50618 20620 50644 20672
rect 50348 20618 50404 20620
rect 50428 20618 50484 20620
rect 50508 20618 50564 20620
rect 50588 20618 50644 20620
rect 50348 19340 50404 19342
rect 50428 19340 50484 19342
rect 50508 19340 50564 19342
rect 50588 19340 50644 19342
rect 50348 19288 50374 19340
rect 50374 19288 50404 19340
rect 50428 19288 50438 19340
rect 50438 19288 50484 19340
rect 50508 19288 50554 19340
rect 50554 19288 50564 19340
rect 50588 19288 50618 19340
rect 50618 19288 50644 19340
rect 50348 19286 50404 19288
rect 50428 19286 50484 19288
rect 50508 19286 50564 19288
rect 50588 19286 50644 19288
rect 50348 18008 50404 18010
rect 50428 18008 50484 18010
rect 50508 18008 50564 18010
rect 50588 18008 50644 18010
rect 50348 17956 50374 18008
rect 50374 17956 50404 18008
rect 50428 17956 50438 18008
rect 50438 17956 50484 18008
rect 50508 17956 50554 18008
rect 50554 17956 50564 18008
rect 50588 17956 50618 18008
rect 50618 17956 50644 18008
rect 50348 17954 50404 17956
rect 50428 17954 50484 17956
rect 50508 17954 50564 17956
rect 50588 17954 50644 17956
rect 50348 16676 50404 16678
rect 50428 16676 50484 16678
rect 50508 16676 50564 16678
rect 50588 16676 50644 16678
rect 50348 16624 50374 16676
rect 50374 16624 50404 16676
rect 50428 16624 50438 16676
rect 50438 16624 50484 16676
rect 50508 16624 50554 16676
rect 50554 16624 50564 16676
rect 50588 16624 50618 16676
rect 50618 16624 50644 16676
rect 50348 16622 50404 16624
rect 50428 16622 50484 16624
rect 50508 16622 50564 16624
rect 50588 16622 50644 16624
rect 50348 15344 50404 15346
rect 50428 15344 50484 15346
rect 50508 15344 50564 15346
rect 50588 15344 50644 15346
rect 50348 15292 50374 15344
rect 50374 15292 50404 15344
rect 50428 15292 50438 15344
rect 50438 15292 50484 15344
rect 50508 15292 50554 15344
rect 50554 15292 50564 15344
rect 50588 15292 50618 15344
rect 50618 15292 50644 15344
rect 50348 15290 50404 15292
rect 50428 15290 50484 15292
rect 50508 15290 50564 15292
rect 50588 15290 50644 15292
rect 50348 14012 50404 14014
rect 50428 14012 50484 14014
rect 50508 14012 50564 14014
rect 50588 14012 50644 14014
rect 50348 13960 50374 14012
rect 50374 13960 50404 14012
rect 50428 13960 50438 14012
rect 50438 13960 50484 14012
rect 50508 13960 50554 14012
rect 50554 13960 50564 14012
rect 50588 13960 50618 14012
rect 50618 13960 50644 14012
rect 50348 13958 50404 13960
rect 50428 13958 50484 13960
rect 50508 13958 50564 13960
rect 50588 13958 50644 13960
rect 50348 12680 50404 12682
rect 50428 12680 50484 12682
rect 50508 12680 50564 12682
rect 50588 12680 50644 12682
rect 50348 12628 50374 12680
rect 50374 12628 50404 12680
rect 50428 12628 50438 12680
rect 50438 12628 50484 12680
rect 50508 12628 50554 12680
rect 50554 12628 50564 12680
rect 50588 12628 50618 12680
rect 50618 12628 50644 12680
rect 50348 12626 50404 12628
rect 50428 12626 50484 12628
rect 50508 12626 50564 12628
rect 50588 12626 50644 12628
rect 50348 11348 50404 11350
rect 50428 11348 50484 11350
rect 50508 11348 50564 11350
rect 50588 11348 50644 11350
rect 50348 11296 50374 11348
rect 50374 11296 50404 11348
rect 50428 11296 50438 11348
rect 50438 11296 50484 11348
rect 50508 11296 50554 11348
rect 50554 11296 50564 11348
rect 50588 11296 50618 11348
rect 50618 11296 50644 11348
rect 50348 11294 50404 11296
rect 50428 11294 50484 11296
rect 50508 11294 50564 11296
rect 50588 11294 50644 11296
rect 50348 10016 50404 10018
rect 50428 10016 50484 10018
rect 50508 10016 50564 10018
rect 50588 10016 50644 10018
rect 50348 9964 50374 10016
rect 50374 9964 50404 10016
rect 50428 9964 50438 10016
rect 50438 9964 50484 10016
rect 50508 9964 50554 10016
rect 50554 9964 50564 10016
rect 50588 9964 50618 10016
rect 50618 9964 50644 10016
rect 50348 9962 50404 9964
rect 50428 9962 50484 9964
rect 50508 9962 50564 9964
rect 50588 9962 50644 9964
rect 50348 8684 50404 8686
rect 50428 8684 50484 8686
rect 50508 8684 50564 8686
rect 50588 8684 50644 8686
rect 50348 8632 50374 8684
rect 50374 8632 50404 8684
rect 50428 8632 50438 8684
rect 50438 8632 50484 8684
rect 50508 8632 50554 8684
rect 50554 8632 50564 8684
rect 50588 8632 50618 8684
rect 50618 8632 50644 8684
rect 50348 8630 50404 8632
rect 50428 8630 50484 8632
rect 50508 8630 50564 8632
rect 50588 8630 50644 8632
rect 50348 7352 50404 7354
rect 50428 7352 50484 7354
rect 50508 7352 50564 7354
rect 50588 7352 50644 7354
rect 50348 7300 50374 7352
rect 50374 7300 50404 7352
rect 50428 7300 50438 7352
rect 50438 7300 50484 7352
rect 50508 7300 50554 7352
rect 50554 7300 50564 7352
rect 50588 7300 50618 7352
rect 50618 7300 50644 7352
rect 50348 7298 50404 7300
rect 50428 7298 50484 7300
rect 50508 7298 50564 7300
rect 50588 7298 50644 7300
rect 50348 6020 50404 6022
rect 50428 6020 50484 6022
rect 50508 6020 50564 6022
rect 50588 6020 50644 6022
rect 50348 5968 50374 6020
rect 50374 5968 50404 6020
rect 50428 5968 50438 6020
rect 50438 5968 50484 6020
rect 50508 5968 50554 6020
rect 50554 5968 50564 6020
rect 50588 5968 50618 6020
rect 50618 5968 50644 6020
rect 50348 5966 50404 5968
rect 50428 5966 50484 5968
rect 50508 5966 50564 5968
rect 50588 5966 50644 5968
rect 50348 4688 50404 4690
rect 50428 4688 50484 4690
rect 50508 4688 50564 4690
rect 50588 4688 50644 4690
rect 50348 4636 50374 4688
rect 50374 4636 50404 4688
rect 50428 4636 50438 4688
rect 50438 4636 50484 4688
rect 50508 4636 50554 4688
rect 50554 4636 50564 4688
rect 50588 4636 50618 4688
rect 50618 4636 50644 4688
rect 50348 4634 50404 4636
rect 50428 4634 50484 4636
rect 50508 4634 50564 4636
rect 50588 4634 50644 4636
rect 50348 3356 50404 3358
rect 50428 3356 50484 3358
rect 50508 3356 50564 3358
rect 50588 3356 50644 3358
rect 50348 3304 50374 3356
rect 50374 3304 50404 3356
rect 50428 3304 50438 3356
rect 50438 3304 50484 3356
rect 50508 3304 50554 3356
rect 50554 3304 50564 3356
rect 50588 3304 50618 3356
rect 50618 3304 50644 3356
rect 50348 3302 50404 3304
rect 50428 3302 50484 3304
rect 50508 3302 50564 3304
rect 50588 3302 50644 3304
<< metal3 >>
rect 4256 57308 4576 57309
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 57243 4576 57244
rect 34976 57308 35296 57309
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 57243 35296 57244
rect 19616 56642 19936 56643
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 56577 19936 56578
rect 50336 56642 50656 56643
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 56577 50656 56578
rect 4256 55976 4576 55977
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 55911 4576 55912
rect 34976 55976 35296 55977
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 55911 35296 55912
rect 19616 55310 19936 55311
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 55245 19936 55246
rect 50336 55310 50656 55311
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 55245 50656 55246
rect 4256 54644 4576 54645
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 54579 4576 54580
rect 34976 54644 35296 54645
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 54579 35296 54580
rect 19616 53978 19936 53979
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 53913 19936 53914
rect 50336 53978 50656 53979
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 53913 50656 53914
rect 4256 53312 4576 53313
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 53247 4576 53248
rect 34976 53312 35296 53313
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 53247 35296 53248
rect 19616 52646 19936 52647
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 52581 19936 52582
rect 50336 52646 50656 52647
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 52581 50656 52582
rect 4256 51980 4576 51981
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 51915 4576 51916
rect 34976 51980 35296 51981
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 51915 35296 51916
rect 19616 51314 19936 51315
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 51249 19936 51250
rect 50336 51314 50656 51315
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 51249 50656 51250
rect 4256 50648 4576 50649
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 50583 4576 50584
rect 34976 50648 35296 50649
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 50583 35296 50584
rect 19616 49982 19936 49983
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 49917 19936 49918
rect 50336 49982 50656 49983
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 49917 50656 49918
rect 4256 49316 4576 49317
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 49251 4576 49252
rect 34976 49316 35296 49317
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 49251 35296 49252
rect 19616 48650 19936 48651
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 48585 19936 48586
rect 50336 48650 50656 48651
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 48585 50656 48586
rect 4256 47984 4576 47985
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 47919 4576 47920
rect 34976 47984 35296 47985
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 47919 35296 47920
rect 19616 47318 19936 47319
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 47253 19936 47254
rect 50336 47318 50656 47319
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 47253 50656 47254
rect 4256 46652 4576 46653
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 46587 4576 46588
rect 34976 46652 35296 46653
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 46587 35296 46588
rect 19616 45986 19936 45987
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 45921 19936 45922
rect 50336 45986 50656 45987
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 45921 50656 45922
rect 4256 45320 4576 45321
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 45255 4576 45256
rect 34976 45320 35296 45321
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 45255 35296 45256
rect 19616 44654 19936 44655
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 44589 19936 44590
rect 50336 44654 50656 44655
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 44589 50656 44590
rect 4256 43988 4576 43989
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 43923 4576 43924
rect 34976 43988 35296 43989
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 43923 35296 43924
rect 19616 43322 19936 43323
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 43257 19936 43258
rect 50336 43322 50656 43323
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 43257 50656 43258
rect 4256 42656 4576 42657
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 42591 4576 42592
rect 34976 42656 35296 42657
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 42591 35296 42592
rect 19616 41990 19936 41991
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 41925 19936 41926
rect 50336 41990 50656 41991
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 41925 50656 41926
rect 4256 41324 4576 41325
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 41259 4576 41260
rect 34976 41324 35296 41325
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 41259 35296 41260
rect 19616 40658 19936 40659
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 40593 19936 40594
rect 50336 40658 50656 40659
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 40593 50656 40594
rect 4256 39992 4576 39993
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 39927 4576 39928
rect 34976 39992 35296 39993
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 39927 35296 39928
rect 19616 39326 19936 39327
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 39261 19936 39262
rect 50336 39326 50656 39327
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 39261 50656 39262
rect 4256 38660 4576 38661
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 38595 4576 38596
rect 34976 38660 35296 38661
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 38595 35296 38596
rect 19616 37994 19936 37995
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 37929 19936 37930
rect 50336 37994 50656 37995
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 37929 50656 37930
rect 4256 37328 4576 37329
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 37263 4576 37264
rect 34976 37328 35296 37329
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 37263 35296 37264
rect 19616 36662 19936 36663
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 36597 19936 36598
rect 50336 36662 50656 36663
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 36597 50656 36598
rect 4256 35996 4576 35997
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 35931 4576 35932
rect 34976 35996 35296 35997
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 35931 35296 35932
rect 19616 35330 19936 35331
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 35265 19936 35266
rect 50336 35330 50656 35331
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 35265 50656 35266
rect 4256 34664 4576 34665
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 34599 4576 34600
rect 34976 34664 35296 34665
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 34599 35296 34600
rect 19616 33998 19936 33999
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 33933 19936 33934
rect 50336 33998 50656 33999
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 33933 50656 33934
rect 4256 33332 4576 33333
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 33267 4576 33268
rect 34976 33332 35296 33333
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 33267 35296 33268
rect 19616 32666 19936 32667
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 32601 19936 32602
rect 50336 32666 50656 32667
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 32601 50656 32602
rect 4256 32000 4576 32001
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 31935 4576 31936
rect 34976 32000 35296 32001
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 31935 35296 31936
rect 19616 31334 19936 31335
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 31269 19936 31270
rect 50336 31334 50656 31335
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 31269 50656 31270
rect 4256 30668 4576 30669
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 30603 4576 30604
rect 34976 30668 35296 30669
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 30603 35296 30604
rect 19616 30002 19936 30003
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 29937 19936 29938
rect 50336 30002 50656 30003
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 29937 50656 29938
rect 4256 29336 4576 29337
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 29271 4576 29272
rect 34976 29336 35296 29337
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 29271 35296 29272
rect 19616 28670 19936 28671
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 28605 19936 28606
rect 50336 28670 50656 28671
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 28605 50656 28606
rect 4256 28004 4576 28005
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 27939 4576 27940
rect 34976 28004 35296 28005
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 27939 35296 27940
rect 19616 27338 19936 27339
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 27273 19936 27274
rect 50336 27338 50656 27339
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 27273 50656 27274
rect 4256 26672 4576 26673
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 26607 4576 26608
rect 34976 26672 35296 26673
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 26607 35296 26608
rect 19616 26006 19936 26007
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 25941 19936 25942
rect 50336 26006 50656 26007
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 25941 50656 25942
rect 4256 25340 4576 25341
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 25275 4576 25276
rect 34976 25340 35296 25341
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 25275 35296 25276
rect 19616 24674 19936 24675
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 24609 19936 24610
rect 50336 24674 50656 24675
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 24609 50656 24610
rect 4256 24008 4576 24009
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 23943 4576 23944
rect 34976 24008 35296 24009
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 23943 35296 23944
rect 19616 23342 19936 23343
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 23277 19936 23278
rect 50336 23342 50656 23343
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 23277 50656 23278
rect 4256 22676 4576 22677
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 22611 4576 22612
rect 34976 22676 35296 22677
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 22611 35296 22612
rect 19616 22010 19936 22011
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 21945 19936 21946
rect 50336 22010 50656 22011
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 21945 50656 21946
rect 4256 21344 4576 21345
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 21279 4576 21280
rect 34976 21344 35296 21345
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 21279 35296 21280
rect 19616 20678 19936 20679
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 20613 19936 20614
rect 50336 20678 50656 20679
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 20613 50656 20614
rect 4256 20012 4576 20013
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 19947 4576 19948
rect 34976 20012 35296 20013
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 19947 35296 19948
rect 19616 19346 19936 19347
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 19281 19936 19282
rect 50336 19346 50656 19347
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 19281 50656 19282
rect 4256 18680 4576 18681
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 18615 4576 18616
rect 34976 18680 35296 18681
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 18615 35296 18616
rect 19616 18014 19936 18015
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 17949 19936 17950
rect 50336 18014 50656 18015
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 17949 50656 17950
rect 4256 17348 4576 17349
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 17283 4576 17284
rect 34976 17348 35296 17349
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 17283 35296 17284
rect 19616 16682 19936 16683
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 16617 19936 16618
rect 50336 16682 50656 16683
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 16617 50656 16618
rect 4256 16016 4576 16017
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 15951 4576 15952
rect 34976 16016 35296 16017
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 15951 35296 15952
rect 19616 15350 19936 15351
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 15285 19936 15286
rect 50336 15350 50656 15351
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 15285 50656 15286
rect 4256 14684 4576 14685
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 14619 4576 14620
rect 34976 14684 35296 14685
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 14619 35296 14620
rect 19616 14018 19936 14019
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 13953 19936 13954
rect 50336 14018 50656 14019
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 13953 50656 13954
rect 4256 13352 4576 13353
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 13287 4576 13288
rect 34976 13352 35296 13353
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 13287 35296 13288
rect 19616 12686 19936 12687
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 12621 19936 12622
rect 50336 12686 50656 12687
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 12621 50656 12622
rect 4256 12020 4576 12021
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 11955 4576 11956
rect 34976 12020 35296 12021
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 11955 35296 11956
rect 19616 11354 19936 11355
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 11289 19936 11290
rect 50336 11354 50656 11355
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 11289 50656 11290
rect 4256 10688 4576 10689
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 10623 4576 10624
rect 34976 10688 35296 10689
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 10623 35296 10624
rect 19616 10022 19936 10023
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 9957 19936 9958
rect 50336 10022 50656 10023
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 9957 50656 9958
rect 4256 9356 4576 9357
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 9291 4576 9292
rect 34976 9356 35296 9357
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 9291 35296 9292
rect 19616 8690 19936 8691
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 8625 19936 8626
rect 50336 8690 50656 8691
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 8625 50656 8626
rect 4256 8024 4576 8025
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 7959 4576 7960
rect 34976 8024 35296 8025
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 7959 35296 7960
rect 19616 7358 19936 7359
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 7293 19936 7294
rect 50336 7358 50656 7359
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 7293 50656 7294
rect 4256 6692 4576 6693
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 6627 4576 6628
rect 34976 6692 35296 6693
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 6627 35296 6628
rect 19616 6026 19936 6027
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 5961 19936 5962
rect 50336 6026 50656 6027
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 5961 50656 5962
rect 4256 5360 4576 5361
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 5295 4576 5296
rect 34976 5360 35296 5361
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 5295 35296 5296
rect 19616 4694 19936 4695
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 4629 19936 4630
rect 50336 4694 50656 4695
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 4629 50656 4630
rect 4256 4028 4576 4029
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 3963 4576 3964
rect 34976 4028 35296 4029
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 3963 35296 3964
rect 33519 3804 33585 3807
rect 33519 3802 33726 3804
rect 33519 3746 33524 3802
rect 33580 3746 33726 3802
rect 33519 3744 33726 3746
rect 33519 3741 33585 3744
rect 19887 3508 19953 3511
rect 19887 3506 20094 3508
rect 19887 3450 19892 3506
rect 19948 3450 20094 3506
rect 19887 3448 20094 3450
rect 19887 3445 19953 3448
rect 19616 3362 19936 3363
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 19616 3297 19936 3298
rect 19791 3212 19857 3215
rect 20034 3212 20094 3448
rect 33666 3363 33726 3744
rect 33666 3358 33777 3363
rect 33666 3302 33716 3358
rect 33772 3302 33777 3358
rect 33666 3300 33777 3302
rect 33711 3297 33777 3300
rect 50336 3362 50656 3363
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 50336 3297 50656 3298
rect 44271 3212 44337 3215
rect 19791 3210 20094 3212
rect 19791 3154 19796 3210
rect 19852 3154 20094 3210
rect 19791 3152 20094 3154
rect 44226 3210 44337 3212
rect 44226 3154 44276 3210
rect 44332 3154 44337 3210
rect 19791 3149 19857 3152
rect 44226 3149 44337 3154
rect 35631 3064 35697 3067
rect 35394 3062 35697 3064
rect 35394 3006 35636 3062
rect 35692 3006 35697 3062
rect 35394 3004 35697 3006
rect 4256 2696 4576 2697
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4256 2631 4576 2632
rect 34976 2696 35296 2697
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 34976 2631 35296 2632
rect 35394 2472 35454 3004
rect 35631 3001 35697 3004
rect 44226 2919 44286 3149
rect 44226 2914 44337 2919
rect 44226 2858 44276 2914
rect 44332 2858 44337 2914
rect 44226 2856 44337 2858
rect 44271 2853 44337 2856
rect 35535 2472 35601 2475
rect 35394 2470 35601 2472
rect 35394 2414 35540 2470
rect 35596 2414 35601 2470
rect 35394 2412 35601 2414
rect 35535 2409 35601 2412
<< via3 >>
rect 4264 57304 4328 57308
rect 4264 57248 4268 57304
rect 4268 57248 4324 57304
rect 4324 57248 4328 57304
rect 4264 57244 4328 57248
rect 4344 57304 4408 57308
rect 4344 57248 4348 57304
rect 4348 57248 4404 57304
rect 4404 57248 4408 57304
rect 4344 57244 4408 57248
rect 4424 57304 4488 57308
rect 4424 57248 4428 57304
rect 4428 57248 4484 57304
rect 4484 57248 4488 57304
rect 4424 57244 4488 57248
rect 4504 57304 4568 57308
rect 4504 57248 4508 57304
rect 4508 57248 4564 57304
rect 4564 57248 4568 57304
rect 4504 57244 4568 57248
rect 34984 57304 35048 57308
rect 34984 57248 34988 57304
rect 34988 57248 35044 57304
rect 35044 57248 35048 57304
rect 34984 57244 35048 57248
rect 35064 57304 35128 57308
rect 35064 57248 35068 57304
rect 35068 57248 35124 57304
rect 35124 57248 35128 57304
rect 35064 57244 35128 57248
rect 35144 57304 35208 57308
rect 35144 57248 35148 57304
rect 35148 57248 35204 57304
rect 35204 57248 35208 57304
rect 35144 57244 35208 57248
rect 35224 57304 35288 57308
rect 35224 57248 35228 57304
rect 35228 57248 35284 57304
rect 35284 57248 35288 57304
rect 35224 57244 35288 57248
rect 19624 56638 19688 56642
rect 19624 56582 19628 56638
rect 19628 56582 19684 56638
rect 19684 56582 19688 56638
rect 19624 56578 19688 56582
rect 19704 56638 19768 56642
rect 19704 56582 19708 56638
rect 19708 56582 19764 56638
rect 19764 56582 19768 56638
rect 19704 56578 19768 56582
rect 19784 56638 19848 56642
rect 19784 56582 19788 56638
rect 19788 56582 19844 56638
rect 19844 56582 19848 56638
rect 19784 56578 19848 56582
rect 19864 56638 19928 56642
rect 19864 56582 19868 56638
rect 19868 56582 19924 56638
rect 19924 56582 19928 56638
rect 19864 56578 19928 56582
rect 50344 56638 50408 56642
rect 50344 56582 50348 56638
rect 50348 56582 50404 56638
rect 50404 56582 50408 56638
rect 50344 56578 50408 56582
rect 50424 56638 50488 56642
rect 50424 56582 50428 56638
rect 50428 56582 50484 56638
rect 50484 56582 50488 56638
rect 50424 56578 50488 56582
rect 50504 56638 50568 56642
rect 50504 56582 50508 56638
rect 50508 56582 50564 56638
rect 50564 56582 50568 56638
rect 50504 56578 50568 56582
rect 50584 56638 50648 56642
rect 50584 56582 50588 56638
rect 50588 56582 50644 56638
rect 50644 56582 50648 56638
rect 50584 56578 50648 56582
rect 4264 55972 4328 55976
rect 4264 55916 4268 55972
rect 4268 55916 4324 55972
rect 4324 55916 4328 55972
rect 4264 55912 4328 55916
rect 4344 55972 4408 55976
rect 4344 55916 4348 55972
rect 4348 55916 4404 55972
rect 4404 55916 4408 55972
rect 4344 55912 4408 55916
rect 4424 55972 4488 55976
rect 4424 55916 4428 55972
rect 4428 55916 4484 55972
rect 4484 55916 4488 55972
rect 4424 55912 4488 55916
rect 4504 55972 4568 55976
rect 4504 55916 4508 55972
rect 4508 55916 4564 55972
rect 4564 55916 4568 55972
rect 4504 55912 4568 55916
rect 34984 55972 35048 55976
rect 34984 55916 34988 55972
rect 34988 55916 35044 55972
rect 35044 55916 35048 55972
rect 34984 55912 35048 55916
rect 35064 55972 35128 55976
rect 35064 55916 35068 55972
rect 35068 55916 35124 55972
rect 35124 55916 35128 55972
rect 35064 55912 35128 55916
rect 35144 55972 35208 55976
rect 35144 55916 35148 55972
rect 35148 55916 35204 55972
rect 35204 55916 35208 55972
rect 35144 55912 35208 55916
rect 35224 55972 35288 55976
rect 35224 55916 35228 55972
rect 35228 55916 35284 55972
rect 35284 55916 35288 55972
rect 35224 55912 35288 55916
rect 19624 55306 19688 55310
rect 19624 55250 19628 55306
rect 19628 55250 19684 55306
rect 19684 55250 19688 55306
rect 19624 55246 19688 55250
rect 19704 55306 19768 55310
rect 19704 55250 19708 55306
rect 19708 55250 19764 55306
rect 19764 55250 19768 55306
rect 19704 55246 19768 55250
rect 19784 55306 19848 55310
rect 19784 55250 19788 55306
rect 19788 55250 19844 55306
rect 19844 55250 19848 55306
rect 19784 55246 19848 55250
rect 19864 55306 19928 55310
rect 19864 55250 19868 55306
rect 19868 55250 19924 55306
rect 19924 55250 19928 55306
rect 19864 55246 19928 55250
rect 50344 55306 50408 55310
rect 50344 55250 50348 55306
rect 50348 55250 50404 55306
rect 50404 55250 50408 55306
rect 50344 55246 50408 55250
rect 50424 55306 50488 55310
rect 50424 55250 50428 55306
rect 50428 55250 50484 55306
rect 50484 55250 50488 55306
rect 50424 55246 50488 55250
rect 50504 55306 50568 55310
rect 50504 55250 50508 55306
rect 50508 55250 50564 55306
rect 50564 55250 50568 55306
rect 50504 55246 50568 55250
rect 50584 55306 50648 55310
rect 50584 55250 50588 55306
rect 50588 55250 50644 55306
rect 50644 55250 50648 55306
rect 50584 55246 50648 55250
rect 4264 54640 4328 54644
rect 4264 54584 4268 54640
rect 4268 54584 4324 54640
rect 4324 54584 4328 54640
rect 4264 54580 4328 54584
rect 4344 54640 4408 54644
rect 4344 54584 4348 54640
rect 4348 54584 4404 54640
rect 4404 54584 4408 54640
rect 4344 54580 4408 54584
rect 4424 54640 4488 54644
rect 4424 54584 4428 54640
rect 4428 54584 4484 54640
rect 4484 54584 4488 54640
rect 4424 54580 4488 54584
rect 4504 54640 4568 54644
rect 4504 54584 4508 54640
rect 4508 54584 4564 54640
rect 4564 54584 4568 54640
rect 4504 54580 4568 54584
rect 34984 54640 35048 54644
rect 34984 54584 34988 54640
rect 34988 54584 35044 54640
rect 35044 54584 35048 54640
rect 34984 54580 35048 54584
rect 35064 54640 35128 54644
rect 35064 54584 35068 54640
rect 35068 54584 35124 54640
rect 35124 54584 35128 54640
rect 35064 54580 35128 54584
rect 35144 54640 35208 54644
rect 35144 54584 35148 54640
rect 35148 54584 35204 54640
rect 35204 54584 35208 54640
rect 35144 54580 35208 54584
rect 35224 54640 35288 54644
rect 35224 54584 35228 54640
rect 35228 54584 35284 54640
rect 35284 54584 35288 54640
rect 35224 54580 35288 54584
rect 19624 53974 19688 53978
rect 19624 53918 19628 53974
rect 19628 53918 19684 53974
rect 19684 53918 19688 53974
rect 19624 53914 19688 53918
rect 19704 53974 19768 53978
rect 19704 53918 19708 53974
rect 19708 53918 19764 53974
rect 19764 53918 19768 53974
rect 19704 53914 19768 53918
rect 19784 53974 19848 53978
rect 19784 53918 19788 53974
rect 19788 53918 19844 53974
rect 19844 53918 19848 53974
rect 19784 53914 19848 53918
rect 19864 53974 19928 53978
rect 19864 53918 19868 53974
rect 19868 53918 19924 53974
rect 19924 53918 19928 53974
rect 19864 53914 19928 53918
rect 50344 53974 50408 53978
rect 50344 53918 50348 53974
rect 50348 53918 50404 53974
rect 50404 53918 50408 53974
rect 50344 53914 50408 53918
rect 50424 53974 50488 53978
rect 50424 53918 50428 53974
rect 50428 53918 50484 53974
rect 50484 53918 50488 53974
rect 50424 53914 50488 53918
rect 50504 53974 50568 53978
rect 50504 53918 50508 53974
rect 50508 53918 50564 53974
rect 50564 53918 50568 53974
rect 50504 53914 50568 53918
rect 50584 53974 50648 53978
rect 50584 53918 50588 53974
rect 50588 53918 50644 53974
rect 50644 53918 50648 53974
rect 50584 53914 50648 53918
rect 4264 53308 4328 53312
rect 4264 53252 4268 53308
rect 4268 53252 4324 53308
rect 4324 53252 4328 53308
rect 4264 53248 4328 53252
rect 4344 53308 4408 53312
rect 4344 53252 4348 53308
rect 4348 53252 4404 53308
rect 4404 53252 4408 53308
rect 4344 53248 4408 53252
rect 4424 53308 4488 53312
rect 4424 53252 4428 53308
rect 4428 53252 4484 53308
rect 4484 53252 4488 53308
rect 4424 53248 4488 53252
rect 4504 53308 4568 53312
rect 4504 53252 4508 53308
rect 4508 53252 4564 53308
rect 4564 53252 4568 53308
rect 4504 53248 4568 53252
rect 34984 53308 35048 53312
rect 34984 53252 34988 53308
rect 34988 53252 35044 53308
rect 35044 53252 35048 53308
rect 34984 53248 35048 53252
rect 35064 53308 35128 53312
rect 35064 53252 35068 53308
rect 35068 53252 35124 53308
rect 35124 53252 35128 53308
rect 35064 53248 35128 53252
rect 35144 53308 35208 53312
rect 35144 53252 35148 53308
rect 35148 53252 35204 53308
rect 35204 53252 35208 53308
rect 35144 53248 35208 53252
rect 35224 53308 35288 53312
rect 35224 53252 35228 53308
rect 35228 53252 35284 53308
rect 35284 53252 35288 53308
rect 35224 53248 35288 53252
rect 19624 52642 19688 52646
rect 19624 52586 19628 52642
rect 19628 52586 19684 52642
rect 19684 52586 19688 52642
rect 19624 52582 19688 52586
rect 19704 52642 19768 52646
rect 19704 52586 19708 52642
rect 19708 52586 19764 52642
rect 19764 52586 19768 52642
rect 19704 52582 19768 52586
rect 19784 52642 19848 52646
rect 19784 52586 19788 52642
rect 19788 52586 19844 52642
rect 19844 52586 19848 52642
rect 19784 52582 19848 52586
rect 19864 52642 19928 52646
rect 19864 52586 19868 52642
rect 19868 52586 19924 52642
rect 19924 52586 19928 52642
rect 19864 52582 19928 52586
rect 50344 52642 50408 52646
rect 50344 52586 50348 52642
rect 50348 52586 50404 52642
rect 50404 52586 50408 52642
rect 50344 52582 50408 52586
rect 50424 52642 50488 52646
rect 50424 52586 50428 52642
rect 50428 52586 50484 52642
rect 50484 52586 50488 52642
rect 50424 52582 50488 52586
rect 50504 52642 50568 52646
rect 50504 52586 50508 52642
rect 50508 52586 50564 52642
rect 50564 52586 50568 52642
rect 50504 52582 50568 52586
rect 50584 52642 50648 52646
rect 50584 52586 50588 52642
rect 50588 52586 50644 52642
rect 50644 52586 50648 52642
rect 50584 52582 50648 52586
rect 4264 51976 4328 51980
rect 4264 51920 4268 51976
rect 4268 51920 4324 51976
rect 4324 51920 4328 51976
rect 4264 51916 4328 51920
rect 4344 51976 4408 51980
rect 4344 51920 4348 51976
rect 4348 51920 4404 51976
rect 4404 51920 4408 51976
rect 4344 51916 4408 51920
rect 4424 51976 4488 51980
rect 4424 51920 4428 51976
rect 4428 51920 4484 51976
rect 4484 51920 4488 51976
rect 4424 51916 4488 51920
rect 4504 51976 4568 51980
rect 4504 51920 4508 51976
rect 4508 51920 4564 51976
rect 4564 51920 4568 51976
rect 4504 51916 4568 51920
rect 34984 51976 35048 51980
rect 34984 51920 34988 51976
rect 34988 51920 35044 51976
rect 35044 51920 35048 51976
rect 34984 51916 35048 51920
rect 35064 51976 35128 51980
rect 35064 51920 35068 51976
rect 35068 51920 35124 51976
rect 35124 51920 35128 51976
rect 35064 51916 35128 51920
rect 35144 51976 35208 51980
rect 35144 51920 35148 51976
rect 35148 51920 35204 51976
rect 35204 51920 35208 51976
rect 35144 51916 35208 51920
rect 35224 51976 35288 51980
rect 35224 51920 35228 51976
rect 35228 51920 35284 51976
rect 35284 51920 35288 51976
rect 35224 51916 35288 51920
rect 19624 51310 19688 51314
rect 19624 51254 19628 51310
rect 19628 51254 19684 51310
rect 19684 51254 19688 51310
rect 19624 51250 19688 51254
rect 19704 51310 19768 51314
rect 19704 51254 19708 51310
rect 19708 51254 19764 51310
rect 19764 51254 19768 51310
rect 19704 51250 19768 51254
rect 19784 51310 19848 51314
rect 19784 51254 19788 51310
rect 19788 51254 19844 51310
rect 19844 51254 19848 51310
rect 19784 51250 19848 51254
rect 19864 51310 19928 51314
rect 19864 51254 19868 51310
rect 19868 51254 19924 51310
rect 19924 51254 19928 51310
rect 19864 51250 19928 51254
rect 50344 51310 50408 51314
rect 50344 51254 50348 51310
rect 50348 51254 50404 51310
rect 50404 51254 50408 51310
rect 50344 51250 50408 51254
rect 50424 51310 50488 51314
rect 50424 51254 50428 51310
rect 50428 51254 50484 51310
rect 50484 51254 50488 51310
rect 50424 51250 50488 51254
rect 50504 51310 50568 51314
rect 50504 51254 50508 51310
rect 50508 51254 50564 51310
rect 50564 51254 50568 51310
rect 50504 51250 50568 51254
rect 50584 51310 50648 51314
rect 50584 51254 50588 51310
rect 50588 51254 50644 51310
rect 50644 51254 50648 51310
rect 50584 51250 50648 51254
rect 4264 50644 4328 50648
rect 4264 50588 4268 50644
rect 4268 50588 4324 50644
rect 4324 50588 4328 50644
rect 4264 50584 4328 50588
rect 4344 50644 4408 50648
rect 4344 50588 4348 50644
rect 4348 50588 4404 50644
rect 4404 50588 4408 50644
rect 4344 50584 4408 50588
rect 4424 50644 4488 50648
rect 4424 50588 4428 50644
rect 4428 50588 4484 50644
rect 4484 50588 4488 50644
rect 4424 50584 4488 50588
rect 4504 50644 4568 50648
rect 4504 50588 4508 50644
rect 4508 50588 4564 50644
rect 4564 50588 4568 50644
rect 4504 50584 4568 50588
rect 34984 50644 35048 50648
rect 34984 50588 34988 50644
rect 34988 50588 35044 50644
rect 35044 50588 35048 50644
rect 34984 50584 35048 50588
rect 35064 50644 35128 50648
rect 35064 50588 35068 50644
rect 35068 50588 35124 50644
rect 35124 50588 35128 50644
rect 35064 50584 35128 50588
rect 35144 50644 35208 50648
rect 35144 50588 35148 50644
rect 35148 50588 35204 50644
rect 35204 50588 35208 50644
rect 35144 50584 35208 50588
rect 35224 50644 35288 50648
rect 35224 50588 35228 50644
rect 35228 50588 35284 50644
rect 35284 50588 35288 50644
rect 35224 50584 35288 50588
rect 19624 49978 19688 49982
rect 19624 49922 19628 49978
rect 19628 49922 19684 49978
rect 19684 49922 19688 49978
rect 19624 49918 19688 49922
rect 19704 49978 19768 49982
rect 19704 49922 19708 49978
rect 19708 49922 19764 49978
rect 19764 49922 19768 49978
rect 19704 49918 19768 49922
rect 19784 49978 19848 49982
rect 19784 49922 19788 49978
rect 19788 49922 19844 49978
rect 19844 49922 19848 49978
rect 19784 49918 19848 49922
rect 19864 49978 19928 49982
rect 19864 49922 19868 49978
rect 19868 49922 19924 49978
rect 19924 49922 19928 49978
rect 19864 49918 19928 49922
rect 50344 49978 50408 49982
rect 50344 49922 50348 49978
rect 50348 49922 50404 49978
rect 50404 49922 50408 49978
rect 50344 49918 50408 49922
rect 50424 49978 50488 49982
rect 50424 49922 50428 49978
rect 50428 49922 50484 49978
rect 50484 49922 50488 49978
rect 50424 49918 50488 49922
rect 50504 49978 50568 49982
rect 50504 49922 50508 49978
rect 50508 49922 50564 49978
rect 50564 49922 50568 49978
rect 50504 49918 50568 49922
rect 50584 49978 50648 49982
rect 50584 49922 50588 49978
rect 50588 49922 50644 49978
rect 50644 49922 50648 49978
rect 50584 49918 50648 49922
rect 4264 49312 4328 49316
rect 4264 49256 4268 49312
rect 4268 49256 4324 49312
rect 4324 49256 4328 49312
rect 4264 49252 4328 49256
rect 4344 49312 4408 49316
rect 4344 49256 4348 49312
rect 4348 49256 4404 49312
rect 4404 49256 4408 49312
rect 4344 49252 4408 49256
rect 4424 49312 4488 49316
rect 4424 49256 4428 49312
rect 4428 49256 4484 49312
rect 4484 49256 4488 49312
rect 4424 49252 4488 49256
rect 4504 49312 4568 49316
rect 4504 49256 4508 49312
rect 4508 49256 4564 49312
rect 4564 49256 4568 49312
rect 4504 49252 4568 49256
rect 34984 49312 35048 49316
rect 34984 49256 34988 49312
rect 34988 49256 35044 49312
rect 35044 49256 35048 49312
rect 34984 49252 35048 49256
rect 35064 49312 35128 49316
rect 35064 49256 35068 49312
rect 35068 49256 35124 49312
rect 35124 49256 35128 49312
rect 35064 49252 35128 49256
rect 35144 49312 35208 49316
rect 35144 49256 35148 49312
rect 35148 49256 35204 49312
rect 35204 49256 35208 49312
rect 35144 49252 35208 49256
rect 35224 49312 35288 49316
rect 35224 49256 35228 49312
rect 35228 49256 35284 49312
rect 35284 49256 35288 49312
rect 35224 49252 35288 49256
rect 19624 48646 19688 48650
rect 19624 48590 19628 48646
rect 19628 48590 19684 48646
rect 19684 48590 19688 48646
rect 19624 48586 19688 48590
rect 19704 48646 19768 48650
rect 19704 48590 19708 48646
rect 19708 48590 19764 48646
rect 19764 48590 19768 48646
rect 19704 48586 19768 48590
rect 19784 48646 19848 48650
rect 19784 48590 19788 48646
rect 19788 48590 19844 48646
rect 19844 48590 19848 48646
rect 19784 48586 19848 48590
rect 19864 48646 19928 48650
rect 19864 48590 19868 48646
rect 19868 48590 19924 48646
rect 19924 48590 19928 48646
rect 19864 48586 19928 48590
rect 50344 48646 50408 48650
rect 50344 48590 50348 48646
rect 50348 48590 50404 48646
rect 50404 48590 50408 48646
rect 50344 48586 50408 48590
rect 50424 48646 50488 48650
rect 50424 48590 50428 48646
rect 50428 48590 50484 48646
rect 50484 48590 50488 48646
rect 50424 48586 50488 48590
rect 50504 48646 50568 48650
rect 50504 48590 50508 48646
rect 50508 48590 50564 48646
rect 50564 48590 50568 48646
rect 50504 48586 50568 48590
rect 50584 48646 50648 48650
rect 50584 48590 50588 48646
rect 50588 48590 50644 48646
rect 50644 48590 50648 48646
rect 50584 48586 50648 48590
rect 4264 47980 4328 47984
rect 4264 47924 4268 47980
rect 4268 47924 4324 47980
rect 4324 47924 4328 47980
rect 4264 47920 4328 47924
rect 4344 47980 4408 47984
rect 4344 47924 4348 47980
rect 4348 47924 4404 47980
rect 4404 47924 4408 47980
rect 4344 47920 4408 47924
rect 4424 47980 4488 47984
rect 4424 47924 4428 47980
rect 4428 47924 4484 47980
rect 4484 47924 4488 47980
rect 4424 47920 4488 47924
rect 4504 47980 4568 47984
rect 4504 47924 4508 47980
rect 4508 47924 4564 47980
rect 4564 47924 4568 47980
rect 4504 47920 4568 47924
rect 34984 47980 35048 47984
rect 34984 47924 34988 47980
rect 34988 47924 35044 47980
rect 35044 47924 35048 47980
rect 34984 47920 35048 47924
rect 35064 47980 35128 47984
rect 35064 47924 35068 47980
rect 35068 47924 35124 47980
rect 35124 47924 35128 47980
rect 35064 47920 35128 47924
rect 35144 47980 35208 47984
rect 35144 47924 35148 47980
rect 35148 47924 35204 47980
rect 35204 47924 35208 47980
rect 35144 47920 35208 47924
rect 35224 47980 35288 47984
rect 35224 47924 35228 47980
rect 35228 47924 35284 47980
rect 35284 47924 35288 47980
rect 35224 47920 35288 47924
rect 19624 47314 19688 47318
rect 19624 47258 19628 47314
rect 19628 47258 19684 47314
rect 19684 47258 19688 47314
rect 19624 47254 19688 47258
rect 19704 47314 19768 47318
rect 19704 47258 19708 47314
rect 19708 47258 19764 47314
rect 19764 47258 19768 47314
rect 19704 47254 19768 47258
rect 19784 47314 19848 47318
rect 19784 47258 19788 47314
rect 19788 47258 19844 47314
rect 19844 47258 19848 47314
rect 19784 47254 19848 47258
rect 19864 47314 19928 47318
rect 19864 47258 19868 47314
rect 19868 47258 19924 47314
rect 19924 47258 19928 47314
rect 19864 47254 19928 47258
rect 50344 47314 50408 47318
rect 50344 47258 50348 47314
rect 50348 47258 50404 47314
rect 50404 47258 50408 47314
rect 50344 47254 50408 47258
rect 50424 47314 50488 47318
rect 50424 47258 50428 47314
rect 50428 47258 50484 47314
rect 50484 47258 50488 47314
rect 50424 47254 50488 47258
rect 50504 47314 50568 47318
rect 50504 47258 50508 47314
rect 50508 47258 50564 47314
rect 50564 47258 50568 47314
rect 50504 47254 50568 47258
rect 50584 47314 50648 47318
rect 50584 47258 50588 47314
rect 50588 47258 50644 47314
rect 50644 47258 50648 47314
rect 50584 47254 50648 47258
rect 4264 46648 4328 46652
rect 4264 46592 4268 46648
rect 4268 46592 4324 46648
rect 4324 46592 4328 46648
rect 4264 46588 4328 46592
rect 4344 46648 4408 46652
rect 4344 46592 4348 46648
rect 4348 46592 4404 46648
rect 4404 46592 4408 46648
rect 4344 46588 4408 46592
rect 4424 46648 4488 46652
rect 4424 46592 4428 46648
rect 4428 46592 4484 46648
rect 4484 46592 4488 46648
rect 4424 46588 4488 46592
rect 4504 46648 4568 46652
rect 4504 46592 4508 46648
rect 4508 46592 4564 46648
rect 4564 46592 4568 46648
rect 4504 46588 4568 46592
rect 34984 46648 35048 46652
rect 34984 46592 34988 46648
rect 34988 46592 35044 46648
rect 35044 46592 35048 46648
rect 34984 46588 35048 46592
rect 35064 46648 35128 46652
rect 35064 46592 35068 46648
rect 35068 46592 35124 46648
rect 35124 46592 35128 46648
rect 35064 46588 35128 46592
rect 35144 46648 35208 46652
rect 35144 46592 35148 46648
rect 35148 46592 35204 46648
rect 35204 46592 35208 46648
rect 35144 46588 35208 46592
rect 35224 46648 35288 46652
rect 35224 46592 35228 46648
rect 35228 46592 35284 46648
rect 35284 46592 35288 46648
rect 35224 46588 35288 46592
rect 19624 45982 19688 45986
rect 19624 45926 19628 45982
rect 19628 45926 19684 45982
rect 19684 45926 19688 45982
rect 19624 45922 19688 45926
rect 19704 45982 19768 45986
rect 19704 45926 19708 45982
rect 19708 45926 19764 45982
rect 19764 45926 19768 45982
rect 19704 45922 19768 45926
rect 19784 45982 19848 45986
rect 19784 45926 19788 45982
rect 19788 45926 19844 45982
rect 19844 45926 19848 45982
rect 19784 45922 19848 45926
rect 19864 45982 19928 45986
rect 19864 45926 19868 45982
rect 19868 45926 19924 45982
rect 19924 45926 19928 45982
rect 19864 45922 19928 45926
rect 50344 45982 50408 45986
rect 50344 45926 50348 45982
rect 50348 45926 50404 45982
rect 50404 45926 50408 45982
rect 50344 45922 50408 45926
rect 50424 45982 50488 45986
rect 50424 45926 50428 45982
rect 50428 45926 50484 45982
rect 50484 45926 50488 45982
rect 50424 45922 50488 45926
rect 50504 45982 50568 45986
rect 50504 45926 50508 45982
rect 50508 45926 50564 45982
rect 50564 45926 50568 45982
rect 50504 45922 50568 45926
rect 50584 45982 50648 45986
rect 50584 45926 50588 45982
rect 50588 45926 50644 45982
rect 50644 45926 50648 45982
rect 50584 45922 50648 45926
rect 4264 45316 4328 45320
rect 4264 45260 4268 45316
rect 4268 45260 4324 45316
rect 4324 45260 4328 45316
rect 4264 45256 4328 45260
rect 4344 45316 4408 45320
rect 4344 45260 4348 45316
rect 4348 45260 4404 45316
rect 4404 45260 4408 45316
rect 4344 45256 4408 45260
rect 4424 45316 4488 45320
rect 4424 45260 4428 45316
rect 4428 45260 4484 45316
rect 4484 45260 4488 45316
rect 4424 45256 4488 45260
rect 4504 45316 4568 45320
rect 4504 45260 4508 45316
rect 4508 45260 4564 45316
rect 4564 45260 4568 45316
rect 4504 45256 4568 45260
rect 34984 45316 35048 45320
rect 34984 45260 34988 45316
rect 34988 45260 35044 45316
rect 35044 45260 35048 45316
rect 34984 45256 35048 45260
rect 35064 45316 35128 45320
rect 35064 45260 35068 45316
rect 35068 45260 35124 45316
rect 35124 45260 35128 45316
rect 35064 45256 35128 45260
rect 35144 45316 35208 45320
rect 35144 45260 35148 45316
rect 35148 45260 35204 45316
rect 35204 45260 35208 45316
rect 35144 45256 35208 45260
rect 35224 45316 35288 45320
rect 35224 45260 35228 45316
rect 35228 45260 35284 45316
rect 35284 45260 35288 45316
rect 35224 45256 35288 45260
rect 19624 44650 19688 44654
rect 19624 44594 19628 44650
rect 19628 44594 19684 44650
rect 19684 44594 19688 44650
rect 19624 44590 19688 44594
rect 19704 44650 19768 44654
rect 19704 44594 19708 44650
rect 19708 44594 19764 44650
rect 19764 44594 19768 44650
rect 19704 44590 19768 44594
rect 19784 44650 19848 44654
rect 19784 44594 19788 44650
rect 19788 44594 19844 44650
rect 19844 44594 19848 44650
rect 19784 44590 19848 44594
rect 19864 44650 19928 44654
rect 19864 44594 19868 44650
rect 19868 44594 19924 44650
rect 19924 44594 19928 44650
rect 19864 44590 19928 44594
rect 50344 44650 50408 44654
rect 50344 44594 50348 44650
rect 50348 44594 50404 44650
rect 50404 44594 50408 44650
rect 50344 44590 50408 44594
rect 50424 44650 50488 44654
rect 50424 44594 50428 44650
rect 50428 44594 50484 44650
rect 50484 44594 50488 44650
rect 50424 44590 50488 44594
rect 50504 44650 50568 44654
rect 50504 44594 50508 44650
rect 50508 44594 50564 44650
rect 50564 44594 50568 44650
rect 50504 44590 50568 44594
rect 50584 44650 50648 44654
rect 50584 44594 50588 44650
rect 50588 44594 50644 44650
rect 50644 44594 50648 44650
rect 50584 44590 50648 44594
rect 4264 43984 4328 43988
rect 4264 43928 4268 43984
rect 4268 43928 4324 43984
rect 4324 43928 4328 43984
rect 4264 43924 4328 43928
rect 4344 43984 4408 43988
rect 4344 43928 4348 43984
rect 4348 43928 4404 43984
rect 4404 43928 4408 43984
rect 4344 43924 4408 43928
rect 4424 43984 4488 43988
rect 4424 43928 4428 43984
rect 4428 43928 4484 43984
rect 4484 43928 4488 43984
rect 4424 43924 4488 43928
rect 4504 43984 4568 43988
rect 4504 43928 4508 43984
rect 4508 43928 4564 43984
rect 4564 43928 4568 43984
rect 4504 43924 4568 43928
rect 34984 43984 35048 43988
rect 34984 43928 34988 43984
rect 34988 43928 35044 43984
rect 35044 43928 35048 43984
rect 34984 43924 35048 43928
rect 35064 43984 35128 43988
rect 35064 43928 35068 43984
rect 35068 43928 35124 43984
rect 35124 43928 35128 43984
rect 35064 43924 35128 43928
rect 35144 43984 35208 43988
rect 35144 43928 35148 43984
rect 35148 43928 35204 43984
rect 35204 43928 35208 43984
rect 35144 43924 35208 43928
rect 35224 43984 35288 43988
rect 35224 43928 35228 43984
rect 35228 43928 35284 43984
rect 35284 43928 35288 43984
rect 35224 43924 35288 43928
rect 19624 43318 19688 43322
rect 19624 43262 19628 43318
rect 19628 43262 19684 43318
rect 19684 43262 19688 43318
rect 19624 43258 19688 43262
rect 19704 43318 19768 43322
rect 19704 43262 19708 43318
rect 19708 43262 19764 43318
rect 19764 43262 19768 43318
rect 19704 43258 19768 43262
rect 19784 43318 19848 43322
rect 19784 43262 19788 43318
rect 19788 43262 19844 43318
rect 19844 43262 19848 43318
rect 19784 43258 19848 43262
rect 19864 43318 19928 43322
rect 19864 43262 19868 43318
rect 19868 43262 19924 43318
rect 19924 43262 19928 43318
rect 19864 43258 19928 43262
rect 50344 43318 50408 43322
rect 50344 43262 50348 43318
rect 50348 43262 50404 43318
rect 50404 43262 50408 43318
rect 50344 43258 50408 43262
rect 50424 43318 50488 43322
rect 50424 43262 50428 43318
rect 50428 43262 50484 43318
rect 50484 43262 50488 43318
rect 50424 43258 50488 43262
rect 50504 43318 50568 43322
rect 50504 43262 50508 43318
rect 50508 43262 50564 43318
rect 50564 43262 50568 43318
rect 50504 43258 50568 43262
rect 50584 43318 50648 43322
rect 50584 43262 50588 43318
rect 50588 43262 50644 43318
rect 50644 43262 50648 43318
rect 50584 43258 50648 43262
rect 4264 42652 4328 42656
rect 4264 42596 4268 42652
rect 4268 42596 4324 42652
rect 4324 42596 4328 42652
rect 4264 42592 4328 42596
rect 4344 42652 4408 42656
rect 4344 42596 4348 42652
rect 4348 42596 4404 42652
rect 4404 42596 4408 42652
rect 4344 42592 4408 42596
rect 4424 42652 4488 42656
rect 4424 42596 4428 42652
rect 4428 42596 4484 42652
rect 4484 42596 4488 42652
rect 4424 42592 4488 42596
rect 4504 42652 4568 42656
rect 4504 42596 4508 42652
rect 4508 42596 4564 42652
rect 4564 42596 4568 42652
rect 4504 42592 4568 42596
rect 34984 42652 35048 42656
rect 34984 42596 34988 42652
rect 34988 42596 35044 42652
rect 35044 42596 35048 42652
rect 34984 42592 35048 42596
rect 35064 42652 35128 42656
rect 35064 42596 35068 42652
rect 35068 42596 35124 42652
rect 35124 42596 35128 42652
rect 35064 42592 35128 42596
rect 35144 42652 35208 42656
rect 35144 42596 35148 42652
rect 35148 42596 35204 42652
rect 35204 42596 35208 42652
rect 35144 42592 35208 42596
rect 35224 42652 35288 42656
rect 35224 42596 35228 42652
rect 35228 42596 35284 42652
rect 35284 42596 35288 42652
rect 35224 42592 35288 42596
rect 19624 41986 19688 41990
rect 19624 41930 19628 41986
rect 19628 41930 19684 41986
rect 19684 41930 19688 41986
rect 19624 41926 19688 41930
rect 19704 41986 19768 41990
rect 19704 41930 19708 41986
rect 19708 41930 19764 41986
rect 19764 41930 19768 41986
rect 19704 41926 19768 41930
rect 19784 41986 19848 41990
rect 19784 41930 19788 41986
rect 19788 41930 19844 41986
rect 19844 41930 19848 41986
rect 19784 41926 19848 41930
rect 19864 41986 19928 41990
rect 19864 41930 19868 41986
rect 19868 41930 19924 41986
rect 19924 41930 19928 41986
rect 19864 41926 19928 41930
rect 50344 41986 50408 41990
rect 50344 41930 50348 41986
rect 50348 41930 50404 41986
rect 50404 41930 50408 41986
rect 50344 41926 50408 41930
rect 50424 41986 50488 41990
rect 50424 41930 50428 41986
rect 50428 41930 50484 41986
rect 50484 41930 50488 41986
rect 50424 41926 50488 41930
rect 50504 41986 50568 41990
rect 50504 41930 50508 41986
rect 50508 41930 50564 41986
rect 50564 41930 50568 41986
rect 50504 41926 50568 41930
rect 50584 41986 50648 41990
rect 50584 41930 50588 41986
rect 50588 41930 50644 41986
rect 50644 41930 50648 41986
rect 50584 41926 50648 41930
rect 4264 41320 4328 41324
rect 4264 41264 4268 41320
rect 4268 41264 4324 41320
rect 4324 41264 4328 41320
rect 4264 41260 4328 41264
rect 4344 41320 4408 41324
rect 4344 41264 4348 41320
rect 4348 41264 4404 41320
rect 4404 41264 4408 41320
rect 4344 41260 4408 41264
rect 4424 41320 4488 41324
rect 4424 41264 4428 41320
rect 4428 41264 4484 41320
rect 4484 41264 4488 41320
rect 4424 41260 4488 41264
rect 4504 41320 4568 41324
rect 4504 41264 4508 41320
rect 4508 41264 4564 41320
rect 4564 41264 4568 41320
rect 4504 41260 4568 41264
rect 34984 41320 35048 41324
rect 34984 41264 34988 41320
rect 34988 41264 35044 41320
rect 35044 41264 35048 41320
rect 34984 41260 35048 41264
rect 35064 41320 35128 41324
rect 35064 41264 35068 41320
rect 35068 41264 35124 41320
rect 35124 41264 35128 41320
rect 35064 41260 35128 41264
rect 35144 41320 35208 41324
rect 35144 41264 35148 41320
rect 35148 41264 35204 41320
rect 35204 41264 35208 41320
rect 35144 41260 35208 41264
rect 35224 41320 35288 41324
rect 35224 41264 35228 41320
rect 35228 41264 35284 41320
rect 35284 41264 35288 41320
rect 35224 41260 35288 41264
rect 19624 40654 19688 40658
rect 19624 40598 19628 40654
rect 19628 40598 19684 40654
rect 19684 40598 19688 40654
rect 19624 40594 19688 40598
rect 19704 40654 19768 40658
rect 19704 40598 19708 40654
rect 19708 40598 19764 40654
rect 19764 40598 19768 40654
rect 19704 40594 19768 40598
rect 19784 40654 19848 40658
rect 19784 40598 19788 40654
rect 19788 40598 19844 40654
rect 19844 40598 19848 40654
rect 19784 40594 19848 40598
rect 19864 40654 19928 40658
rect 19864 40598 19868 40654
rect 19868 40598 19924 40654
rect 19924 40598 19928 40654
rect 19864 40594 19928 40598
rect 50344 40654 50408 40658
rect 50344 40598 50348 40654
rect 50348 40598 50404 40654
rect 50404 40598 50408 40654
rect 50344 40594 50408 40598
rect 50424 40654 50488 40658
rect 50424 40598 50428 40654
rect 50428 40598 50484 40654
rect 50484 40598 50488 40654
rect 50424 40594 50488 40598
rect 50504 40654 50568 40658
rect 50504 40598 50508 40654
rect 50508 40598 50564 40654
rect 50564 40598 50568 40654
rect 50504 40594 50568 40598
rect 50584 40654 50648 40658
rect 50584 40598 50588 40654
rect 50588 40598 50644 40654
rect 50644 40598 50648 40654
rect 50584 40594 50648 40598
rect 4264 39988 4328 39992
rect 4264 39932 4268 39988
rect 4268 39932 4324 39988
rect 4324 39932 4328 39988
rect 4264 39928 4328 39932
rect 4344 39988 4408 39992
rect 4344 39932 4348 39988
rect 4348 39932 4404 39988
rect 4404 39932 4408 39988
rect 4344 39928 4408 39932
rect 4424 39988 4488 39992
rect 4424 39932 4428 39988
rect 4428 39932 4484 39988
rect 4484 39932 4488 39988
rect 4424 39928 4488 39932
rect 4504 39988 4568 39992
rect 4504 39932 4508 39988
rect 4508 39932 4564 39988
rect 4564 39932 4568 39988
rect 4504 39928 4568 39932
rect 34984 39988 35048 39992
rect 34984 39932 34988 39988
rect 34988 39932 35044 39988
rect 35044 39932 35048 39988
rect 34984 39928 35048 39932
rect 35064 39988 35128 39992
rect 35064 39932 35068 39988
rect 35068 39932 35124 39988
rect 35124 39932 35128 39988
rect 35064 39928 35128 39932
rect 35144 39988 35208 39992
rect 35144 39932 35148 39988
rect 35148 39932 35204 39988
rect 35204 39932 35208 39988
rect 35144 39928 35208 39932
rect 35224 39988 35288 39992
rect 35224 39932 35228 39988
rect 35228 39932 35284 39988
rect 35284 39932 35288 39988
rect 35224 39928 35288 39932
rect 19624 39322 19688 39326
rect 19624 39266 19628 39322
rect 19628 39266 19684 39322
rect 19684 39266 19688 39322
rect 19624 39262 19688 39266
rect 19704 39322 19768 39326
rect 19704 39266 19708 39322
rect 19708 39266 19764 39322
rect 19764 39266 19768 39322
rect 19704 39262 19768 39266
rect 19784 39322 19848 39326
rect 19784 39266 19788 39322
rect 19788 39266 19844 39322
rect 19844 39266 19848 39322
rect 19784 39262 19848 39266
rect 19864 39322 19928 39326
rect 19864 39266 19868 39322
rect 19868 39266 19924 39322
rect 19924 39266 19928 39322
rect 19864 39262 19928 39266
rect 50344 39322 50408 39326
rect 50344 39266 50348 39322
rect 50348 39266 50404 39322
rect 50404 39266 50408 39322
rect 50344 39262 50408 39266
rect 50424 39322 50488 39326
rect 50424 39266 50428 39322
rect 50428 39266 50484 39322
rect 50484 39266 50488 39322
rect 50424 39262 50488 39266
rect 50504 39322 50568 39326
rect 50504 39266 50508 39322
rect 50508 39266 50564 39322
rect 50564 39266 50568 39322
rect 50504 39262 50568 39266
rect 50584 39322 50648 39326
rect 50584 39266 50588 39322
rect 50588 39266 50644 39322
rect 50644 39266 50648 39322
rect 50584 39262 50648 39266
rect 4264 38656 4328 38660
rect 4264 38600 4268 38656
rect 4268 38600 4324 38656
rect 4324 38600 4328 38656
rect 4264 38596 4328 38600
rect 4344 38656 4408 38660
rect 4344 38600 4348 38656
rect 4348 38600 4404 38656
rect 4404 38600 4408 38656
rect 4344 38596 4408 38600
rect 4424 38656 4488 38660
rect 4424 38600 4428 38656
rect 4428 38600 4484 38656
rect 4484 38600 4488 38656
rect 4424 38596 4488 38600
rect 4504 38656 4568 38660
rect 4504 38600 4508 38656
rect 4508 38600 4564 38656
rect 4564 38600 4568 38656
rect 4504 38596 4568 38600
rect 34984 38656 35048 38660
rect 34984 38600 34988 38656
rect 34988 38600 35044 38656
rect 35044 38600 35048 38656
rect 34984 38596 35048 38600
rect 35064 38656 35128 38660
rect 35064 38600 35068 38656
rect 35068 38600 35124 38656
rect 35124 38600 35128 38656
rect 35064 38596 35128 38600
rect 35144 38656 35208 38660
rect 35144 38600 35148 38656
rect 35148 38600 35204 38656
rect 35204 38600 35208 38656
rect 35144 38596 35208 38600
rect 35224 38656 35288 38660
rect 35224 38600 35228 38656
rect 35228 38600 35284 38656
rect 35284 38600 35288 38656
rect 35224 38596 35288 38600
rect 19624 37990 19688 37994
rect 19624 37934 19628 37990
rect 19628 37934 19684 37990
rect 19684 37934 19688 37990
rect 19624 37930 19688 37934
rect 19704 37990 19768 37994
rect 19704 37934 19708 37990
rect 19708 37934 19764 37990
rect 19764 37934 19768 37990
rect 19704 37930 19768 37934
rect 19784 37990 19848 37994
rect 19784 37934 19788 37990
rect 19788 37934 19844 37990
rect 19844 37934 19848 37990
rect 19784 37930 19848 37934
rect 19864 37990 19928 37994
rect 19864 37934 19868 37990
rect 19868 37934 19924 37990
rect 19924 37934 19928 37990
rect 19864 37930 19928 37934
rect 50344 37990 50408 37994
rect 50344 37934 50348 37990
rect 50348 37934 50404 37990
rect 50404 37934 50408 37990
rect 50344 37930 50408 37934
rect 50424 37990 50488 37994
rect 50424 37934 50428 37990
rect 50428 37934 50484 37990
rect 50484 37934 50488 37990
rect 50424 37930 50488 37934
rect 50504 37990 50568 37994
rect 50504 37934 50508 37990
rect 50508 37934 50564 37990
rect 50564 37934 50568 37990
rect 50504 37930 50568 37934
rect 50584 37990 50648 37994
rect 50584 37934 50588 37990
rect 50588 37934 50644 37990
rect 50644 37934 50648 37990
rect 50584 37930 50648 37934
rect 4264 37324 4328 37328
rect 4264 37268 4268 37324
rect 4268 37268 4324 37324
rect 4324 37268 4328 37324
rect 4264 37264 4328 37268
rect 4344 37324 4408 37328
rect 4344 37268 4348 37324
rect 4348 37268 4404 37324
rect 4404 37268 4408 37324
rect 4344 37264 4408 37268
rect 4424 37324 4488 37328
rect 4424 37268 4428 37324
rect 4428 37268 4484 37324
rect 4484 37268 4488 37324
rect 4424 37264 4488 37268
rect 4504 37324 4568 37328
rect 4504 37268 4508 37324
rect 4508 37268 4564 37324
rect 4564 37268 4568 37324
rect 4504 37264 4568 37268
rect 34984 37324 35048 37328
rect 34984 37268 34988 37324
rect 34988 37268 35044 37324
rect 35044 37268 35048 37324
rect 34984 37264 35048 37268
rect 35064 37324 35128 37328
rect 35064 37268 35068 37324
rect 35068 37268 35124 37324
rect 35124 37268 35128 37324
rect 35064 37264 35128 37268
rect 35144 37324 35208 37328
rect 35144 37268 35148 37324
rect 35148 37268 35204 37324
rect 35204 37268 35208 37324
rect 35144 37264 35208 37268
rect 35224 37324 35288 37328
rect 35224 37268 35228 37324
rect 35228 37268 35284 37324
rect 35284 37268 35288 37324
rect 35224 37264 35288 37268
rect 19624 36658 19688 36662
rect 19624 36602 19628 36658
rect 19628 36602 19684 36658
rect 19684 36602 19688 36658
rect 19624 36598 19688 36602
rect 19704 36658 19768 36662
rect 19704 36602 19708 36658
rect 19708 36602 19764 36658
rect 19764 36602 19768 36658
rect 19704 36598 19768 36602
rect 19784 36658 19848 36662
rect 19784 36602 19788 36658
rect 19788 36602 19844 36658
rect 19844 36602 19848 36658
rect 19784 36598 19848 36602
rect 19864 36658 19928 36662
rect 19864 36602 19868 36658
rect 19868 36602 19924 36658
rect 19924 36602 19928 36658
rect 19864 36598 19928 36602
rect 50344 36658 50408 36662
rect 50344 36602 50348 36658
rect 50348 36602 50404 36658
rect 50404 36602 50408 36658
rect 50344 36598 50408 36602
rect 50424 36658 50488 36662
rect 50424 36602 50428 36658
rect 50428 36602 50484 36658
rect 50484 36602 50488 36658
rect 50424 36598 50488 36602
rect 50504 36658 50568 36662
rect 50504 36602 50508 36658
rect 50508 36602 50564 36658
rect 50564 36602 50568 36658
rect 50504 36598 50568 36602
rect 50584 36658 50648 36662
rect 50584 36602 50588 36658
rect 50588 36602 50644 36658
rect 50644 36602 50648 36658
rect 50584 36598 50648 36602
rect 4264 35992 4328 35996
rect 4264 35936 4268 35992
rect 4268 35936 4324 35992
rect 4324 35936 4328 35992
rect 4264 35932 4328 35936
rect 4344 35992 4408 35996
rect 4344 35936 4348 35992
rect 4348 35936 4404 35992
rect 4404 35936 4408 35992
rect 4344 35932 4408 35936
rect 4424 35992 4488 35996
rect 4424 35936 4428 35992
rect 4428 35936 4484 35992
rect 4484 35936 4488 35992
rect 4424 35932 4488 35936
rect 4504 35992 4568 35996
rect 4504 35936 4508 35992
rect 4508 35936 4564 35992
rect 4564 35936 4568 35992
rect 4504 35932 4568 35936
rect 34984 35992 35048 35996
rect 34984 35936 34988 35992
rect 34988 35936 35044 35992
rect 35044 35936 35048 35992
rect 34984 35932 35048 35936
rect 35064 35992 35128 35996
rect 35064 35936 35068 35992
rect 35068 35936 35124 35992
rect 35124 35936 35128 35992
rect 35064 35932 35128 35936
rect 35144 35992 35208 35996
rect 35144 35936 35148 35992
rect 35148 35936 35204 35992
rect 35204 35936 35208 35992
rect 35144 35932 35208 35936
rect 35224 35992 35288 35996
rect 35224 35936 35228 35992
rect 35228 35936 35284 35992
rect 35284 35936 35288 35992
rect 35224 35932 35288 35936
rect 19624 35326 19688 35330
rect 19624 35270 19628 35326
rect 19628 35270 19684 35326
rect 19684 35270 19688 35326
rect 19624 35266 19688 35270
rect 19704 35326 19768 35330
rect 19704 35270 19708 35326
rect 19708 35270 19764 35326
rect 19764 35270 19768 35326
rect 19704 35266 19768 35270
rect 19784 35326 19848 35330
rect 19784 35270 19788 35326
rect 19788 35270 19844 35326
rect 19844 35270 19848 35326
rect 19784 35266 19848 35270
rect 19864 35326 19928 35330
rect 19864 35270 19868 35326
rect 19868 35270 19924 35326
rect 19924 35270 19928 35326
rect 19864 35266 19928 35270
rect 50344 35326 50408 35330
rect 50344 35270 50348 35326
rect 50348 35270 50404 35326
rect 50404 35270 50408 35326
rect 50344 35266 50408 35270
rect 50424 35326 50488 35330
rect 50424 35270 50428 35326
rect 50428 35270 50484 35326
rect 50484 35270 50488 35326
rect 50424 35266 50488 35270
rect 50504 35326 50568 35330
rect 50504 35270 50508 35326
rect 50508 35270 50564 35326
rect 50564 35270 50568 35326
rect 50504 35266 50568 35270
rect 50584 35326 50648 35330
rect 50584 35270 50588 35326
rect 50588 35270 50644 35326
rect 50644 35270 50648 35326
rect 50584 35266 50648 35270
rect 4264 34660 4328 34664
rect 4264 34604 4268 34660
rect 4268 34604 4324 34660
rect 4324 34604 4328 34660
rect 4264 34600 4328 34604
rect 4344 34660 4408 34664
rect 4344 34604 4348 34660
rect 4348 34604 4404 34660
rect 4404 34604 4408 34660
rect 4344 34600 4408 34604
rect 4424 34660 4488 34664
rect 4424 34604 4428 34660
rect 4428 34604 4484 34660
rect 4484 34604 4488 34660
rect 4424 34600 4488 34604
rect 4504 34660 4568 34664
rect 4504 34604 4508 34660
rect 4508 34604 4564 34660
rect 4564 34604 4568 34660
rect 4504 34600 4568 34604
rect 34984 34660 35048 34664
rect 34984 34604 34988 34660
rect 34988 34604 35044 34660
rect 35044 34604 35048 34660
rect 34984 34600 35048 34604
rect 35064 34660 35128 34664
rect 35064 34604 35068 34660
rect 35068 34604 35124 34660
rect 35124 34604 35128 34660
rect 35064 34600 35128 34604
rect 35144 34660 35208 34664
rect 35144 34604 35148 34660
rect 35148 34604 35204 34660
rect 35204 34604 35208 34660
rect 35144 34600 35208 34604
rect 35224 34660 35288 34664
rect 35224 34604 35228 34660
rect 35228 34604 35284 34660
rect 35284 34604 35288 34660
rect 35224 34600 35288 34604
rect 19624 33994 19688 33998
rect 19624 33938 19628 33994
rect 19628 33938 19684 33994
rect 19684 33938 19688 33994
rect 19624 33934 19688 33938
rect 19704 33994 19768 33998
rect 19704 33938 19708 33994
rect 19708 33938 19764 33994
rect 19764 33938 19768 33994
rect 19704 33934 19768 33938
rect 19784 33994 19848 33998
rect 19784 33938 19788 33994
rect 19788 33938 19844 33994
rect 19844 33938 19848 33994
rect 19784 33934 19848 33938
rect 19864 33994 19928 33998
rect 19864 33938 19868 33994
rect 19868 33938 19924 33994
rect 19924 33938 19928 33994
rect 19864 33934 19928 33938
rect 50344 33994 50408 33998
rect 50344 33938 50348 33994
rect 50348 33938 50404 33994
rect 50404 33938 50408 33994
rect 50344 33934 50408 33938
rect 50424 33994 50488 33998
rect 50424 33938 50428 33994
rect 50428 33938 50484 33994
rect 50484 33938 50488 33994
rect 50424 33934 50488 33938
rect 50504 33994 50568 33998
rect 50504 33938 50508 33994
rect 50508 33938 50564 33994
rect 50564 33938 50568 33994
rect 50504 33934 50568 33938
rect 50584 33994 50648 33998
rect 50584 33938 50588 33994
rect 50588 33938 50644 33994
rect 50644 33938 50648 33994
rect 50584 33934 50648 33938
rect 4264 33328 4328 33332
rect 4264 33272 4268 33328
rect 4268 33272 4324 33328
rect 4324 33272 4328 33328
rect 4264 33268 4328 33272
rect 4344 33328 4408 33332
rect 4344 33272 4348 33328
rect 4348 33272 4404 33328
rect 4404 33272 4408 33328
rect 4344 33268 4408 33272
rect 4424 33328 4488 33332
rect 4424 33272 4428 33328
rect 4428 33272 4484 33328
rect 4484 33272 4488 33328
rect 4424 33268 4488 33272
rect 4504 33328 4568 33332
rect 4504 33272 4508 33328
rect 4508 33272 4564 33328
rect 4564 33272 4568 33328
rect 4504 33268 4568 33272
rect 34984 33328 35048 33332
rect 34984 33272 34988 33328
rect 34988 33272 35044 33328
rect 35044 33272 35048 33328
rect 34984 33268 35048 33272
rect 35064 33328 35128 33332
rect 35064 33272 35068 33328
rect 35068 33272 35124 33328
rect 35124 33272 35128 33328
rect 35064 33268 35128 33272
rect 35144 33328 35208 33332
rect 35144 33272 35148 33328
rect 35148 33272 35204 33328
rect 35204 33272 35208 33328
rect 35144 33268 35208 33272
rect 35224 33328 35288 33332
rect 35224 33272 35228 33328
rect 35228 33272 35284 33328
rect 35284 33272 35288 33328
rect 35224 33268 35288 33272
rect 19624 32662 19688 32666
rect 19624 32606 19628 32662
rect 19628 32606 19684 32662
rect 19684 32606 19688 32662
rect 19624 32602 19688 32606
rect 19704 32662 19768 32666
rect 19704 32606 19708 32662
rect 19708 32606 19764 32662
rect 19764 32606 19768 32662
rect 19704 32602 19768 32606
rect 19784 32662 19848 32666
rect 19784 32606 19788 32662
rect 19788 32606 19844 32662
rect 19844 32606 19848 32662
rect 19784 32602 19848 32606
rect 19864 32662 19928 32666
rect 19864 32606 19868 32662
rect 19868 32606 19924 32662
rect 19924 32606 19928 32662
rect 19864 32602 19928 32606
rect 50344 32662 50408 32666
rect 50344 32606 50348 32662
rect 50348 32606 50404 32662
rect 50404 32606 50408 32662
rect 50344 32602 50408 32606
rect 50424 32662 50488 32666
rect 50424 32606 50428 32662
rect 50428 32606 50484 32662
rect 50484 32606 50488 32662
rect 50424 32602 50488 32606
rect 50504 32662 50568 32666
rect 50504 32606 50508 32662
rect 50508 32606 50564 32662
rect 50564 32606 50568 32662
rect 50504 32602 50568 32606
rect 50584 32662 50648 32666
rect 50584 32606 50588 32662
rect 50588 32606 50644 32662
rect 50644 32606 50648 32662
rect 50584 32602 50648 32606
rect 4264 31996 4328 32000
rect 4264 31940 4268 31996
rect 4268 31940 4324 31996
rect 4324 31940 4328 31996
rect 4264 31936 4328 31940
rect 4344 31996 4408 32000
rect 4344 31940 4348 31996
rect 4348 31940 4404 31996
rect 4404 31940 4408 31996
rect 4344 31936 4408 31940
rect 4424 31996 4488 32000
rect 4424 31940 4428 31996
rect 4428 31940 4484 31996
rect 4484 31940 4488 31996
rect 4424 31936 4488 31940
rect 4504 31996 4568 32000
rect 4504 31940 4508 31996
rect 4508 31940 4564 31996
rect 4564 31940 4568 31996
rect 4504 31936 4568 31940
rect 34984 31996 35048 32000
rect 34984 31940 34988 31996
rect 34988 31940 35044 31996
rect 35044 31940 35048 31996
rect 34984 31936 35048 31940
rect 35064 31996 35128 32000
rect 35064 31940 35068 31996
rect 35068 31940 35124 31996
rect 35124 31940 35128 31996
rect 35064 31936 35128 31940
rect 35144 31996 35208 32000
rect 35144 31940 35148 31996
rect 35148 31940 35204 31996
rect 35204 31940 35208 31996
rect 35144 31936 35208 31940
rect 35224 31996 35288 32000
rect 35224 31940 35228 31996
rect 35228 31940 35284 31996
rect 35284 31940 35288 31996
rect 35224 31936 35288 31940
rect 19624 31330 19688 31334
rect 19624 31274 19628 31330
rect 19628 31274 19684 31330
rect 19684 31274 19688 31330
rect 19624 31270 19688 31274
rect 19704 31330 19768 31334
rect 19704 31274 19708 31330
rect 19708 31274 19764 31330
rect 19764 31274 19768 31330
rect 19704 31270 19768 31274
rect 19784 31330 19848 31334
rect 19784 31274 19788 31330
rect 19788 31274 19844 31330
rect 19844 31274 19848 31330
rect 19784 31270 19848 31274
rect 19864 31330 19928 31334
rect 19864 31274 19868 31330
rect 19868 31274 19924 31330
rect 19924 31274 19928 31330
rect 19864 31270 19928 31274
rect 50344 31330 50408 31334
rect 50344 31274 50348 31330
rect 50348 31274 50404 31330
rect 50404 31274 50408 31330
rect 50344 31270 50408 31274
rect 50424 31330 50488 31334
rect 50424 31274 50428 31330
rect 50428 31274 50484 31330
rect 50484 31274 50488 31330
rect 50424 31270 50488 31274
rect 50504 31330 50568 31334
rect 50504 31274 50508 31330
rect 50508 31274 50564 31330
rect 50564 31274 50568 31330
rect 50504 31270 50568 31274
rect 50584 31330 50648 31334
rect 50584 31274 50588 31330
rect 50588 31274 50644 31330
rect 50644 31274 50648 31330
rect 50584 31270 50648 31274
rect 4264 30664 4328 30668
rect 4264 30608 4268 30664
rect 4268 30608 4324 30664
rect 4324 30608 4328 30664
rect 4264 30604 4328 30608
rect 4344 30664 4408 30668
rect 4344 30608 4348 30664
rect 4348 30608 4404 30664
rect 4404 30608 4408 30664
rect 4344 30604 4408 30608
rect 4424 30664 4488 30668
rect 4424 30608 4428 30664
rect 4428 30608 4484 30664
rect 4484 30608 4488 30664
rect 4424 30604 4488 30608
rect 4504 30664 4568 30668
rect 4504 30608 4508 30664
rect 4508 30608 4564 30664
rect 4564 30608 4568 30664
rect 4504 30604 4568 30608
rect 34984 30664 35048 30668
rect 34984 30608 34988 30664
rect 34988 30608 35044 30664
rect 35044 30608 35048 30664
rect 34984 30604 35048 30608
rect 35064 30664 35128 30668
rect 35064 30608 35068 30664
rect 35068 30608 35124 30664
rect 35124 30608 35128 30664
rect 35064 30604 35128 30608
rect 35144 30664 35208 30668
rect 35144 30608 35148 30664
rect 35148 30608 35204 30664
rect 35204 30608 35208 30664
rect 35144 30604 35208 30608
rect 35224 30664 35288 30668
rect 35224 30608 35228 30664
rect 35228 30608 35284 30664
rect 35284 30608 35288 30664
rect 35224 30604 35288 30608
rect 19624 29998 19688 30002
rect 19624 29942 19628 29998
rect 19628 29942 19684 29998
rect 19684 29942 19688 29998
rect 19624 29938 19688 29942
rect 19704 29998 19768 30002
rect 19704 29942 19708 29998
rect 19708 29942 19764 29998
rect 19764 29942 19768 29998
rect 19704 29938 19768 29942
rect 19784 29998 19848 30002
rect 19784 29942 19788 29998
rect 19788 29942 19844 29998
rect 19844 29942 19848 29998
rect 19784 29938 19848 29942
rect 19864 29998 19928 30002
rect 19864 29942 19868 29998
rect 19868 29942 19924 29998
rect 19924 29942 19928 29998
rect 19864 29938 19928 29942
rect 50344 29998 50408 30002
rect 50344 29942 50348 29998
rect 50348 29942 50404 29998
rect 50404 29942 50408 29998
rect 50344 29938 50408 29942
rect 50424 29998 50488 30002
rect 50424 29942 50428 29998
rect 50428 29942 50484 29998
rect 50484 29942 50488 29998
rect 50424 29938 50488 29942
rect 50504 29998 50568 30002
rect 50504 29942 50508 29998
rect 50508 29942 50564 29998
rect 50564 29942 50568 29998
rect 50504 29938 50568 29942
rect 50584 29998 50648 30002
rect 50584 29942 50588 29998
rect 50588 29942 50644 29998
rect 50644 29942 50648 29998
rect 50584 29938 50648 29942
rect 4264 29332 4328 29336
rect 4264 29276 4268 29332
rect 4268 29276 4324 29332
rect 4324 29276 4328 29332
rect 4264 29272 4328 29276
rect 4344 29332 4408 29336
rect 4344 29276 4348 29332
rect 4348 29276 4404 29332
rect 4404 29276 4408 29332
rect 4344 29272 4408 29276
rect 4424 29332 4488 29336
rect 4424 29276 4428 29332
rect 4428 29276 4484 29332
rect 4484 29276 4488 29332
rect 4424 29272 4488 29276
rect 4504 29332 4568 29336
rect 4504 29276 4508 29332
rect 4508 29276 4564 29332
rect 4564 29276 4568 29332
rect 4504 29272 4568 29276
rect 34984 29332 35048 29336
rect 34984 29276 34988 29332
rect 34988 29276 35044 29332
rect 35044 29276 35048 29332
rect 34984 29272 35048 29276
rect 35064 29332 35128 29336
rect 35064 29276 35068 29332
rect 35068 29276 35124 29332
rect 35124 29276 35128 29332
rect 35064 29272 35128 29276
rect 35144 29332 35208 29336
rect 35144 29276 35148 29332
rect 35148 29276 35204 29332
rect 35204 29276 35208 29332
rect 35144 29272 35208 29276
rect 35224 29332 35288 29336
rect 35224 29276 35228 29332
rect 35228 29276 35284 29332
rect 35284 29276 35288 29332
rect 35224 29272 35288 29276
rect 19624 28666 19688 28670
rect 19624 28610 19628 28666
rect 19628 28610 19684 28666
rect 19684 28610 19688 28666
rect 19624 28606 19688 28610
rect 19704 28666 19768 28670
rect 19704 28610 19708 28666
rect 19708 28610 19764 28666
rect 19764 28610 19768 28666
rect 19704 28606 19768 28610
rect 19784 28666 19848 28670
rect 19784 28610 19788 28666
rect 19788 28610 19844 28666
rect 19844 28610 19848 28666
rect 19784 28606 19848 28610
rect 19864 28666 19928 28670
rect 19864 28610 19868 28666
rect 19868 28610 19924 28666
rect 19924 28610 19928 28666
rect 19864 28606 19928 28610
rect 50344 28666 50408 28670
rect 50344 28610 50348 28666
rect 50348 28610 50404 28666
rect 50404 28610 50408 28666
rect 50344 28606 50408 28610
rect 50424 28666 50488 28670
rect 50424 28610 50428 28666
rect 50428 28610 50484 28666
rect 50484 28610 50488 28666
rect 50424 28606 50488 28610
rect 50504 28666 50568 28670
rect 50504 28610 50508 28666
rect 50508 28610 50564 28666
rect 50564 28610 50568 28666
rect 50504 28606 50568 28610
rect 50584 28666 50648 28670
rect 50584 28610 50588 28666
rect 50588 28610 50644 28666
rect 50644 28610 50648 28666
rect 50584 28606 50648 28610
rect 4264 28000 4328 28004
rect 4264 27944 4268 28000
rect 4268 27944 4324 28000
rect 4324 27944 4328 28000
rect 4264 27940 4328 27944
rect 4344 28000 4408 28004
rect 4344 27944 4348 28000
rect 4348 27944 4404 28000
rect 4404 27944 4408 28000
rect 4344 27940 4408 27944
rect 4424 28000 4488 28004
rect 4424 27944 4428 28000
rect 4428 27944 4484 28000
rect 4484 27944 4488 28000
rect 4424 27940 4488 27944
rect 4504 28000 4568 28004
rect 4504 27944 4508 28000
rect 4508 27944 4564 28000
rect 4564 27944 4568 28000
rect 4504 27940 4568 27944
rect 34984 28000 35048 28004
rect 34984 27944 34988 28000
rect 34988 27944 35044 28000
rect 35044 27944 35048 28000
rect 34984 27940 35048 27944
rect 35064 28000 35128 28004
rect 35064 27944 35068 28000
rect 35068 27944 35124 28000
rect 35124 27944 35128 28000
rect 35064 27940 35128 27944
rect 35144 28000 35208 28004
rect 35144 27944 35148 28000
rect 35148 27944 35204 28000
rect 35204 27944 35208 28000
rect 35144 27940 35208 27944
rect 35224 28000 35288 28004
rect 35224 27944 35228 28000
rect 35228 27944 35284 28000
rect 35284 27944 35288 28000
rect 35224 27940 35288 27944
rect 19624 27334 19688 27338
rect 19624 27278 19628 27334
rect 19628 27278 19684 27334
rect 19684 27278 19688 27334
rect 19624 27274 19688 27278
rect 19704 27334 19768 27338
rect 19704 27278 19708 27334
rect 19708 27278 19764 27334
rect 19764 27278 19768 27334
rect 19704 27274 19768 27278
rect 19784 27334 19848 27338
rect 19784 27278 19788 27334
rect 19788 27278 19844 27334
rect 19844 27278 19848 27334
rect 19784 27274 19848 27278
rect 19864 27334 19928 27338
rect 19864 27278 19868 27334
rect 19868 27278 19924 27334
rect 19924 27278 19928 27334
rect 19864 27274 19928 27278
rect 50344 27334 50408 27338
rect 50344 27278 50348 27334
rect 50348 27278 50404 27334
rect 50404 27278 50408 27334
rect 50344 27274 50408 27278
rect 50424 27334 50488 27338
rect 50424 27278 50428 27334
rect 50428 27278 50484 27334
rect 50484 27278 50488 27334
rect 50424 27274 50488 27278
rect 50504 27334 50568 27338
rect 50504 27278 50508 27334
rect 50508 27278 50564 27334
rect 50564 27278 50568 27334
rect 50504 27274 50568 27278
rect 50584 27334 50648 27338
rect 50584 27278 50588 27334
rect 50588 27278 50644 27334
rect 50644 27278 50648 27334
rect 50584 27274 50648 27278
rect 4264 26668 4328 26672
rect 4264 26612 4268 26668
rect 4268 26612 4324 26668
rect 4324 26612 4328 26668
rect 4264 26608 4328 26612
rect 4344 26668 4408 26672
rect 4344 26612 4348 26668
rect 4348 26612 4404 26668
rect 4404 26612 4408 26668
rect 4344 26608 4408 26612
rect 4424 26668 4488 26672
rect 4424 26612 4428 26668
rect 4428 26612 4484 26668
rect 4484 26612 4488 26668
rect 4424 26608 4488 26612
rect 4504 26668 4568 26672
rect 4504 26612 4508 26668
rect 4508 26612 4564 26668
rect 4564 26612 4568 26668
rect 4504 26608 4568 26612
rect 34984 26668 35048 26672
rect 34984 26612 34988 26668
rect 34988 26612 35044 26668
rect 35044 26612 35048 26668
rect 34984 26608 35048 26612
rect 35064 26668 35128 26672
rect 35064 26612 35068 26668
rect 35068 26612 35124 26668
rect 35124 26612 35128 26668
rect 35064 26608 35128 26612
rect 35144 26668 35208 26672
rect 35144 26612 35148 26668
rect 35148 26612 35204 26668
rect 35204 26612 35208 26668
rect 35144 26608 35208 26612
rect 35224 26668 35288 26672
rect 35224 26612 35228 26668
rect 35228 26612 35284 26668
rect 35284 26612 35288 26668
rect 35224 26608 35288 26612
rect 19624 26002 19688 26006
rect 19624 25946 19628 26002
rect 19628 25946 19684 26002
rect 19684 25946 19688 26002
rect 19624 25942 19688 25946
rect 19704 26002 19768 26006
rect 19704 25946 19708 26002
rect 19708 25946 19764 26002
rect 19764 25946 19768 26002
rect 19704 25942 19768 25946
rect 19784 26002 19848 26006
rect 19784 25946 19788 26002
rect 19788 25946 19844 26002
rect 19844 25946 19848 26002
rect 19784 25942 19848 25946
rect 19864 26002 19928 26006
rect 19864 25946 19868 26002
rect 19868 25946 19924 26002
rect 19924 25946 19928 26002
rect 19864 25942 19928 25946
rect 50344 26002 50408 26006
rect 50344 25946 50348 26002
rect 50348 25946 50404 26002
rect 50404 25946 50408 26002
rect 50344 25942 50408 25946
rect 50424 26002 50488 26006
rect 50424 25946 50428 26002
rect 50428 25946 50484 26002
rect 50484 25946 50488 26002
rect 50424 25942 50488 25946
rect 50504 26002 50568 26006
rect 50504 25946 50508 26002
rect 50508 25946 50564 26002
rect 50564 25946 50568 26002
rect 50504 25942 50568 25946
rect 50584 26002 50648 26006
rect 50584 25946 50588 26002
rect 50588 25946 50644 26002
rect 50644 25946 50648 26002
rect 50584 25942 50648 25946
rect 4264 25336 4328 25340
rect 4264 25280 4268 25336
rect 4268 25280 4324 25336
rect 4324 25280 4328 25336
rect 4264 25276 4328 25280
rect 4344 25336 4408 25340
rect 4344 25280 4348 25336
rect 4348 25280 4404 25336
rect 4404 25280 4408 25336
rect 4344 25276 4408 25280
rect 4424 25336 4488 25340
rect 4424 25280 4428 25336
rect 4428 25280 4484 25336
rect 4484 25280 4488 25336
rect 4424 25276 4488 25280
rect 4504 25336 4568 25340
rect 4504 25280 4508 25336
rect 4508 25280 4564 25336
rect 4564 25280 4568 25336
rect 4504 25276 4568 25280
rect 34984 25336 35048 25340
rect 34984 25280 34988 25336
rect 34988 25280 35044 25336
rect 35044 25280 35048 25336
rect 34984 25276 35048 25280
rect 35064 25336 35128 25340
rect 35064 25280 35068 25336
rect 35068 25280 35124 25336
rect 35124 25280 35128 25336
rect 35064 25276 35128 25280
rect 35144 25336 35208 25340
rect 35144 25280 35148 25336
rect 35148 25280 35204 25336
rect 35204 25280 35208 25336
rect 35144 25276 35208 25280
rect 35224 25336 35288 25340
rect 35224 25280 35228 25336
rect 35228 25280 35284 25336
rect 35284 25280 35288 25336
rect 35224 25276 35288 25280
rect 19624 24670 19688 24674
rect 19624 24614 19628 24670
rect 19628 24614 19684 24670
rect 19684 24614 19688 24670
rect 19624 24610 19688 24614
rect 19704 24670 19768 24674
rect 19704 24614 19708 24670
rect 19708 24614 19764 24670
rect 19764 24614 19768 24670
rect 19704 24610 19768 24614
rect 19784 24670 19848 24674
rect 19784 24614 19788 24670
rect 19788 24614 19844 24670
rect 19844 24614 19848 24670
rect 19784 24610 19848 24614
rect 19864 24670 19928 24674
rect 19864 24614 19868 24670
rect 19868 24614 19924 24670
rect 19924 24614 19928 24670
rect 19864 24610 19928 24614
rect 50344 24670 50408 24674
rect 50344 24614 50348 24670
rect 50348 24614 50404 24670
rect 50404 24614 50408 24670
rect 50344 24610 50408 24614
rect 50424 24670 50488 24674
rect 50424 24614 50428 24670
rect 50428 24614 50484 24670
rect 50484 24614 50488 24670
rect 50424 24610 50488 24614
rect 50504 24670 50568 24674
rect 50504 24614 50508 24670
rect 50508 24614 50564 24670
rect 50564 24614 50568 24670
rect 50504 24610 50568 24614
rect 50584 24670 50648 24674
rect 50584 24614 50588 24670
rect 50588 24614 50644 24670
rect 50644 24614 50648 24670
rect 50584 24610 50648 24614
rect 4264 24004 4328 24008
rect 4264 23948 4268 24004
rect 4268 23948 4324 24004
rect 4324 23948 4328 24004
rect 4264 23944 4328 23948
rect 4344 24004 4408 24008
rect 4344 23948 4348 24004
rect 4348 23948 4404 24004
rect 4404 23948 4408 24004
rect 4344 23944 4408 23948
rect 4424 24004 4488 24008
rect 4424 23948 4428 24004
rect 4428 23948 4484 24004
rect 4484 23948 4488 24004
rect 4424 23944 4488 23948
rect 4504 24004 4568 24008
rect 4504 23948 4508 24004
rect 4508 23948 4564 24004
rect 4564 23948 4568 24004
rect 4504 23944 4568 23948
rect 34984 24004 35048 24008
rect 34984 23948 34988 24004
rect 34988 23948 35044 24004
rect 35044 23948 35048 24004
rect 34984 23944 35048 23948
rect 35064 24004 35128 24008
rect 35064 23948 35068 24004
rect 35068 23948 35124 24004
rect 35124 23948 35128 24004
rect 35064 23944 35128 23948
rect 35144 24004 35208 24008
rect 35144 23948 35148 24004
rect 35148 23948 35204 24004
rect 35204 23948 35208 24004
rect 35144 23944 35208 23948
rect 35224 24004 35288 24008
rect 35224 23948 35228 24004
rect 35228 23948 35284 24004
rect 35284 23948 35288 24004
rect 35224 23944 35288 23948
rect 19624 23338 19688 23342
rect 19624 23282 19628 23338
rect 19628 23282 19684 23338
rect 19684 23282 19688 23338
rect 19624 23278 19688 23282
rect 19704 23338 19768 23342
rect 19704 23282 19708 23338
rect 19708 23282 19764 23338
rect 19764 23282 19768 23338
rect 19704 23278 19768 23282
rect 19784 23338 19848 23342
rect 19784 23282 19788 23338
rect 19788 23282 19844 23338
rect 19844 23282 19848 23338
rect 19784 23278 19848 23282
rect 19864 23338 19928 23342
rect 19864 23282 19868 23338
rect 19868 23282 19924 23338
rect 19924 23282 19928 23338
rect 19864 23278 19928 23282
rect 50344 23338 50408 23342
rect 50344 23282 50348 23338
rect 50348 23282 50404 23338
rect 50404 23282 50408 23338
rect 50344 23278 50408 23282
rect 50424 23338 50488 23342
rect 50424 23282 50428 23338
rect 50428 23282 50484 23338
rect 50484 23282 50488 23338
rect 50424 23278 50488 23282
rect 50504 23338 50568 23342
rect 50504 23282 50508 23338
rect 50508 23282 50564 23338
rect 50564 23282 50568 23338
rect 50504 23278 50568 23282
rect 50584 23338 50648 23342
rect 50584 23282 50588 23338
rect 50588 23282 50644 23338
rect 50644 23282 50648 23338
rect 50584 23278 50648 23282
rect 4264 22672 4328 22676
rect 4264 22616 4268 22672
rect 4268 22616 4324 22672
rect 4324 22616 4328 22672
rect 4264 22612 4328 22616
rect 4344 22672 4408 22676
rect 4344 22616 4348 22672
rect 4348 22616 4404 22672
rect 4404 22616 4408 22672
rect 4344 22612 4408 22616
rect 4424 22672 4488 22676
rect 4424 22616 4428 22672
rect 4428 22616 4484 22672
rect 4484 22616 4488 22672
rect 4424 22612 4488 22616
rect 4504 22672 4568 22676
rect 4504 22616 4508 22672
rect 4508 22616 4564 22672
rect 4564 22616 4568 22672
rect 4504 22612 4568 22616
rect 34984 22672 35048 22676
rect 34984 22616 34988 22672
rect 34988 22616 35044 22672
rect 35044 22616 35048 22672
rect 34984 22612 35048 22616
rect 35064 22672 35128 22676
rect 35064 22616 35068 22672
rect 35068 22616 35124 22672
rect 35124 22616 35128 22672
rect 35064 22612 35128 22616
rect 35144 22672 35208 22676
rect 35144 22616 35148 22672
rect 35148 22616 35204 22672
rect 35204 22616 35208 22672
rect 35144 22612 35208 22616
rect 35224 22672 35288 22676
rect 35224 22616 35228 22672
rect 35228 22616 35284 22672
rect 35284 22616 35288 22672
rect 35224 22612 35288 22616
rect 19624 22006 19688 22010
rect 19624 21950 19628 22006
rect 19628 21950 19684 22006
rect 19684 21950 19688 22006
rect 19624 21946 19688 21950
rect 19704 22006 19768 22010
rect 19704 21950 19708 22006
rect 19708 21950 19764 22006
rect 19764 21950 19768 22006
rect 19704 21946 19768 21950
rect 19784 22006 19848 22010
rect 19784 21950 19788 22006
rect 19788 21950 19844 22006
rect 19844 21950 19848 22006
rect 19784 21946 19848 21950
rect 19864 22006 19928 22010
rect 19864 21950 19868 22006
rect 19868 21950 19924 22006
rect 19924 21950 19928 22006
rect 19864 21946 19928 21950
rect 50344 22006 50408 22010
rect 50344 21950 50348 22006
rect 50348 21950 50404 22006
rect 50404 21950 50408 22006
rect 50344 21946 50408 21950
rect 50424 22006 50488 22010
rect 50424 21950 50428 22006
rect 50428 21950 50484 22006
rect 50484 21950 50488 22006
rect 50424 21946 50488 21950
rect 50504 22006 50568 22010
rect 50504 21950 50508 22006
rect 50508 21950 50564 22006
rect 50564 21950 50568 22006
rect 50504 21946 50568 21950
rect 50584 22006 50648 22010
rect 50584 21950 50588 22006
rect 50588 21950 50644 22006
rect 50644 21950 50648 22006
rect 50584 21946 50648 21950
rect 4264 21340 4328 21344
rect 4264 21284 4268 21340
rect 4268 21284 4324 21340
rect 4324 21284 4328 21340
rect 4264 21280 4328 21284
rect 4344 21340 4408 21344
rect 4344 21284 4348 21340
rect 4348 21284 4404 21340
rect 4404 21284 4408 21340
rect 4344 21280 4408 21284
rect 4424 21340 4488 21344
rect 4424 21284 4428 21340
rect 4428 21284 4484 21340
rect 4484 21284 4488 21340
rect 4424 21280 4488 21284
rect 4504 21340 4568 21344
rect 4504 21284 4508 21340
rect 4508 21284 4564 21340
rect 4564 21284 4568 21340
rect 4504 21280 4568 21284
rect 34984 21340 35048 21344
rect 34984 21284 34988 21340
rect 34988 21284 35044 21340
rect 35044 21284 35048 21340
rect 34984 21280 35048 21284
rect 35064 21340 35128 21344
rect 35064 21284 35068 21340
rect 35068 21284 35124 21340
rect 35124 21284 35128 21340
rect 35064 21280 35128 21284
rect 35144 21340 35208 21344
rect 35144 21284 35148 21340
rect 35148 21284 35204 21340
rect 35204 21284 35208 21340
rect 35144 21280 35208 21284
rect 35224 21340 35288 21344
rect 35224 21284 35228 21340
rect 35228 21284 35284 21340
rect 35284 21284 35288 21340
rect 35224 21280 35288 21284
rect 19624 20674 19688 20678
rect 19624 20618 19628 20674
rect 19628 20618 19684 20674
rect 19684 20618 19688 20674
rect 19624 20614 19688 20618
rect 19704 20674 19768 20678
rect 19704 20618 19708 20674
rect 19708 20618 19764 20674
rect 19764 20618 19768 20674
rect 19704 20614 19768 20618
rect 19784 20674 19848 20678
rect 19784 20618 19788 20674
rect 19788 20618 19844 20674
rect 19844 20618 19848 20674
rect 19784 20614 19848 20618
rect 19864 20674 19928 20678
rect 19864 20618 19868 20674
rect 19868 20618 19924 20674
rect 19924 20618 19928 20674
rect 19864 20614 19928 20618
rect 50344 20674 50408 20678
rect 50344 20618 50348 20674
rect 50348 20618 50404 20674
rect 50404 20618 50408 20674
rect 50344 20614 50408 20618
rect 50424 20674 50488 20678
rect 50424 20618 50428 20674
rect 50428 20618 50484 20674
rect 50484 20618 50488 20674
rect 50424 20614 50488 20618
rect 50504 20674 50568 20678
rect 50504 20618 50508 20674
rect 50508 20618 50564 20674
rect 50564 20618 50568 20674
rect 50504 20614 50568 20618
rect 50584 20674 50648 20678
rect 50584 20618 50588 20674
rect 50588 20618 50644 20674
rect 50644 20618 50648 20674
rect 50584 20614 50648 20618
rect 4264 20008 4328 20012
rect 4264 19952 4268 20008
rect 4268 19952 4324 20008
rect 4324 19952 4328 20008
rect 4264 19948 4328 19952
rect 4344 20008 4408 20012
rect 4344 19952 4348 20008
rect 4348 19952 4404 20008
rect 4404 19952 4408 20008
rect 4344 19948 4408 19952
rect 4424 20008 4488 20012
rect 4424 19952 4428 20008
rect 4428 19952 4484 20008
rect 4484 19952 4488 20008
rect 4424 19948 4488 19952
rect 4504 20008 4568 20012
rect 4504 19952 4508 20008
rect 4508 19952 4564 20008
rect 4564 19952 4568 20008
rect 4504 19948 4568 19952
rect 34984 20008 35048 20012
rect 34984 19952 34988 20008
rect 34988 19952 35044 20008
rect 35044 19952 35048 20008
rect 34984 19948 35048 19952
rect 35064 20008 35128 20012
rect 35064 19952 35068 20008
rect 35068 19952 35124 20008
rect 35124 19952 35128 20008
rect 35064 19948 35128 19952
rect 35144 20008 35208 20012
rect 35144 19952 35148 20008
rect 35148 19952 35204 20008
rect 35204 19952 35208 20008
rect 35144 19948 35208 19952
rect 35224 20008 35288 20012
rect 35224 19952 35228 20008
rect 35228 19952 35284 20008
rect 35284 19952 35288 20008
rect 35224 19948 35288 19952
rect 19624 19342 19688 19346
rect 19624 19286 19628 19342
rect 19628 19286 19684 19342
rect 19684 19286 19688 19342
rect 19624 19282 19688 19286
rect 19704 19342 19768 19346
rect 19704 19286 19708 19342
rect 19708 19286 19764 19342
rect 19764 19286 19768 19342
rect 19704 19282 19768 19286
rect 19784 19342 19848 19346
rect 19784 19286 19788 19342
rect 19788 19286 19844 19342
rect 19844 19286 19848 19342
rect 19784 19282 19848 19286
rect 19864 19342 19928 19346
rect 19864 19286 19868 19342
rect 19868 19286 19924 19342
rect 19924 19286 19928 19342
rect 19864 19282 19928 19286
rect 50344 19342 50408 19346
rect 50344 19286 50348 19342
rect 50348 19286 50404 19342
rect 50404 19286 50408 19342
rect 50344 19282 50408 19286
rect 50424 19342 50488 19346
rect 50424 19286 50428 19342
rect 50428 19286 50484 19342
rect 50484 19286 50488 19342
rect 50424 19282 50488 19286
rect 50504 19342 50568 19346
rect 50504 19286 50508 19342
rect 50508 19286 50564 19342
rect 50564 19286 50568 19342
rect 50504 19282 50568 19286
rect 50584 19342 50648 19346
rect 50584 19286 50588 19342
rect 50588 19286 50644 19342
rect 50644 19286 50648 19342
rect 50584 19282 50648 19286
rect 4264 18676 4328 18680
rect 4264 18620 4268 18676
rect 4268 18620 4324 18676
rect 4324 18620 4328 18676
rect 4264 18616 4328 18620
rect 4344 18676 4408 18680
rect 4344 18620 4348 18676
rect 4348 18620 4404 18676
rect 4404 18620 4408 18676
rect 4344 18616 4408 18620
rect 4424 18676 4488 18680
rect 4424 18620 4428 18676
rect 4428 18620 4484 18676
rect 4484 18620 4488 18676
rect 4424 18616 4488 18620
rect 4504 18676 4568 18680
rect 4504 18620 4508 18676
rect 4508 18620 4564 18676
rect 4564 18620 4568 18676
rect 4504 18616 4568 18620
rect 34984 18676 35048 18680
rect 34984 18620 34988 18676
rect 34988 18620 35044 18676
rect 35044 18620 35048 18676
rect 34984 18616 35048 18620
rect 35064 18676 35128 18680
rect 35064 18620 35068 18676
rect 35068 18620 35124 18676
rect 35124 18620 35128 18676
rect 35064 18616 35128 18620
rect 35144 18676 35208 18680
rect 35144 18620 35148 18676
rect 35148 18620 35204 18676
rect 35204 18620 35208 18676
rect 35144 18616 35208 18620
rect 35224 18676 35288 18680
rect 35224 18620 35228 18676
rect 35228 18620 35284 18676
rect 35284 18620 35288 18676
rect 35224 18616 35288 18620
rect 19624 18010 19688 18014
rect 19624 17954 19628 18010
rect 19628 17954 19684 18010
rect 19684 17954 19688 18010
rect 19624 17950 19688 17954
rect 19704 18010 19768 18014
rect 19704 17954 19708 18010
rect 19708 17954 19764 18010
rect 19764 17954 19768 18010
rect 19704 17950 19768 17954
rect 19784 18010 19848 18014
rect 19784 17954 19788 18010
rect 19788 17954 19844 18010
rect 19844 17954 19848 18010
rect 19784 17950 19848 17954
rect 19864 18010 19928 18014
rect 19864 17954 19868 18010
rect 19868 17954 19924 18010
rect 19924 17954 19928 18010
rect 19864 17950 19928 17954
rect 50344 18010 50408 18014
rect 50344 17954 50348 18010
rect 50348 17954 50404 18010
rect 50404 17954 50408 18010
rect 50344 17950 50408 17954
rect 50424 18010 50488 18014
rect 50424 17954 50428 18010
rect 50428 17954 50484 18010
rect 50484 17954 50488 18010
rect 50424 17950 50488 17954
rect 50504 18010 50568 18014
rect 50504 17954 50508 18010
rect 50508 17954 50564 18010
rect 50564 17954 50568 18010
rect 50504 17950 50568 17954
rect 50584 18010 50648 18014
rect 50584 17954 50588 18010
rect 50588 17954 50644 18010
rect 50644 17954 50648 18010
rect 50584 17950 50648 17954
rect 4264 17344 4328 17348
rect 4264 17288 4268 17344
rect 4268 17288 4324 17344
rect 4324 17288 4328 17344
rect 4264 17284 4328 17288
rect 4344 17344 4408 17348
rect 4344 17288 4348 17344
rect 4348 17288 4404 17344
rect 4404 17288 4408 17344
rect 4344 17284 4408 17288
rect 4424 17344 4488 17348
rect 4424 17288 4428 17344
rect 4428 17288 4484 17344
rect 4484 17288 4488 17344
rect 4424 17284 4488 17288
rect 4504 17344 4568 17348
rect 4504 17288 4508 17344
rect 4508 17288 4564 17344
rect 4564 17288 4568 17344
rect 4504 17284 4568 17288
rect 34984 17344 35048 17348
rect 34984 17288 34988 17344
rect 34988 17288 35044 17344
rect 35044 17288 35048 17344
rect 34984 17284 35048 17288
rect 35064 17344 35128 17348
rect 35064 17288 35068 17344
rect 35068 17288 35124 17344
rect 35124 17288 35128 17344
rect 35064 17284 35128 17288
rect 35144 17344 35208 17348
rect 35144 17288 35148 17344
rect 35148 17288 35204 17344
rect 35204 17288 35208 17344
rect 35144 17284 35208 17288
rect 35224 17344 35288 17348
rect 35224 17288 35228 17344
rect 35228 17288 35284 17344
rect 35284 17288 35288 17344
rect 35224 17284 35288 17288
rect 19624 16678 19688 16682
rect 19624 16622 19628 16678
rect 19628 16622 19684 16678
rect 19684 16622 19688 16678
rect 19624 16618 19688 16622
rect 19704 16678 19768 16682
rect 19704 16622 19708 16678
rect 19708 16622 19764 16678
rect 19764 16622 19768 16678
rect 19704 16618 19768 16622
rect 19784 16678 19848 16682
rect 19784 16622 19788 16678
rect 19788 16622 19844 16678
rect 19844 16622 19848 16678
rect 19784 16618 19848 16622
rect 19864 16678 19928 16682
rect 19864 16622 19868 16678
rect 19868 16622 19924 16678
rect 19924 16622 19928 16678
rect 19864 16618 19928 16622
rect 50344 16678 50408 16682
rect 50344 16622 50348 16678
rect 50348 16622 50404 16678
rect 50404 16622 50408 16678
rect 50344 16618 50408 16622
rect 50424 16678 50488 16682
rect 50424 16622 50428 16678
rect 50428 16622 50484 16678
rect 50484 16622 50488 16678
rect 50424 16618 50488 16622
rect 50504 16678 50568 16682
rect 50504 16622 50508 16678
rect 50508 16622 50564 16678
rect 50564 16622 50568 16678
rect 50504 16618 50568 16622
rect 50584 16678 50648 16682
rect 50584 16622 50588 16678
rect 50588 16622 50644 16678
rect 50644 16622 50648 16678
rect 50584 16618 50648 16622
rect 4264 16012 4328 16016
rect 4264 15956 4268 16012
rect 4268 15956 4324 16012
rect 4324 15956 4328 16012
rect 4264 15952 4328 15956
rect 4344 16012 4408 16016
rect 4344 15956 4348 16012
rect 4348 15956 4404 16012
rect 4404 15956 4408 16012
rect 4344 15952 4408 15956
rect 4424 16012 4488 16016
rect 4424 15956 4428 16012
rect 4428 15956 4484 16012
rect 4484 15956 4488 16012
rect 4424 15952 4488 15956
rect 4504 16012 4568 16016
rect 4504 15956 4508 16012
rect 4508 15956 4564 16012
rect 4564 15956 4568 16012
rect 4504 15952 4568 15956
rect 34984 16012 35048 16016
rect 34984 15956 34988 16012
rect 34988 15956 35044 16012
rect 35044 15956 35048 16012
rect 34984 15952 35048 15956
rect 35064 16012 35128 16016
rect 35064 15956 35068 16012
rect 35068 15956 35124 16012
rect 35124 15956 35128 16012
rect 35064 15952 35128 15956
rect 35144 16012 35208 16016
rect 35144 15956 35148 16012
rect 35148 15956 35204 16012
rect 35204 15956 35208 16012
rect 35144 15952 35208 15956
rect 35224 16012 35288 16016
rect 35224 15956 35228 16012
rect 35228 15956 35284 16012
rect 35284 15956 35288 16012
rect 35224 15952 35288 15956
rect 19624 15346 19688 15350
rect 19624 15290 19628 15346
rect 19628 15290 19684 15346
rect 19684 15290 19688 15346
rect 19624 15286 19688 15290
rect 19704 15346 19768 15350
rect 19704 15290 19708 15346
rect 19708 15290 19764 15346
rect 19764 15290 19768 15346
rect 19704 15286 19768 15290
rect 19784 15346 19848 15350
rect 19784 15290 19788 15346
rect 19788 15290 19844 15346
rect 19844 15290 19848 15346
rect 19784 15286 19848 15290
rect 19864 15346 19928 15350
rect 19864 15290 19868 15346
rect 19868 15290 19924 15346
rect 19924 15290 19928 15346
rect 19864 15286 19928 15290
rect 50344 15346 50408 15350
rect 50344 15290 50348 15346
rect 50348 15290 50404 15346
rect 50404 15290 50408 15346
rect 50344 15286 50408 15290
rect 50424 15346 50488 15350
rect 50424 15290 50428 15346
rect 50428 15290 50484 15346
rect 50484 15290 50488 15346
rect 50424 15286 50488 15290
rect 50504 15346 50568 15350
rect 50504 15290 50508 15346
rect 50508 15290 50564 15346
rect 50564 15290 50568 15346
rect 50504 15286 50568 15290
rect 50584 15346 50648 15350
rect 50584 15290 50588 15346
rect 50588 15290 50644 15346
rect 50644 15290 50648 15346
rect 50584 15286 50648 15290
rect 4264 14680 4328 14684
rect 4264 14624 4268 14680
rect 4268 14624 4324 14680
rect 4324 14624 4328 14680
rect 4264 14620 4328 14624
rect 4344 14680 4408 14684
rect 4344 14624 4348 14680
rect 4348 14624 4404 14680
rect 4404 14624 4408 14680
rect 4344 14620 4408 14624
rect 4424 14680 4488 14684
rect 4424 14624 4428 14680
rect 4428 14624 4484 14680
rect 4484 14624 4488 14680
rect 4424 14620 4488 14624
rect 4504 14680 4568 14684
rect 4504 14624 4508 14680
rect 4508 14624 4564 14680
rect 4564 14624 4568 14680
rect 4504 14620 4568 14624
rect 34984 14680 35048 14684
rect 34984 14624 34988 14680
rect 34988 14624 35044 14680
rect 35044 14624 35048 14680
rect 34984 14620 35048 14624
rect 35064 14680 35128 14684
rect 35064 14624 35068 14680
rect 35068 14624 35124 14680
rect 35124 14624 35128 14680
rect 35064 14620 35128 14624
rect 35144 14680 35208 14684
rect 35144 14624 35148 14680
rect 35148 14624 35204 14680
rect 35204 14624 35208 14680
rect 35144 14620 35208 14624
rect 35224 14680 35288 14684
rect 35224 14624 35228 14680
rect 35228 14624 35284 14680
rect 35284 14624 35288 14680
rect 35224 14620 35288 14624
rect 19624 14014 19688 14018
rect 19624 13958 19628 14014
rect 19628 13958 19684 14014
rect 19684 13958 19688 14014
rect 19624 13954 19688 13958
rect 19704 14014 19768 14018
rect 19704 13958 19708 14014
rect 19708 13958 19764 14014
rect 19764 13958 19768 14014
rect 19704 13954 19768 13958
rect 19784 14014 19848 14018
rect 19784 13958 19788 14014
rect 19788 13958 19844 14014
rect 19844 13958 19848 14014
rect 19784 13954 19848 13958
rect 19864 14014 19928 14018
rect 19864 13958 19868 14014
rect 19868 13958 19924 14014
rect 19924 13958 19928 14014
rect 19864 13954 19928 13958
rect 50344 14014 50408 14018
rect 50344 13958 50348 14014
rect 50348 13958 50404 14014
rect 50404 13958 50408 14014
rect 50344 13954 50408 13958
rect 50424 14014 50488 14018
rect 50424 13958 50428 14014
rect 50428 13958 50484 14014
rect 50484 13958 50488 14014
rect 50424 13954 50488 13958
rect 50504 14014 50568 14018
rect 50504 13958 50508 14014
rect 50508 13958 50564 14014
rect 50564 13958 50568 14014
rect 50504 13954 50568 13958
rect 50584 14014 50648 14018
rect 50584 13958 50588 14014
rect 50588 13958 50644 14014
rect 50644 13958 50648 14014
rect 50584 13954 50648 13958
rect 4264 13348 4328 13352
rect 4264 13292 4268 13348
rect 4268 13292 4324 13348
rect 4324 13292 4328 13348
rect 4264 13288 4328 13292
rect 4344 13348 4408 13352
rect 4344 13292 4348 13348
rect 4348 13292 4404 13348
rect 4404 13292 4408 13348
rect 4344 13288 4408 13292
rect 4424 13348 4488 13352
rect 4424 13292 4428 13348
rect 4428 13292 4484 13348
rect 4484 13292 4488 13348
rect 4424 13288 4488 13292
rect 4504 13348 4568 13352
rect 4504 13292 4508 13348
rect 4508 13292 4564 13348
rect 4564 13292 4568 13348
rect 4504 13288 4568 13292
rect 34984 13348 35048 13352
rect 34984 13292 34988 13348
rect 34988 13292 35044 13348
rect 35044 13292 35048 13348
rect 34984 13288 35048 13292
rect 35064 13348 35128 13352
rect 35064 13292 35068 13348
rect 35068 13292 35124 13348
rect 35124 13292 35128 13348
rect 35064 13288 35128 13292
rect 35144 13348 35208 13352
rect 35144 13292 35148 13348
rect 35148 13292 35204 13348
rect 35204 13292 35208 13348
rect 35144 13288 35208 13292
rect 35224 13348 35288 13352
rect 35224 13292 35228 13348
rect 35228 13292 35284 13348
rect 35284 13292 35288 13348
rect 35224 13288 35288 13292
rect 19624 12682 19688 12686
rect 19624 12626 19628 12682
rect 19628 12626 19684 12682
rect 19684 12626 19688 12682
rect 19624 12622 19688 12626
rect 19704 12682 19768 12686
rect 19704 12626 19708 12682
rect 19708 12626 19764 12682
rect 19764 12626 19768 12682
rect 19704 12622 19768 12626
rect 19784 12682 19848 12686
rect 19784 12626 19788 12682
rect 19788 12626 19844 12682
rect 19844 12626 19848 12682
rect 19784 12622 19848 12626
rect 19864 12682 19928 12686
rect 19864 12626 19868 12682
rect 19868 12626 19924 12682
rect 19924 12626 19928 12682
rect 19864 12622 19928 12626
rect 50344 12682 50408 12686
rect 50344 12626 50348 12682
rect 50348 12626 50404 12682
rect 50404 12626 50408 12682
rect 50344 12622 50408 12626
rect 50424 12682 50488 12686
rect 50424 12626 50428 12682
rect 50428 12626 50484 12682
rect 50484 12626 50488 12682
rect 50424 12622 50488 12626
rect 50504 12682 50568 12686
rect 50504 12626 50508 12682
rect 50508 12626 50564 12682
rect 50564 12626 50568 12682
rect 50504 12622 50568 12626
rect 50584 12682 50648 12686
rect 50584 12626 50588 12682
rect 50588 12626 50644 12682
rect 50644 12626 50648 12682
rect 50584 12622 50648 12626
rect 4264 12016 4328 12020
rect 4264 11960 4268 12016
rect 4268 11960 4324 12016
rect 4324 11960 4328 12016
rect 4264 11956 4328 11960
rect 4344 12016 4408 12020
rect 4344 11960 4348 12016
rect 4348 11960 4404 12016
rect 4404 11960 4408 12016
rect 4344 11956 4408 11960
rect 4424 12016 4488 12020
rect 4424 11960 4428 12016
rect 4428 11960 4484 12016
rect 4484 11960 4488 12016
rect 4424 11956 4488 11960
rect 4504 12016 4568 12020
rect 4504 11960 4508 12016
rect 4508 11960 4564 12016
rect 4564 11960 4568 12016
rect 4504 11956 4568 11960
rect 34984 12016 35048 12020
rect 34984 11960 34988 12016
rect 34988 11960 35044 12016
rect 35044 11960 35048 12016
rect 34984 11956 35048 11960
rect 35064 12016 35128 12020
rect 35064 11960 35068 12016
rect 35068 11960 35124 12016
rect 35124 11960 35128 12016
rect 35064 11956 35128 11960
rect 35144 12016 35208 12020
rect 35144 11960 35148 12016
rect 35148 11960 35204 12016
rect 35204 11960 35208 12016
rect 35144 11956 35208 11960
rect 35224 12016 35288 12020
rect 35224 11960 35228 12016
rect 35228 11960 35284 12016
rect 35284 11960 35288 12016
rect 35224 11956 35288 11960
rect 19624 11350 19688 11354
rect 19624 11294 19628 11350
rect 19628 11294 19684 11350
rect 19684 11294 19688 11350
rect 19624 11290 19688 11294
rect 19704 11350 19768 11354
rect 19704 11294 19708 11350
rect 19708 11294 19764 11350
rect 19764 11294 19768 11350
rect 19704 11290 19768 11294
rect 19784 11350 19848 11354
rect 19784 11294 19788 11350
rect 19788 11294 19844 11350
rect 19844 11294 19848 11350
rect 19784 11290 19848 11294
rect 19864 11350 19928 11354
rect 19864 11294 19868 11350
rect 19868 11294 19924 11350
rect 19924 11294 19928 11350
rect 19864 11290 19928 11294
rect 50344 11350 50408 11354
rect 50344 11294 50348 11350
rect 50348 11294 50404 11350
rect 50404 11294 50408 11350
rect 50344 11290 50408 11294
rect 50424 11350 50488 11354
rect 50424 11294 50428 11350
rect 50428 11294 50484 11350
rect 50484 11294 50488 11350
rect 50424 11290 50488 11294
rect 50504 11350 50568 11354
rect 50504 11294 50508 11350
rect 50508 11294 50564 11350
rect 50564 11294 50568 11350
rect 50504 11290 50568 11294
rect 50584 11350 50648 11354
rect 50584 11294 50588 11350
rect 50588 11294 50644 11350
rect 50644 11294 50648 11350
rect 50584 11290 50648 11294
rect 4264 10684 4328 10688
rect 4264 10628 4268 10684
rect 4268 10628 4324 10684
rect 4324 10628 4328 10684
rect 4264 10624 4328 10628
rect 4344 10684 4408 10688
rect 4344 10628 4348 10684
rect 4348 10628 4404 10684
rect 4404 10628 4408 10684
rect 4344 10624 4408 10628
rect 4424 10684 4488 10688
rect 4424 10628 4428 10684
rect 4428 10628 4484 10684
rect 4484 10628 4488 10684
rect 4424 10624 4488 10628
rect 4504 10684 4568 10688
rect 4504 10628 4508 10684
rect 4508 10628 4564 10684
rect 4564 10628 4568 10684
rect 4504 10624 4568 10628
rect 34984 10684 35048 10688
rect 34984 10628 34988 10684
rect 34988 10628 35044 10684
rect 35044 10628 35048 10684
rect 34984 10624 35048 10628
rect 35064 10684 35128 10688
rect 35064 10628 35068 10684
rect 35068 10628 35124 10684
rect 35124 10628 35128 10684
rect 35064 10624 35128 10628
rect 35144 10684 35208 10688
rect 35144 10628 35148 10684
rect 35148 10628 35204 10684
rect 35204 10628 35208 10684
rect 35144 10624 35208 10628
rect 35224 10684 35288 10688
rect 35224 10628 35228 10684
rect 35228 10628 35284 10684
rect 35284 10628 35288 10684
rect 35224 10624 35288 10628
rect 19624 10018 19688 10022
rect 19624 9962 19628 10018
rect 19628 9962 19684 10018
rect 19684 9962 19688 10018
rect 19624 9958 19688 9962
rect 19704 10018 19768 10022
rect 19704 9962 19708 10018
rect 19708 9962 19764 10018
rect 19764 9962 19768 10018
rect 19704 9958 19768 9962
rect 19784 10018 19848 10022
rect 19784 9962 19788 10018
rect 19788 9962 19844 10018
rect 19844 9962 19848 10018
rect 19784 9958 19848 9962
rect 19864 10018 19928 10022
rect 19864 9962 19868 10018
rect 19868 9962 19924 10018
rect 19924 9962 19928 10018
rect 19864 9958 19928 9962
rect 50344 10018 50408 10022
rect 50344 9962 50348 10018
rect 50348 9962 50404 10018
rect 50404 9962 50408 10018
rect 50344 9958 50408 9962
rect 50424 10018 50488 10022
rect 50424 9962 50428 10018
rect 50428 9962 50484 10018
rect 50484 9962 50488 10018
rect 50424 9958 50488 9962
rect 50504 10018 50568 10022
rect 50504 9962 50508 10018
rect 50508 9962 50564 10018
rect 50564 9962 50568 10018
rect 50504 9958 50568 9962
rect 50584 10018 50648 10022
rect 50584 9962 50588 10018
rect 50588 9962 50644 10018
rect 50644 9962 50648 10018
rect 50584 9958 50648 9962
rect 4264 9352 4328 9356
rect 4264 9296 4268 9352
rect 4268 9296 4324 9352
rect 4324 9296 4328 9352
rect 4264 9292 4328 9296
rect 4344 9352 4408 9356
rect 4344 9296 4348 9352
rect 4348 9296 4404 9352
rect 4404 9296 4408 9352
rect 4344 9292 4408 9296
rect 4424 9352 4488 9356
rect 4424 9296 4428 9352
rect 4428 9296 4484 9352
rect 4484 9296 4488 9352
rect 4424 9292 4488 9296
rect 4504 9352 4568 9356
rect 4504 9296 4508 9352
rect 4508 9296 4564 9352
rect 4564 9296 4568 9352
rect 4504 9292 4568 9296
rect 34984 9352 35048 9356
rect 34984 9296 34988 9352
rect 34988 9296 35044 9352
rect 35044 9296 35048 9352
rect 34984 9292 35048 9296
rect 35064 9352 35128 9356
rect 35064 9296 35068 9352
rect 35068 9296 35124 9352
rect 35124 9296 35128 9352
rect 35064 9292 35128 9296
rect 35144 9352 35208 9356
rect 35144 9296 35148 9352
rect 35148 9296 35204 9352
rect 35204 9296 35208 9352
rect 35144 9292 35208 9296
rect 35224 9352 35288 9356
rect 35224 9296 35228 9352
rect 35228 9296 35284 9352
rect 35284 9296 35288 9352
rect 35224 9292 35288 9296
rect 19624 8686 19688 8690
rect 19624 8630 19628 8686
rect 19628 8630 19684 8686
rect 19684 8630 19688 8686
rect 19624 8626 19688 8630
rect 19704 8686 19768 8690
rect 19704 8630 19708 8686
rect 19708 8630 19764 8686
rect 19764 8630 19768 8686
rect 19704 8626 19768 8630
rect 19784 8686 19848 8690
rect 19784 8630 19788 8686
rect 19788 8630 19844 8686
rect 19844 8630 19848 8686
rect 19784 8626 19848 8630
rect 19864 8686 19928 8690
rect 19864 8630 19868 8686
rect 19868 8630 19924 8686
rect 19924 8630 19928 8686
rect 19864 8626 19928 8630
rect 50344 8686 50408 8690
rect 50344 8630 50348 8686
rect 50348 8630 50404 8686
rect 50404 8630 50408 8686
rect 50344 8626 50408 8630
rect 50424 8686 50488 8690
rect 50424 8630 50428 8686
rect 50428 8630 50484 8686
rect 50484 8630 50488 8686
rect 50424 8626 50488 8630
rect 50504 8686 50568 8690
rect 50504 8630 50508 8686
rect 50508 8630 50564 8686
rect 50564 8630 50568 8686
rect 50504 8626 50568 8630
rect 50584 8686 50648 8690
rect 50584 8630 50588 8686
rect 50588 8630 50644 8686
rect 50644 8630 50648 8686
rect 50584 8626 50648 8630
rect 4264 8020 4328 8024
rect 4264 7964 4268 8020
rect 4268 7964 4324 8020
rect 4324 7964 4328 8020
rect 4264 7960 4328 7964
rect 4344 8020 4408 8024
rect 4344 7964 4348 8020
rect 4348 7964 4404 8020
rect 4404 7964 4408 8020
rect 4344 7960 4408 7964
rect 4424 8020 4488 8024
rect 4424 7964 4428 8020
rect 4428 7964 4484 8020
rect 4484 7964 4488 8020
rect 4424 7960 4488 7964
rect 4504 8020 4568 8024
rect 4504 7964 4508 8020
rect 4508 7964 4564 8020
rect 4564 7964 4568 8020
rect 4504 7960 4568 7964
rect 34984 8020 35048 8024
rect 34984 7964 34988 8020
rect 34988 7964 35044 8020
rect 35044 7964 35048 8020
rect 34984 7960 35048 7964
rect 35064 8020 35128 8024
rect 35064 7964 35068 8020
rect 35068 7964 35124 8020
rect 35124 7964 35128 8020
rect 35064 7960 35128 7964
rect 35144 8020 35208 8024
rect 35144 7964 35148 8020
rect 35148 7964 35204 8020
rect 35204 7964 35208 8020
rect 35144 7960 35208 7964
rect 35224 8020 35288 8024
rect 35224 7964 35228 8020
rect 35228 7964 35284 8020
rect 35284 7964 35288 8020
rect 35224 7960 35288 7964
rect 19624 7354 19688 7358
rect 19624 7298 19628 7354
rect 19628 7298 19684 7354
rect 19684 7298 19688 7354
rect 19624 7294 19688 7298
rect 19704 7354 19768 7358
rect 19704 7298 19708 7354
rect 19708 7298 19764 7354
rect 19764 7298 19768 7354
rect 19704 7294 19768 7298
rect 19784 7354 19848 7358
rect 19784 7298 19788 7354
rect 19788 7298 19844 7354
rect 19844 7298 19848 7354
rect 19784 7294 19848 7298
rect 19864 7354 19928 7358
rect 19864 7298 19868 7354
rect 19868 7298 19924 7354
rect 19924 7298 19928 7354
rect 19864 7294 19928 7298
rect 50344 7354 50408 7358
rect 50344 7298 50348 7354
rect 50348 7298 50404 7354
rect 50404 7298 50408 7354
rect 50344 7294 50408 7298
rect 50424 7354 50488 7358
rect 50424 7298 50428 7354
rect 50428 7298 50484 7354
rect 50484 7298 50488 7354
rect 50424 7294 50488 7298
rect 50504 7354 50568 7358
rect 50504 7298 50508 7354
rect 50508 7298 50564 7354
rect 50564 7298 50568 7354
rect 50504 7294 50568 7298
rect 50584 7354 50648 7358
rect 50584 7298 50588 7354
rect 50588 7298 50644 7354
rect 50644 7298 50648 7354
rect 50584 7294 50648 7298
rect 4264 6688 4328 6692
rect 4264 6632 4268 6688
rect 4268 6632 4324 6688
rect 4324 6632 4328 6688
rect 4264 6628 4328 6632
rect 4344 6688 4408 6692
rect 4344 6632 4348 6688
rect 4348 6632 4404 6688
rect 4404 6632 4408 6688
rect 4344 6628 4408 6632
rect 4424 6688 4488 6692
rect 4424 6632 4428 6688
rect 4428 6632 4484 6688
rect 4484 6632 4488 6688
rect 4424 6628 4488 6632
rect 4504 6688 4568 6692
rect 4504 6632 4508 6688
rect 4508 6632 4564 6688
rect 4564 6632 4568 6688
rect 4504 6628 4568 6632
rect 34984 6688 35048 6692
rect 34984 6632 34988 6688
rect 34988 6632 35044 6688
rect 35044 6632 35048 6688
rect 34984 6628 35048 6632
rect 35064 6688 35128 6692
rect 35064 6632 35068 6688
rect 35068 6632 35124 6688
rect 35124 6632 35128 6688
rect 35064 6628 35128 6632
rect 35144 6688 35208 6692
rect 35144 6632 35148 6688
rect 35148 6632 35204 6688
rect 35204 6632 35208 6688
rect 35144 6628 35208 6632
rect 35224 6688 35288 6692
rect 35224 6632 35228 6688
rect 35228 6632 35284 6688
rect 35284 6632 35288 6688
rect 35224 6628 35288 6632
rect 19624 6022 19688 6026
rect 19624 5966 19628 6022
rect 19628 5966 19684 6022
rect 19684 5966 19688 6022
rect 19624 5962 19688 5966
rect 19704 6022 19768 6026
rect 19704 5966 19708 6022
rect 19708 5966 19764 6022
rect 19764 5966 19768 6022
rect 19704 5962 19768 5966
rect 19784 6022 19848 6026
rect 19784 5966 19788 6022
rect 19788 5966 19844 6022
rect 19844 5966 19848 6022
rect 19784 5962 19848 5966
rect 19864 6022 19928 6026
rect 19864 5966 19868 6022
rect 19868 5966 19924 6022
rect 19924 5966 19928 6022
rect 19864 5962 19928 5966
rect 50344 6022 50408 6026
rect 50344 5966 50348 6022
rect 50348 5966 50404 6022
rect 50404 5966 50408 6022
rect 50344 5962 50408 5966
rect 50424 6022 50488 6026
rect 50424 5966 50428 6022
rect 50428 5966 50484 6022
rect 50484 5966 50488 6022
rect 50424 5962 50488 5966
rect 50504 6022 50568 6026
rect 50504 5966 50508 6022
rect 50508 5966 50564 6022
rect 50564 5966 50568 6022
rect 50504 5962 50568 5966
rect 50584 6022 50648 6026
rect 50584 5966 50588 6022
rect 50588 5966 50644 6022
rect 50644 5966 50648 6022
rect 50584 5962 50648 5966
rect 4264 5356 4328 5360
rect 4264 5300 4268 5356
rect 4268 5300 4324 5356
rect 4324 5300 4328 5356
rect 4264 5296 4328 5300
rect 4344 5356 4408 5360
rect 4344 5300 4348 5356
rect 4348 5300 4404 5356
rect 4404 5300 4408 5356
rect 4344 5296 4408 5300
rect 4424 5356 4488 5360
rect 4424 5300 4428 5356
rect 4428 5300 4484 5356
rect 4484 5300 4488 5356
rect 4424 5296 4488 5300
rect 4504 5356 4568 5360
rect 4504 5300 4508 5356
rect 4508 5300 4564 5356
rect 4564 5300 4568 5356
rect 4504 5296 4568 5300
rect 34984 5356 35048 5360
rect 34984 5300 34988 5356
rect 34988 5300 35044 5356
rect 35044 5300 35048 5356
rect 34984 5296 35048 5300
rect 35064 5356 35128 5360
rect 35064 5300 35068 5356
rect 35068 5300 35124 5356
rect 35124 5300 35128 5356
rect 35064 5296 35128 5300
rect 35144 5356 35208 5360
rect 35144 5300 35148 5356
rect 35148 5300 35204 5356
rect 35204 5300 35208 5356
rect 35144 5296 35208 5300
rect 35224 5356 35288 5360
rect 35224 5300 35228 5356
rect 35228 5300 35284 5356
rect 35284 5300 35288 5356
rect 35224 5296 35288 5300
rect 19624 4690 19688 4694
rect 19624 4634 19628 4690
rect 19628 4634 19684 4690
rect 19684 4634 19688 4690
rect 19624 4630 19688 4634
rect 19704 4690 19768 4694
rect 19704 4634 19708 4690
rect 19708 4634 19764 4690
rect 19764 4634 19768 4690
rect 19704 4630 19768 4634
rect 19784 4690 19848 4694
rect 19784 4634 19788 4690
rect 19788 4634 19844 4690
rect 19844 4634 19848 4690
rect 19784 4630 19848 4634
rect 19864 4690 19928 4694
rect 19864 4634 19868 4690
rect 19868 4634 19924 4690
rect 19924 4634 19928 4690
rect 19864 4630 19928 4634
rect 50344 4690 50408 4694
rect 50344 4634 50348 4690
rect 50348 4634 50404 4690
rect 50404 4634 50408 4690
rect 50344 4630 50408 4634
rect 50424 4690 50488 4694
rect 50424 4634 50428 4690
rect 50428 4634 50484 4690
rect 50484 4634 50488 4690
rect 50424 4630 50488 4634
rect 50504 4690 50568 4694
rect 50504 4634 50508 4690
rect 50508 4634 50564 4690
rect 50564 4634 50568 4690
rect 50504 4630 50568 4634
rect 50584 4690 50648 4694
rect 50584 4634 50588 4690
rect 50588 4634 50644 4690
rect 50644 4634 50648 4690
rect 50584 4630 50648 4634
rect 4264 4024 4328 4028
rect 4264 3968 4268 4024
rect 4268 3968 4324 4024
rect 4324 3968 4328 4024
rect 4264 3964 4328 3968
rect 4344 4024 4408 4028
rect 4344 3968 4348 4024
rect 4348 3968 4404 4024
rect 4404 3968 4408 4024
rect 4344 3964 4408 3968
rect 4424 4024 4488 4028
rect 4424 3968 4428 4024
rect 4428 3968 4484 4024
rect 4484 3968 4488 4024
rect 4424 3964 4488 3968
rect 4504 4024 4568 4028
rect 4504 3968 4508 4024
rect 4508 3968 4564 4024
rect 4564 3968 4568 4024
rect 4504 3964 4568 3968
rect 34984 4024 35048 4028
rect 34984 3968 34988 4024
rect 34988 3968 35044 4024
rect 35044 3968 35048 4024
rect 34984 3964 35048 3968
rect 35064 4024 35128 4028
rect 35064 3968 35068 4024
rect 35068 3968 35124 4024
rect 35124 3968 35128 4024
rect 35064 3964 35128 3968
rect 35144 4024 35208 4028
rect 35144 3968 35148 4024
rect 35148 3968 35204 4024
rect 35204 3968 35208 4024
rect 35144 3964 35208 3968
rect 35224 4024 35288 4028
rect 35224 3968 35228 4024
rect 35228 3968 35284 4024
rect 35284 3968 35288 4024
rect 35224 3964 35288 3968
rect 19624 3358 19688 3362
rect 19624 3302 19628 3358
rect 19628 3302 19684 3358
rect 19684 3302 19688 3358
rect 19624 3298 19688 3302
rect 19704 3358 19768 3362
rect 19704 3302 19708 3358
rect 19708 3302 19764 3358
rect 19764 3302 19768 3358
rect 19704 3298 19768 3302
rect 19784 3358 19848 3362
rect 19784 3302 19788 3358
rect 19788 3302 19844 3358
rect 19844 3302 19848 3358
rect 19784 3298 19848 3302
rect 19864 3358 19928 3362
rect 19864 3302 19868 3358
rect 19868 3302 19924 3358
rect 19924 3302 19928 3358
rect 19864 3298 19928 3302
rect 50344 3358 50408 3362
rect 50344 3302 50348 3358
rect 50348 3302 50404 3358
rect 50404 3302 50408 3358
rect 50344 3298 50408 3302
rect 50424 3358 50488 3362
rect 50424 3302 50428 3358
rect 50428 3302 50484 3358
rect 50484 3302 50488 3358
rect 50424 3298 50488 3302
rect 50504 3358 50568 3362
rect 50504 3302 50508 3358
rect 50508 3302 50564 3358
rect 50564 3302 50568 3358
rect 50504 3298 50568 3302
rect 50584 3358 50648 3362
rect 50584 3302 50588 3358
rect 50588 3302 50644 3358
rect 50644 3302 50648 3358
rect 50584 3298 50648 3302
rect 4264 2692 4328 2696
rect 4264 2636 4268 2692
rect 4268 2636 4324 2692
rect 4324 2636 4328 2692
rect 4264 2632 4328 2636
rect 4344 2692 4408 2696
rect 4344 2636 4348 2692
rect 4348 2636 4404 2692
rect 4404 2636 4408 2692
rect 4344 2632 4408 2636
rect 4424 2692 4488 2696
rect 4424 2636 4428 2692
rect 4428 2636 4484 2692
rect 4484 2636 4488 2692
rect 4424 2632 4488 2636
rect 4504 2692 4568 2696
rect 4504 2636 4508 2692
rect 4508 2636 4564 2692
rect 4564 2636 4568 2692
rect 4504 2632 4568 2636
rect 34984 2692 35048 2696
rect 34984 2636 34988 2692
rect 34988 2636 35044 2692
rect 35044 2636 35048 2692
rect 34984 2632 35048 2636
rect 35064 2692 35128 2696
rect 35064 2636 35068 2692
rect 35068 2636 35124 2692
rect 35124 2636 35128 2692
rect 35064 2632 35128 2636
rect 35144 2692 35208 2696
rect 35144 2636 35148 2692
rect 35148 2636 35204 2692
rect 35204 2636 35208 2692
rect 35144 2632 35208 2636
rect 35224 2692 35288 2696
rect 35224 2636 35228 2692
rect 35228 2636 35284 2692
rect 35284 2636 35288 2692
rect 35224 2632 35288 2636
<< metal4 >>
rect 4256 57308 4576 57324
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 55976 4576 57244
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 54644 4576 55912
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 53312 4576 54580
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 51980 4576 53248
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 50648 4576 51916
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 49316 4576 50584
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 47984 4576 49252
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 46652 4576 47920
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 45320 4576 46588
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 43988 4576 45256
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 42656 4576 43924
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 41324 4576 42592
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 39992 4576 41260
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 38660 4576 39928
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 37328 4576 38596
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 35996 4576 37264
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 34664 4576 35932
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 33332 4576 34600
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 32000 4576 33268
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 30668 4576 31936
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 29336 4576 30604
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 28004 4576 29272
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 26672 4576 27940
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 25340 4576 26608
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 24008 4576 25276
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 22676 4576 23944
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 21344 4576 22612
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 20012 4576 21280
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 18680 4576 19948
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 17348 4576 18616
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 16016 4576 17284
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 14684 4576 15952
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 13352 4576 14620
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 12020 4576 13288
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 10688 4576 11956
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 9356 4576 10624
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 8024 4576 9292
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 6692 4576 7960
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 5360 4576 6628
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 4028 4576 5296
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 2696 4576 3964
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 56642 19936 57324
rect 34976 57308 35296 57324
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 55310 19936 56578
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 53978 19936 55246
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 52646 19936 53914
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 51314 19936 52582
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 49982 19936 51250
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 48650 19936 49918
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 47318 19936 48586
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 45986 19936 47254
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 44654 19936 45922
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 43322 19936 44590
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 41990 19936 43258
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 40658 19936 41926
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 39326 19936 40594
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 37994 19936 39262
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 36662 19936 37930
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 35330 19936 36598
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 33998 19936 35266
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 32666 19936 33934
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 31334 19936 32602
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 30002 19936 31270
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 28670 19936 29938
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 27338 19936 28606
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 26006 19936 27274
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 24674 19936 25942
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 23342 19936 24610
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 22010 19936 23278
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 20678 19936 21946
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 19346 19936 20614
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 18014 19936 19282
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 16682 19936 17950
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 15350 19936 16618
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 14018 19936 15286
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 12686 19936 13954
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 11354 19936 12622
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 10022 19936 11290
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 8690 19936 9958
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 7358 19936 8626
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 6026 19936 7294
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 4694 19936 5962
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 3362 19936 4630
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 4256 2616 4576 2632
rect 19616 2616 19936 3298
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 55976 35296 57244
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 54644 35296 55912
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 53312 35296 54580
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 51980 35296 53248
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 50648 35296 51916
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 49316 35296 50584
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 47984 35296 49252
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 46652 35296 47920
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 45320 35296 46588
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 43988 35296 45256
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 42656 35296 43924
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 41324 35296 42592
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 39992 35296 41260
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 38660 35296 39928
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 37328 35296 38596
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 35996 35296 37264
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 34664 35296 35932
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 33332 35296 34600
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 32000 35296 33268
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 30668 35296 31936
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 29336 35296 30604
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 28004 35296 29272
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 26672 35296 27940
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 25340 35296 26608
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 24008 35296 25276
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 22676 35296 23944
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 21344 35296 22612
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 20012 35296 21280
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 18680 35296 19948
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 17348 35296 18616
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 16016 35296 17284
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 14684 35296 15952
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 13352 35296 14620
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 12020 35296 13288
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 10688 35296 11956
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 9356 35296 10624
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 8024 35296 9292
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 6692 35296 7960
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 5360 35296 6628
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 4028 35296 5296
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 2696 35296 3964
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 56642 50656 57324
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 55310 50656 56578
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 53978 50656 55246
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 52646 50656 53914
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 51314 50656 52582
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 49982 50656 51250
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 48650 50656 49918
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 47318 50656 48586
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 45986 50656 47254
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 44654 50656 45922
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 43322 50656 44590
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 41990 50656 43258
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 40658 50656 41926
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 39326 50656 40594
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 37994 50656 39262
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 36662 50656 37930
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 35330 50656 36598
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 33998 50656 35266
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 32666 50656 33934
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 31334 50656 32602
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 30002 50656 31270
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 28670 50656 29938
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 27338 50656 28606
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 26006 50656 27274
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 24674 50656 25942
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 23342 50656 24610
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 22010 50656 23278
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 20678 50656 21946
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 19346 50656 20614
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 18014 50656 19282
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 16682 50656 17950
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 15350 50656 16618
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 14018 50656 15286
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 12686 50656 13954
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 11354 50656 12622
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 10022 50656 11290
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 8690 50656 9958
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 7358 50656 8626
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 6026 50656 7294
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 4694 50656 5962
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 3362 50656 4630
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 34976 2616 35296 2632
rect 50336 2616 50656 3298
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
use sky130_fd_sc_ls__decap_4  FILLER_1_8 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1920 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_8
timestamp 1621261055
transform 1 0 1920 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input296 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input295
timestamp 1621261055
transform 1 0 1536 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_2
timestamp 1621261055
transform 1 0 1152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_0
timestamp 1621261055
transform 1 0 1152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_16
timestamp 1621261055
transform 1 0 2688 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_16
timestamp 1621261055
transform 1 0 2688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input319
timestamp 1621261055
transform 1 0 2304 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input297
timestamp 1621261055
transform 1 0 2304 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_24
timestamp 1621261055
transform 1 0 3456 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_24
timestamp 1621261055
transform 1 0 3456 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input323
timestamp 1621261055
transform 1 0 3072 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input322
timestamp 1621261055
transform 1 0 3072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_32
timestamp 1621261055
transform 1 0 4224 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3936 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input324
timestamp 1621261055
transform 1 0 3840 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_164 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3840 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 4704 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input325
timestamp 1621261055
transform 1 0 4608 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_40
timestamp 1621261055
transform 1 0 4992 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input298
timestamp 1621261055
transform 1 0 4896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_44
timestamp 1621261055
transform 1 0 5376 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_43
timestamp 1621261055
transform 1 0 5280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input300
timestamp 1621261055
transform 1 0 5568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input299
timestamp 1621261055
transform 1 0 5664 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_50
timestamp 1621261055
transform 1 0 5952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_51
timestamp 1621261055
transform 1 0 6048 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_56
timestamp 1621261055
transform 1 0 6528 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 6336 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_57
timestamp 1621261055
transform 1 0 6624 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_55
timestamp 1621261055
transform 1 0 6432 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_185
timestamp 1621261055
transform 1 0 6432 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_165
timestamp 1621261055
transform 1 0 6528 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input302
timestamp 1621261055
transform 1 0 6912 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input301
timestamp 1621261055
transform 1 0 7008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_64
timestamp 1621261055
transform 1 0 7296 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_65
timestamp 1621261055
transform 1 0 7392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_72
timestamp 1621261055
transform 1 0 8064 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_73
timestamp 1621261055
transform 1 0 8160 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input304
timestamp 1621261055
transform 1 0 7680 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input303
timestamp 1621261055
transform 1 0 7776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_80
timestamp 1621261055
transform 1 0 8832 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_83
timestamp 1621261055
transform 1 0 9120 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_81
timestamp 1621261055
transform 1 0 8928 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input306
timestamp 1621261055
transform 1 0 8448 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_88
timestamp 1621261055
transform 1 0 9600 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_85
timestamp 1621261055
transform 1 0 9312 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input311
timestamp 1621261055
transform 1 0 9984 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input309
timestamp 1621261055
transform 1 0 9216 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input307
timestamp 1621261055
transform 1 0 9696 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_166
timestamp 1621261055
transform 1 0 9216 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_96
timestamp 1621261055
transform 1 0 10368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_93
timestamp 1621261055
transform 1 0 10080 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input310
timestamp 1621261055
transform 1 0 10464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_104
timestamp 1621261055
transform 1 0 11136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_101
timestamp 1621261055
transform 1 0 10848 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input313
timestamp 1621261055
transform 1 0 10752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_1_111
timestamp 1621261055
transform 1 0 11808 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_108
timestamp 1621261055
transform 1 0 11520 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_113
timestamp 1621261055
transform 1 0 12000 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_0_111
timestamp 1621261055
transform 1 0 11808 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_109
timestamp 1621261055
transform 1 0 11616 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_186
timestamp 1621261055
transform 1 0 11712 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_167
timestamp 1621261055
transform 1 0 11904 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_123
timestamp 1621261055
transform 1 0 12960 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_121
timestamp 1621261055
transform 1 0 12768 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input167
timestamp 1621261055
transform 1 0 12576 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input39 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 12960 0 -1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_1_132
timestamp 1621261055
transform 1 0 13824 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_128
timestamp 1621261055
transform 1 0 13440 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input100
timestamp 1621261055
transform 1 0 13824 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input78
timestamp 1621261055
transform 1 0 13344 0 1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_0_136
timestamp 1621261055
transform 1 0 14208 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input89
timestamp 1621261055
transform 1 0 14208 0 1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_168
timestamp 1621261055
transform 1 0 14592 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_149
timestamp 1621261055
transform 1 0 15456 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_141
timestamp 1621261055
transform 1 0 14688 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_141
timestamp 1621261055
transform 1 0 14688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input122
timestamp 1621261055
transform 1 0 15072 0 -1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_2  input111 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 15072 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_1_157
timestamp 1621261055
transform 1 0 16224 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_158
timestamp 1621261055
transform 1 0 16320 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_150
timestamp 1621261055
transform 1 0 15552 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input133
timestamp 1621261055
transform 1 0 15840 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_164
timestamp 1621261055
transform 1 0 16896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input50
timestamp 1621261055
transform 1 0 16512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_187
timestamp 1621261055
transform 1 0 16992 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_166
timestamp 1621261055
transform 1 0 17088 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_169
timestamp 1621261055
transform 1 0 17376 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input70
timestamp 1621261055
transform 1 0 17472 0 1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input61
timestamp 1621261055
transform 1 0 17760 0 -1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_169
timestamp 1621261055
transform 1 0 17280 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_175
timestamp 1621261055
transform 1 0 17952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_178
timestamp 1621261055
transform 1 0 18240 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input72
timestamp 1621261055
transform 1 0 18336 0 1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input71
timestamp 1621261055
transform 1 0 18624 0 -1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_1_184
timestamp 1621261055
transform 1 0 18816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_187
timestamp 1621261055
transform 1 0 19104 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input73
timestamp 1621261055
transform 1 0 19200 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_198
timestamp 1621261055
transform 1 0 20160 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_196
timestamp 1621261055
transform 1 0 19968 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_192
timestamp 1621261055
transform 1 0 19584 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_197
timestamp 1621261055
transform 1 0 20064 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_195
timestamp 1621261055
transform 1 0 19872 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_170
timestamp 1621261055
transform 1 0 19968 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_204
timestamp 1621261055
transform 1 0 20736 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_206
timestamp 1621261055
transform 1 0 20928 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input79
timestamp 1621261055
transform 1 0 20256 0 1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input77
timestamp 1621261055
transform 1 0 20448 0 -1 3330
box -38 -49 518 715
use sky130_fd_sc_ls__decap_8  FILLER_1_212
timestamp 1621261055
transform 1 0 21504 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_0_214
timestamp 1621261055
transform 1 0 21696 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input80
timestamp 1621261055
transform 1 0 21120 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input75 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 21312 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_221
timestamp 1621261055
transform 1 0 22368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_222
timestamp 1621261055
transform 1 0 22464 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_188
timestamp 1621261055
transform 1 0 22272 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_171
timestamp 1621261055
transform 1 0 22656 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_229
timestamp 1621261055
transform 1 0 23136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_225
timestamp 1621261055
transform 1 0 22752 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input84
timestamp 1621261055
transform 1 0 22752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input82
timestamp 1621261055
transform 1 0 23136 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_233
timestamp 1621261055
transform 1 0 23520 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input86
timestamp 1621261055
transform 1 0 23520 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_237
timestamp 1621261055
transform 1 0 23904 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input85
timestamp 1621261055
transform 1 0 23904 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_245
timestamp 1621261055
transform 1 0 24672 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_241
timestamp 1621261055
transform 1 0 24288 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input88
timestamp 1621261055
transform 1 0 24288 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _158_ $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 24672 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_248
timestamp 1621261055
transform 1 0 24960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input91
timestamp 1621261055
transform 1 0 25056 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_253
timestamp 1621261055
transform 1 0 25440 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_253
timestamp 1621261055
transform 1 0 25440 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_172
timestamp 1621261055
transform 1 0 25344 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input92
timestamp 1621261055
transform 1 0 25824 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input90
timestamp 1621261055
transform 1 0 25824 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_261
timestamp 1621261055
transform 1 0 26208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_261
timestamp 1621261055
transform 1 0 26208 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_269
timestamp 1621261055
transform 1 0 26976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_269
timestamp 1621261055
transform 1 0 26976 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input95
timestamp 1621261055
transform 1 0 26592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input93
timestamp 1621261055
transform 1 0 26592 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_276
timestamp 1621261055
transform 1 0 27648 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_273
timestamp 1621261055
transform 1 0 27360 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_281
timestamp 1621261055
transform 1 0 28128 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_279
timestamp 1621261055
transform 1 0 27936 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_277
timestamp 1621261055
transform 1 0 27744 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input99
timestamp 1621261055
transform 1 0 28032 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_189
timestamp 1621261055
transform 1 0 27552 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_173
timestamp 1621261055
transform 1 0 28032 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_284
timestamp 1621261055
transform 1 0 28416 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_289
timestamp 1621261055
transform 1 0 28896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input102
timestamp 1621261055
transform 1 0 28800 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input98
timestamp 1621261055
transform 1 0 28512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_292
timestamp 1621261055
transform 1 0 29184 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_297
timestamp 1621261055
transform 1 0 29664 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input104
timestamp 1621261055
transform 1 0 29568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input101
timestamp 1621261055
transform 1 0 29280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_300
timestamp 1621261055
transform 1 0 29952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_305
timestamp 1621261055
transform 1 0 30432 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input106
timestamp 1621261055
transform 1 0 30336 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_308
timestamp 1621261055
transform 1 0 30720 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_309
timestamp 1621261055
transform 1 0 30816 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_307
timestamp 1621261055
transform 1 0 30624 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input108
timestamp 1621261055
transform 1 0 31104 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input107
timestamp 1621261055
transform 1 0 31200 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_174
timestamp 1621261055
transform 1 0 30720 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_316
timestamp 1621261055
transform 1 0 31488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_317
timestamp 1621261055
transform 1 0 31584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input112
timestamp 1621261055
transform 1 0 31872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input109
timestamp 1621261055
transform 1 0 31968 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_328
timestamp 1621261055
transform 1 0 32640 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_324
timestamp 1621261055
transform 1 0 32256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_325
timestamp 1621261055
transform 1 0 32352 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_190
timestamp 1621261055
transform 1 0 32832 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_331
timestamp 1621261055
transform 1 0 32928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_337
timestamp 1621261055
transform 1 0 33504 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_335
timestamp 1621261055
transform 1 0 33312 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_333
timestamp 1621261055
transform 1 0 33120 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input115
timestamp 1621261055
transform 1 0 33312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_175
timestamp 1621261055
transform 1 0 33408 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_347
timestamp 1621261055
transform 1 0 34464 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_339
timestamp 1621261055
transform 1 0 33696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_345
timestamp 1621261055
transform 1 0 34272 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input118
timestamp 1621261055
transform 1 0 34080 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input114
timestamp 1621261055
transform 1 0 33888 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_355
timestamp 1621261055
transform 1 0 35232 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_353
timestamp 1621261055
transform 1 0 35040 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input120
timestamp 1621261055
transform 1 0 34848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input117
timestamp 1621261055
transform 1 0 34656 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_363
timestamp 1621261055
transform 1 0 36000 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_363
timestamp 1621261055
transform 1 0 36000 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_361
timestamp 1621261055
transform 1 0 35808 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input123
timestamp 1621261055
transform 1 0 35616 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_371
timestamp 1621261055
transform 1 0 36768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_365
timestamp 1621261055
transform 1 0 36192 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input125
timestamp 1621261055
transform 1 0 36384 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input124
timestamp 1621261055
transform 1 0 36576 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_176
timestamp 1621261055
transform 1 0 36096 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_379
timestamp 1621261055
transform 1 0 37536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_373
timestamp 1621261055
transform 1 0 36960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input127
timestamp 1621261055
transform 1 0 37152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input126
timestamp 1621261055
transform 1 0 37344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_386
timestamp 1621261055
transform 1 0 38208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_383
timestamp 1621261055
transform 1 0 37920 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_389
timestamp 1621261055
transform 1 0 38496 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_381
timestamp 1621261055
transform 1 0 37728 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_191
timestamp 1621261055
transform 1 0 38112 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_394
timestamp 1621261055
transform 1 0 38976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_393
timestamp 1621261055
transform 1 0 38880 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_391
timestamp 1621261055
transform 1 0 38688 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input131
timestamp 1621261055
transform 1 0 38592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_177
timestamp 1621261055
transform 1 0 38784 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_402
timestamp 1621261055
transform 1 0 39744 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_401
timestamp 1621261055
transform 1 0 39648 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input134
timestamp 1621261055
transform 1 0 39360 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input130
timestamp 1621261055
transform 1 0 39264 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_410
timestamp 1621261055
transform 1 0 40512 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_409
timestamp 1621261055
transform 1 0 40416 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input136
timestamp 1621261055
transform 1 0 40128 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input132
timestamp 1621261055
transform 1 0 40032 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_418
timestamp 1621261055
transform 1 0 41280 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_421
timestamp 1621261055
transform 1 0 41568 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_419
timestamp 1621261055
transform 1 0 41376 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_417
timestamp 1621261055
transform 1 0 41184 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input140
timestamp 1621261055
transform 1 0 41664 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input138
timestamp 1621261055
transform 1 0 40896 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_178
timestamp 1621261055
transform 1 0 41472 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_426
timestamp 1621261055
transform 1 0 42048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_429
timestamp 1621261055
transform 1 0 42336 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input139
timestamp 1621261055
transform 1 0 41952 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_434
timestamp 1621261055
transform 1 0 42816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_437
timestamp 1621261055
transform 1 0 43104 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input142
timestamp 1621261055
transform 1 0 42432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input141
timestamp 1621261055
transform 1 0 42720 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_441
timestamp 1621261055
transform 1 0 43488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_438
timestamp 1621261055
transform 1 0 43200 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_445
timestamp 1621261055
transform 1 0 43872 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input146
timestamp 1621261055
transform 1 0 43872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_192
timestamp 1621261055
transform 1 0 43392 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_449
timestamp 1621261055
transform 1 0 44256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_449
timestamp 1621261055
transform 1 0 44256 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_447
timestamp 1621261055
transform 1 0 44064 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input149
timestamp 1621261055
transform 1 0 44640 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input147
timestamp 1621261055
transform 1 0 44640 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_179
timestamp 1621261055
transform 1 0 44160 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_457
timestamp 1621261055
transform 1 0 45024 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_457
timestamp 1621261055
transform 1 0 45024 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input151
timestamp 1621261055
transform 1 0 45408 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input150
timestamp 1621261055
transform 1 0 45408 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_465
timestamp 1621261055
transform 1 0 45792 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_465
timestamp 1621261055
transform 1 0 45792 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input153
timestamp 1621261055
transform 1 0 46176 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _108_
timestamp 1621261055
transform 1 0 46176 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_473
timestamp 1621261055
transform 1 0 46560 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_477
timestamp 1621261055
transform 1 0 46944 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_472
timestamp 1621261055
transform 1 0 46464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input156
timestamp 1621261055
transform 1 0 46944 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_180
timestamp 1621261055
transform 1 0 46848 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_481
timestamp 1621261055
transform 1 0 47328 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_485
timestamp 1621261055
transform 1 0 47712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input159
timestamp 1621261055
transform 1 0 47712 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input154
timestamp 1621261055
transform 1 0 47328 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_493
timestamp 1621261055
transform 1 0 48480 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_489
timestamp 1621261055
transform 1 0 48096 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_493
timestamp 1621261055
transform 1 0 48480 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input157
timestamp 1621261055
transform 1 0 48096 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_193
timestamp 1621261055
transform 1 0 48672 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_496
timestamp 1621261055
transform 1 0 48768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_503
timestamp 1621261055
transform 1 0 49440 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_501
timestamp 1621261055
transform 1 0 49248 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input162
timestamp 1621261055
transform 1 0 49152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_512
timestamp 1621261055
transform 1 0 50304 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_504
timestamp 1621261055
transform 1 0 49536 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_505
timestamp 1621261055
transform 1 0 49632 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input40
timestamp 1621261055
transform 1 0 50016 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_181
timestamp 1621261055
transform 1 0 49536 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_517
timestamp 1621261055
transform 1 0 50784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_521
timestamp 1621261055
transform 1 0 51168 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_513
timestamp 1621261055
transform 1 0 50400 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input43
timestamp 1621261055
transform 1 0 51168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input42
timestamp 1621261055
transform 1 0 50400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input41
timestamp 1621261055
transform 1 0 50784 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_525
timestamp 1621261055
transform 1 0 51552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_528
timestamp 1621261055
transform 1 0 51840 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_16 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform -1 0 51552 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _214_
timestamp 1621261055
transform -1 0 51840 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_533
timestamp 1621261055
transform 1 0 52320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_533
timestamp 1621261055
transform 1 0 52320 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input44
timestamp 1621261055
transform 1 0 51936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_182
timestamp 1621261055
transform 1 0 52224 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_541
timestamp 1621261055
transform 1 0 53088 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_541
timestamp 1621261055
transform 1 0 53088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input47
timestamp 1621261055
transform 1 0 53472 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input46
timestamp 1621261055
transform 1 0 52704 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input45
timestamp 1621261055
transform 1 0 52704 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_551
timestamp 1621261055
transform 1 0 54048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_549
timestamp 1621261055
transform 1 0 53856 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_549
timestamp 1621261055
transform 1 0 53856 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_194
timestamp 1621261055
transform 1 0 53952 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _110_
timestamp 1621261055
transform 1 0 54240 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_559
timestamp 1621261055
transform 1 0 54816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_561
timestamp 1621261055
transform 1 0 55008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_556
timestamp 1621261055
transform 1 0 54528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input51
timestamp 1621261055
transform 1 0 54432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_183
timestamp 1621261055
transform 1 0 54912 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_567
timestamp 1621261055
transform 1 0 55584 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_569
timestamp 1621261055
transform 1 0 55776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input54
timestamp 1621261055
transform 1 0 55200 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input52
timestamp 1621261055
transform 1 0 55392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_575
timestamp 1621261055
transform 1 0 56352 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_577
timestamp 1621261055
transform 1 0 56544 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input56
timestamp 1621261055
transform 1 0 55968 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input55
timestamp 1621261055
transform 1 0 56160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_583
timestamp 1621261055
transform 1 0 57120 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_584
timestamp 1621261055
transform 1 0 57216 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input59
timestamp 1621261055
transform 1 0 57504 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input58
timestamp 1621261055
transform 1 0 56736 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _109_
timestamp 1621261055
transform 1 0 56928 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_591
timestamp 1621261055
transform 1 0 57888 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_589
timestamp 1621261055
transform 1 0 57696 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_184
timestamp 1621261055
transform 1 0 57600 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_1
timestamp 1621261055
transform -1 0 58848 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_3
timestamp 1621261055
transform -1 0 58848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_595
timestamp 1621261055
transform 1 0 58272 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input308
timestamp 1621261055
transform 1 0 1536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_4
timestamp 1621261055
transform 1 0 1152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_8
timestamp 1621261055
transform 1 0 1920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input330
timestamp 1621261055
transform 1 0 2304 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_16
timestamp 1621261055
transform 1 0 2688 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_24
timestamp 1621261055
transform 1 0 3456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input341
timestamp 1621261055
transform 1 0 3072 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_195
timestamp 1621261055
transform 1 0 3840 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_29
timestamp 1621261055
transform 1 0 3936 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input326
timestamp 1621261055
transform 1 0 4320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input305
timestamp 1621261055
transform 1 0 7392 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input328
timestamp 1621261055
transform 1 0 5088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input331
timestamp 1621261055
transform 1 0 5856 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input333
timestamp 1621261055
transform 1 0 6624 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_37
timestamp 1621261055
transform 1 0 4704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_45
timestamp 1621261055
transform 1 0 5472 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_53
timestamp 1621261055
transform 1 0 6240 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_61
timestamp 1621261055
transform 1 0 7008 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_196
timestamp 1621261055
transform 1 0 9120 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input312
timestamp 1621261055
transform 1 0 9600 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input314
timestamp 1621261055
transform 1 0 10368 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input335
timestamp 1621261055
transform 1 0 8160 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_69
timestamp 1621261055
transform 1 0 7776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_77
timestamp 1621261055
transform 1 0 8544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_81
timestamp 1621261055
transform 1 0 8928 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_84
timestamp 1621261055
transform 1 0 9216 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_92
timestamp 1621261055
transform 1 0 9984 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input206
timestamp 1621261055
transform 1 0 13536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input315
timestamp 1621261055
transform 1 0 11136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input316
timestamp 1621261055
transform 1 0 11904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input317
timestamp 1621261055
transform 1 0 12672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_100
timestamp 1621261055
transform 1 0 10752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_108
timestamp 1621261055
transform 1 0 11520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_116
timestamp 1621261055
transform 1 0 12288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_124
timestamp 1621261055
transform 1 0 13056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_128
timestamp 1621261055
transform 1 0 13440 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_139
timestamp 1621261055
transform 1 0 14496 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_2_137
timestamp 1621261055
transform 1 0 14304 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_133
timestamp 1621261055
transform 1 0 13920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_197
timestamp 1621261055
transform 1 0 14400 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_147
timestamp 1621261055
transform 1 0 15264 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input144
timestamp 1621261055
transform 1 0 15456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_153
timestamp 1621261055
transform 1 0 15840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input155
timestamp 1621261055
transform 1 0 16224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_161
timestamp 1621261055
transform 1 0 16608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input166
timestamp 1621261055
transform 1 0 16992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_169
timestamp 1621261055
transform 1 0 17376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input178
timestamp 1621261055
transform 1 0 17760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_177
timestamp 1621261055
transform 1 0 18144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_183
timestamp 1621261055
transform 1 0 18720 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_181
timestamp 1621261055
transform 1 0 18528 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input74
timestamp 1621261055
transform 1 0 18816 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_188
timestamp 1621261055
transform 1 0 19200 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_192
timestamp 1621261055
transform 1 0 19584 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_198
timestamp 1621261055
transform 1 0 19680 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_194
timestamp 1621261055
transform 1 0 19776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input76
timestamp 1621261055
transform 1 0 20160 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _119_
timestamp 1621261055
transform 1 0 22560 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input81
timestamp 1621261055
transform 1 0 21024 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input83
timestamp 1621261055
transform 1 0 21792 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input87
timestamp 1621261055
transform 1 0 23232 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_202
timestamp 1621261055
transform 1 0 20544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_206
timestamp 1621261055
transform 1 0 20928 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_211
timestamp 1621261055
transform 1 0 21408 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_219
timestamp 1621261055
transform 1 0 22176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_226
timestamp 1621261055
transform 1 0 22848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_199
timestamp 1621261055
transform 1 0 24960 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input94
timestamp 1621261055
transform 1 0 25440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input96
timestamp 1621261055
transform 1 0 26208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input211
timestamp 1621261055
transform 1 0 24000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_234
timestamp 1621261055
transform 1 0 23616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_242
timestamp 1621261055
transform 1 0 24384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_246
timestamp 1621261055
transform 1 0 24768 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_249
timestamp 1621261055
transform 1 0 25056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_257
timestamp 1621261055
transform 1 0 25824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input97
timestamp 1621261055
transform 1 0 26976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input103
timestamp 1621261055
transform 1 0 28320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input105
timestamp 1621261055
transform 1 0 29088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_265
timestamp 1621261055
transform 1 0 26592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_273
timestamp 1621261055
transform 1 0 27360 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_281
timestamp 1621261055
transform 1 0 28128 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_287
timestamp 1621261055
transform 1 0 28704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_295
timestamp 1621261055
transform 1 0 29472 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_304
timestamp 1621261055
transform 1 0 30336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_200
timestamp 1621261055
transform 1 0 30240 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_308
timestamp 1621261055
transform 1 0 30720 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input110
timestamp 1621261055
transform 1 0 30912 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_314
timestamp 1621261055
transform 1 0 31296 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input113
timestamp 1621261055
transform 1 0 31680 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_322
timestamp 1621261055
transform 1 0 32064 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_328
timestamp 1621261055
transform 1 0 32640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_326
timestamp 1621261055
transform 1 0 32448 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input116
timestamp 1621261055
transform 1 0 32736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_201
timestamp 1621261055
transform 1 0 35520 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input119
timestamp 1621261055
transform 1 0 33888 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input121
timestamp 1621261055
transform 1 0 34656 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input247
timestamp 1621261055
transform 1 0 36000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_333
timestamp 1621261055
transform 1 0 33120 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_345
timestamp 1621261055
transform 1 0 34272 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_353
timestamp 1621261055
transform 1 0 35040 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_357
timestamp 1621261055
transform 1 0 35424 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_359
timestamp 1621261055
transform 1 0 35616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _005_
timestamp 1621261055
transform 1 0 38304 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input128
timestamp 1621261055
transform 1 0 36768 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input129
timestamp 1621261055
transform 1 0 37536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input135
timestamp 1621261055
transform 1 0 38976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_6
timestamp 1621261055
transform 1 0 38112 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_367
timestamp 1621261055
transform 1 0 36384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_375
timestamp 1621261055
transform 1 0 37152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_383
timestamp 1621261055
transform 1 0 37920 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_390
timestamp 1621261055
transform 1 0 38592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_398
timestamp 1621261055
transform 1 0 39360 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input137
timestamp 1621261055
transform 1 0 39744 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_410
timestamp 1621261055
transform 1 0 40512 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_406
timestamp 1621261055
transform 1 0 40128 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_414
timestamp 1621261055
transform 1 0 40896 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_412
timestamp 1621261055
transform 1 0 40704 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_202
timestamp 1621261055
transform 1 0 40800 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _060_
timestamp 1621261055
transform 1 0 41280 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_2_421
timestamp 1621261055
transform 1 0 41568 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_429
timestamp 1621261055
transform 1 0 42336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input143
timestamp 1621261055
transform 1 0 41952 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input145
timestamp 1621261055
transform 1 0 42720 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input148
timestamp 1621261055
transform 1 0 43488 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input152
timestamp 1621261055
transform 1 0 44928 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_437
timestamp 1621261055
transform 1 0 43104 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_445
timestamp 1621261055
transform 1 0 43872 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_453
timestamp 1621261055
transform 1 0 44640 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_455
timestamp 1621261055
transform 1 0 44832 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_460
timestamp 1621261055
transform 1 0 45312 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_203
timestamp 1621261055
transform 1 0 46080 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input158
timestamp 1621261055
transform 1 0 46752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input160
timestamp 1621261055
transform 1 0 47520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input161
timestamp 1621261055
transform 1 0 48288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_469
timestamp 1621261055
transform 1 0 46176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_473
timestamp 1621261055
transform 1 0 46560 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_479
timestamp 1621261055
transform 1 0 47136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_487
timestamp 1621261055
transform 1 0 47904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_495
timestamp 1621261055
transform 1 0 48672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_204
timestamp 1621261055
transform 1 0 51360 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input163
timestamp 1621261055
transform 1 0 49056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input164
timestamp 1621261055
transform 1 0 49824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input168
timestamp 1621261055
transform 1 0 50592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input171
timestamp 1621261055
transform 1 0 51840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_503
timestamp 1621261055
transform 1 0 49440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_511
timestamp 1621261055
transform 1 0 50208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_519
timestamp 1621261055
transform 1 0 50976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_524
timestamp 1621261055
transform 1 0 51456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _165_
timestamp 1621261055
transform 1 0 54912 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input48
timestamp 1621261055
transform 1 0 52608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input49
timestamp 1621261055
transform 1 0 53376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input53
timestamp 1621261055
transform 1 0 54144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_532
timestamp 1621261055
transform 1 0 52224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_540
timestamp 1621261055
transform 1 0 52992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_548
timestamp 1621261055
transform 1 0 53760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_556
timestamp 1621261055
transform 1 0 54528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_205
timestamp 1621261055
transform 1 0 56640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input57
timestamp 1621261055
transform 1 0 55584 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input60
timestamp 1621261055
transform 1 0 57120 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_563
timestamp 1621261055
transform 1 0 55200 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_571
timestamp 1621261055
transform 1 0 55968 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_575
timestamp 1621261055
transform 1 0 56352 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_577
timestamp 1621261055
transform 1 0 56544 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_579
timestamp 1621261055
transform 1 0 56736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_587
timestamp 1621261055
transform 1 0 57504 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_5
timestamp 1621261055
transform -1 0 58848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_595
timestamp 1621261055
transform 1 0 58272 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input329
timestamp 1621261055
transform 1 0 1536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_6
timestamp 1621261055
transform 1 0 1152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_8
timestamp 1621261055
transform 1 0 1920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input352
timestamp 1621261055
transform 1 0 2304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_16
timestamp 1621261055
transform 1 0 2688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_24
timestamp 1621261055
transform 1 0 3456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input355
timestamp 1621261055
transform 1 0 3072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_28
timestamp 1621261055
transform 1 0 3840 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_30
timestamp 1621261055
transform 1 0 4032 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input327
timestamp 1621261055
transform 1 0 4128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_35
timestamp 1621261055
transform 1 0 4512 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_3_48
timestamp 1621261055
transform 1 0 5760 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_43
timestamp 1621261055
transform 1 0 5280 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input332
timestamp 1621261055
transform 1 0 5376 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_56
timestamp 1621261055
transform 1 0 6528 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_54
timestamp 1621261055
transform 1 0 6336 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_52
timestamp 1621261055
transform 1 0 6144 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_206
timestamp 1621261055
transform 1 0 6432 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_64
timestamp 1621261055
transform 1 0 7296 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input334
timestamp 1621261055
transform 1 0 6912 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input336
timestamp 1621261055
transform 1 0 7680 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input338
timestamp 1621261055
transform 1 0 8448 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input340
timestamp 1621261055
transform 1 0 9216 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input342
timestamp 1621261055
transform 1 0 9984 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_72
timestamp 1621261055
transform 1 0 8064 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_80
timestamp 1621261055
transform 1 0 8832 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_88
timestamp 1621261055
transform 1 0 9600 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_96
timestamp 1621261055
transform 1 0 10368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input344
timestamp 1621261055
transform 1 0 10752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_108
timestamp 1621261055
transform 1 0 11520 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_104
timestamp 1621261055
transform 1 0 11136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_111
timestamp 1621261055
transform 1 0 11808 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_207
timestamp 1621261055
transform 1 0 11712 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input318
timestamp 1621261055
transform 1 0 12192 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_119
timestamp 1621261055
transform 1 0 12576 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input320
timestamp 1621261055
transform 1 0 12960 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_127
timestamp 1621261055
transform 1 0 13344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_131
timestamp 1621261055
transform 1 0 13728 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_208
timestamp 1621261055
transform 1 0 16992 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input217
timestamp 1621261055
transform 1 0 13920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input228
timestamp 1621261055
transform 1 0 14688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input239
timestamp 1621261055
transform 1 0 15456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input261
timestamp 1621261055
transform 1 0 16224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_137
timestamp 1621261055
transform 1 0 14304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_145
timestamp 1621261055
transform 1 0 15072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_153
timestamp 1621261055
transform 1 0 15840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_161
timestamp 1621261055
transform 1 0 16608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input189
timestamp 1621261055
transform 1 0 17472 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input198
timestamp 1621261055
transform 1 0 18240 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input200
timestamp 1621261055
transform 1 0 19008 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input202
timestamp 1621261055
transform 1 0 19776 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_166
timestamp 1621261055
transform 1 0 17088 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_174
timestamp 1621261055
transform 1 0 17856 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_182
timestamp 1621261055
transform 1 0 18624 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_190
timestamp 1621261055
transform 1 0 19392 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_198
timestamp 1621261055
transform 1 0 20160 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_209
timestamp 1621261055
transform 1 0 22272 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input203
timestamp 1621261055
transform 1 0 20544 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input205
timestamp 1621261055
transform 1 0 21312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input209
timestamp 1621261055
transform 1 0 22752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_206
timestamp 1621261055
transform 1 0 20928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_214
timestamp 1621261055
transform 1 0 21696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_218
timestamp 1621261055
transform 1 0 22080 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_221
timestamp 1621261055
transform 1 0 22368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_229
timestamp 1621261055
transform 1 0 23136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input212
timestamp 1621261055
transform 1 0 23520 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input214
timestamp 1621261055
transform 1 0 24288 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input216
timestamp 1621261055
transform 1 0 25056 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input218
timestamp 1621261055
transform 1 0 25824 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_237
timestamp 1621261055
transform 1 0 23904 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_245
timestamp 1621261055
transform 1 0 24672 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_253
timestamp 1621261055
transform 1 0 25440 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_261
timestamp 1621261055
transform 1 0 26208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input220
timestamp 1621261055
transform 1 0 26592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_273
timestamp 1621261055
transform 1 0 27360 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_269
timestamp 1621261055
transform 1 0 26976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_276
timestamp 1621261055
transform 1 0 27648 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_210
timestamp 1621261055
transform 1 0 27552 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input224
timestamp 1621261055
transform 1 0 28032 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_284
timestamp 1621261055
transform 1 0 28416 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input227
timestamp 1621261055
transform 1 0 28800 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_292
timestamp 1621261055
transform 1 0 29184 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input230
timestamp 1621261055
transform 1 0 29568 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_211
timestamp 1621261055
transform 1 0 32832 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input232
timestamp 1621261055
transform 1 0 30336 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input233
timestamp 1621261055
transform 1 0 31104 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input236
timestamp 1621261055
transform 1 0 31872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_300
timestamp 1621261055
transform 1 0 29952 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_308
timestamp 1621261055
transform 1 0 30720 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_316
timestamp 1621261055
transform 1 0 31488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_324
timestamp 1621261055
transform 1 0 32256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_328
timestamp 1621261055
transform 1 0 32640 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input241
timestamp 1621261055
transform 1 0 33312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input243
timestamp 1621261055
transform 1 0 34080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input245
timestamp 1621261055
transform 1 0 34848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input248
timestamp 1621261055
transform 1 0 35616 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_331
timestamp 1621261055
transform 1 0 32928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_339
timestamp 1621261055
transform 1 0 33696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_347
timestamp 1621261055
transform 1 0 34464 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_355
timestamp 1621261055
transform 1 0 35232 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_363
timestamp 1621261055
transform 1 0 36000 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_212
timestamp 1621261055
transform 1 0 38112 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input249
timestamp 1621261055
transform 1 0 36384 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input252
timestamp 1621261055
transform 1 0 37152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input256
timestamp 1621261055
transform 1 0 38592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_371
timestamp 1621261055
transform 1 0 36768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_379
timestamp 1621261055
transform 1 0 37536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_383
timestamp 1621261055
transform 1 0 37920 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_386
timestamp 1621261055
transform 1 0 38208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_394
timestamp 1621261055
transform 1 0 38976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input258
timestamp 1621261055
transform 1 0 39360 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input260
timestamp 1621261055
transform 1 0 40128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input264
timestamp 1621261055
transform 1 0 40896 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input265
timestamp 1621261055
transform 1 0 41664 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_402
timestamp 1621261055
transform 1 0 39744 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_410
timestamp 1621261055
transform 1 0 40512 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_418
timestamp 1621261055
transform 1 0 41280 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_426
timestamp 1621261055
transform 1 0 42048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input268
timestamp 1621261055
transform 1 0 42432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_438
timestamp 1621261055
transform 1 0 43200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_434
timestamp 1621261055
transform 1 0 42816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_441
timestamp 1621261055
transform 1 0 43488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_213
timestamp 1621261055
transform 1 0 43392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input271
timestamp 1621261055
transform 1 0 43872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_449
timestamp 1621261055
transform 1 0 44256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input274
timestamp 1621261055
transform 1 0 44640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_457
timestamp 1621261055
transform 1 0 45024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input276
timestamp 1621261055
transform 1 0 45408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_214
timestamp 1621261055
transform 1 0 48672 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input278
timestamp 1621261055
transform 1 0 46176 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input280
timestamp 1621261055
transform 1 0 46944 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input284
timestamp 1621261055
transform 1 0 47712 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_465
timestamp 1621261055
transform 1 0 45792 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_473
timestamp 1621261055
transform 1 0 46560 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_481
timestamp 1621261055
transform 1 0 47328 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_489
timestamp 1621261055
transform 1 0 48096 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_493
timestamp 1621261055
transform 1 0 48480 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_496
timestamp 1621261055
transform 1 0 48768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_500
timestamp 1621261055
transform 1 0 49152 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input165
timestamp 1621261055
transform 1 0 49344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_506
timestamp 1621261055
transform 1 0 49728 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_510
timestamp 1621261055
transform 1 0 50112 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input169
timestamp 1621261055
transform 1 0 50304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_516
timestamp 1621261055
transform 1 0 50688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input170
timestamp 1621261055
transform 1 0 51072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_524
timestamp 1621261055
transform 1 0 51456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input172
timestamp 1621261055
transform 1 0 51840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_215
timestamp 1621261055
transform 1 0 53952 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input173
timestamp 1621261055
transform 1 0 52608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input177
timestamp 1621261055
transform 1 0 54432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_532
timestamp 1621261055
transform 1 0 52224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_540
timestamp 1621261055
transform 1 0 52992 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_548
timestamp 1621261055
transform 1 0 53760 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_551
timestamp 1621261055
transform 1 0 54048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_559
timestamp 1621261055
transform 1 0 54816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_565
timestamp 1621261055
transform 1 0 55392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_563
timestamp 1621261055
transform 1 0 55200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_570
timestamp 1621261055
transform 1 0 55872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input68
timestamp 1621261055
transform 1 0 55488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input64
timestamp 1621261055
transform 1 0 56256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_578
timestamp 1621261055
transform 1 0 56640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input62
timestamp 1621261055
transform 1 0 57024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_586
timestamp 1621261055
transform 1 0 57408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_593
timestamp 1621261055
transform 1 0 58080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _197_
timestamp 1621261055
transform 1 0 57792 0 1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_7
timestamp 1621261055
transform -1 0 58848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_8
timestamp 1621261055
transform 1 0 1920 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input362
timestamp 1621261055
transform 1 0 1536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_8
timestamp 1621261055
transform 1 0 1152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_16
timestamp 1621261055
transform 1 0 2688 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input356
timestamp 1621261055
transform 1 0 2784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_25
timestamp 1621261055
transform 1 0 3552 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_21
timestamp 1621261055
transform 1 0 3168 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_29
timestamp 1621261055
transform 1 0 3936 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_27
timestamp 1621261055
transform 1 0 3744 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input358
timestamp 1621261055
transform 1 0 4320 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_216
timestamp 1621261055
transform 1 0 3840 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input337
timestamp 1621261055
transform 1 0 7200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input360
timestamp 1621261055
transform 1 0 5088 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output574
timestamp 1621261055
transform 1 0 5856 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_37
timestamp 1621261055
transform 1 0 4704 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_45
timestamp 1621261055
transform 1 0 5472 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_53
timestamp 1621261055
transform 1 0 6240 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_61
timestamp 1621261055
transform 1 0 7008 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_217
timestamp 1621261055
transform 1 0 9120 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input339
timestamp 1621261055
transform 1 0 7968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input343
timestamp 1621261055
transform 1 0 9600 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input345
timestamp 1621261055
transform 1 0 10368 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_67
timestamp 1621261055
transform 1 0 7584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_75
timestamp 1621261055
transform 1 0 8352 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_4_84
timestamp 1621261055
transform 1 0 9216 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_92
timestamp 1621261055
transform 1 0 9984 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_100
timestamp 1621261055
transform 1 0 10752 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_108
timestamp 1621261055
transform 1 0 11520 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input347
timestamp 1621261055
transform 1 0 11136 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_57
timestamp 1621261055
transform 1 0 11712 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _053_
timestamp 1621261055
transform 1 0 11904 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_4_115
timestamp 1621261055
transform 1 0 12192 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_123
timestamp 1621261055
transform 1 0 12960 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input321
timestamp 1621261055
transform 1 0 12576 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input351
timestamp 1621261055
transform 1 0 13344 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_131
timestamp 1621261055
transform 1 0 13728 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_135
timestamp 1621261055
transform 1 0 14112 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_139
timestamp 1621261055
transform 1 0 14496 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_137
timestamp 1621261055
transform 1 0 14304 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_218
timestamp 1621261055
transform 1 0 14400 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_4_143
timestamp 1621261055
transform 1 0 14880 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input250
timestamp 1621261055
transform 1 0 14976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_148
timestamp 1621261055
transform 1 0 15360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_156
timestamp 1621261055
transform 1 0 16128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input272
timestamp 1621261055
transform 1 0 15744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input283
timestamp 1621261055
transform 1 0 16512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_164
timestamp 1621261055
transform 1 0 16896 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_42
timestamp 1621261055
transform 1 0 17088 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _047_
timestamp 1621261055
transform 1 0 17280 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_4_171
timestamp 1621261055
transform 1 0 17568 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_179
timestamp 1621261055
transform 1 0 18336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input199
timestamp 1621261055
transform 1 0 17952 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input201
timestamp 1621261055
transform 1 0 18720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_187
timestamp 1621261055
transform 1 0 19104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_191
timestamp 1621261055
transform 1 0 19488 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_219
timestamp 1621261055
transform 1 0 19680 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_194
timestamp 1621261055
transform 1 0 19776 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input204
timestamp 1621261055
transform 1 0 20160 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input207
timestamp 1621261055
transform 1 0 20928 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input208
timestamp 1621261055
transform 1 0 21696 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input210
timestamp 1621261055
transform 1 0 22464 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input213
timestamp 1621261055
transform 1 0 23232 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_202
timestamp 1621261055
transform 1 0 20544 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_210
timestamp 1621261055
transform 1 0 21312 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_218
timestamp 1621261055
transform 1 0 22080 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_226
timestamp 1621261055
transform 1 0 22848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_220
timestamp 1621261055
transform 1 0 24960 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input215
timestamp 1621261055
transform 1 0 24000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input219
timestamp 1621261055
transform 1 0 25440 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input221
timestamp 1621261055
transform 1 0 26208 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_234
timestamp 1621261055
transform 1 0 23616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_242
timestamp 1621261055
transform 1 0 24384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_246
timestamp 1621261055
transform 1 0 24768 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_249
timestamp 1621261055
transform 1 0 25056 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_257
timestamp 1621261055
transform 1 0 25824 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input223
timestamp 1621261055
transform 1 0 26976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input226
timestamp 1621261055
transform 1 0 27744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input229
timestamp 1621261055
transform 1 0 28512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input231
timestamp 1621261055
transform 1 0 29280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_265
timestamp 1621261055
transform 1 0 26592 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_273
timestamp 1621261055
transform 1 0 27360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_281
timestamp 1621261055
transform 1 0 28128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_289
timestamp 1621261055
transform 1 0 28896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_297
timestamp 1621261055
transform 1 0 29664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_221
timestamp 1621261055
transform 1 0 30240 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input235
timestamp 1621261055
transform 1 0 30720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input237
timestamp 1621261055
transform 1 0 31488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input240
timestamp 1621261055
transform 1 0 32256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_301
timestamp 1621261055
transform 1 0 30048 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_304
timestamp 1621261055
transform 1 0 30336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_312
timestamp 1621261055
transform 1 0 31104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_320
timestamp 1621261055
transform 1 0 31872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_328
timestamp 1621261055
transform 1 0 32640 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input242
timestamp 1621261055
transform 1 0 33024 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_336
timestamp 1621261055
transform 1 0 33408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_344
timestamp 1621261055
transform 1 0 34176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input244
timestamp 1621261055
transform 1 0 33792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input246
timestamp 1621261055
transform 1 0 34560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_352
timestamp 1621261055
transform 1 0 34944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_356
timestamp 1621261055
transform 1 0 35328 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_222
timestamp 1621261055
transform 1 0 35520 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_359
timestamp 1621261055
transform 1 0 35616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input251
timestamp 1621261055
transform 1 0 36000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input253
timestamp 1621261055
transform 1 0 36768 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input255
timestamp 1621261055
transform 1 0 37536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input257
timestamp 1621261055
transform 1 0 38304 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input259
timestamp 1621261055
transform 1 0 39072 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_367
timestamp 1621261055
transform 1 0 36384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_375
timestamp 1621261055
transform 1 0 37152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_383
timestamp 1621261055
transform 1 0 37920 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_391
timestamp 1621261055
transform 1 0 38688 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_399
timestamp 1621261055
transform 1 0 39456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input263
timestamp 1621261055
transform 1 0 39840 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_407
timestamp 1621261055
transform 1 0 40224 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_414
timestamp 1621261055
transform 1 0 40896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_411
timestamp 1621261055
transform 1 0 40608 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_223
timestamp 1621261055
transform 1 0 40800 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input267
timestamp 1621261055
transform 1 0 41280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_422
timestamp 1621261055
transform 1 0 41664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_428
timestamp 1621261055
transform 1 0 42240 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_426
timestamp 1621261055
transform 1 0 42048 0 -1 5994
box -38 -49 230 715
use OAI21X1  OAI21X1
timestamp 1623610208
transform 1 0 42336 0 -1 5994
box 0 -48 1152 714
use sky130_fd_sc_ls__clkbuf_1  input273
timestamp 1621261055
transform 1 0 43872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input277
timestamp 1621261055
transform 1 0 44640 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_441
timestamp 1621261055
transform 1 0 43488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_449
timestamp 1621261055
transform 1 0 44256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_457
timestamp 1621261055
transform 1 0 45024 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_465
timestamp 1621261055
transform 1 0 45792 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_469
timestamp 1621261055
transform 1 0 46176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_467
timestamp 1621261055
transform 1 0 45984 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_224
timestamp 1621261055
transform 1 0 46080 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input282
timestamp 1621261055
transform 1 0 46560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_477
timestamp 1621261055
transform 1 0 46944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input285
timestamp 1621261055
transform 1 0 47328 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_485
timestamp 1621261055
transform 1 0 47712 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input287
timestamp 1621261055
transform 1 0 48096 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_493
timestamp 1621261055
transform 1 0 48480 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input289
timestamp 1621261055
transform 1 0 48864 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_501
timestamp 1621261055
transform 1 0 49248 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_509
timestamp 1621261055
transform 1 0 50016 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input290
timestamp 1621261055
transform 1 0 49632 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input292
timestamp 1621261055
transform 1 0 50400 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_517
timestamp 1621261055
transform 1 0 50784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_521
timestamp 1621261055
transform 1 0 51168 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_225
timestamp 1621261055
transform 1 0 51360 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_528
timestamp 1621261055
transform 1 0 51840 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_524
timestamp 1621261055
transform 1 0 51456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_530
timestamp 1621261055
transform 1 0 52032 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input174
timestamp 1621261055
transform 1 0 52128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_535
timestamp 1621261055
transform 1 0 52512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input175
timestamp 1621261055
transform 1 0 52896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_543
timestamp 1621261055
transform 1 0 53280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input176
timestamp 1621261055
transform 1 0 53664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_551
timestamp 1621261055
transform 1 0 54048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input179
timestamp 1621261055
transform 1 0 54432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_559
timestamp 1621261055
transform 1 0 54816 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_4
timestamp 1621261055
transform 1 0 55008 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _016_
timestamp 1621261055
transform 1 0 55200 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_4_566
timestamp 1621261055
transform 1 0 55488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input69
timestamp 1621261055
transform 1 0 55872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_574
timestamp 1621261055
transform 1 0 56256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_579
timestamp 1621261055
transform 1 0 56736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_226
timestamp 1621261055
transform 1 0 56640 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_4_585
timestamp 1621261055
transform 1 0 57312 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_583
timestamp 1621261055
transform 1 0 57120 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input63
timestamp 1621261055
transform 1 0 57408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_594
timestamp 1621261055
transform 1 0 58176 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_590
timestamp 1621261055
transform 1 0 57792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_9
timestamp 1621261055
transform -1 0 58848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_596
timestamp 1621261055
transform 1 0 58368 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input363
timestamp 1621261055
transform 1 0 1536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_10
timestamp 1621261055
transform 1 0 1152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_8
timestamp 1621261055
transform 1 0 1920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input364
timestamp 1621261055
transform 1 0 2304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_16
timestamp 1621261055
transform 1 0 2688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_20
timestamp 1621261055
transform 1 0 3072 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input357
timestamp 1621261055
transform 1 0 3168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_25
timestamp 1621261055
transform 1 0 3552 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_33
timestamp 1621261055
transform 1 0 4320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input359
timestamp 1621261055
transform 1 0 3936 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_227
timestamp 1621261055
transform 1 0 6432 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input361
timestamp 1621261055
transform 1 0 4704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output575
timestamp 1621261055
transform 1 0 5472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output577
timestamp 1621261055
transform 1 0 6912 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_41
timestamp 1621261055
transform 1 0 5088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_49
timestamp 1621261055
transform 1 0 5856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_53
timestamp 1621261055
transform 1 0 6240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_56
timestamp 1621261055
transform 1 0 6528 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_64
timestamp 1621261055
transform 1 0 7296 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output579
timestamp 1621261055
transform 1 0 7680 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_72
timestamp 1621261055
transform 1 0 8064 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_201
timestamp 1621261055
transform 1 0 8256 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_80
timestamp 1621261055
transform 1 0 8832 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output581
timestamp 1621261055
transform 1 0 8448 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_205
timestamp 1621261055
transform 1 0 9024 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output583
timestamp 1621261055
transform 1 0 9216 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_88
timestamp 1621261055
transform 1 0 9600 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_92
timestamp 1621261055
transform 1 0 9984 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input346
timestamp 1621261055
transform 1 0 10080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_97
timestamp 1621261055
transform 1 0 10464 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input348
timestamp 1621261055
transform 1 0 10848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_105
timestamp 1621261055
transform 1 0 11232 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_111
timestamp 1621261055
transform 1 0 11808 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_109
timestamp 1621261055
transform 1 0 11616 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_228
timestamp 1621261055
transform 1 0 11712 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input350
timestamp 1621261055
transform 1 0 12192 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_119
timestamp 1621261055
transform 1 0 12576 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input353
timestamp 1621261055
transform 1 0 12960 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_127
timestamp 1621261055
transform 1 0 13344 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output444
timestamp 1621261055
transform 1 0 13728 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_135
timestamp 1621261055
transform 1 0 14112 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output494
timestamp 1621261055
transform 1 0 14496 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_143
timestamp 1621261055
transform 1 0 14880 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_128
timestamp 1621261055
transform 1 0 15072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_151
timestamp 1621261055
transform 1 0 15648 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output505
timestamp 1621261055
transform 1 0 15264 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_155
timestamp 1621261055
transform 1 0 16032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input294
timestamp 1621261055
transform 1 0 16224 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_161
timestamp 1621261055
transform 1 0 16608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_229
timestamp 1621261055
transform 1 0 16992 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_166
timestamp 1621261055
transform 1 0 17088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_174
timestamp 1621261055
transform 1 0 17856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output455
timestamp 1621261055
transform 1 0 17472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output475
timestamp 1621261055
transform 1 0 18240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_182
timestamp 1621261055
transform 1 0 18624 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_104
timestamp 1621261055
transform 1 0 18816 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output477
timestamp 1621261055
transform 1 0 19008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_190
timestamp 1621261055
transform 1 0 19392 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_106
timestamp 1621261055
transform 1 0 19584 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_198
timestamp 1621261055
transform 1 0 20160 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output479
timestamp 1621261055
transform 1 0 19776 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_108
timestamp 1621261055
transform 1 0 20352 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output480
timestamp 1621261055
transform 1 0 20544 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_206
timestamp 1621261055
transform 1 0 20928 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_112
timestamp 1621261055
transform 1 0 21120 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output482
timestamp 1621261055
transform 1 0 21312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_214
timestamp 1621261055
transform 1 0 21696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_221
timestamp 1621261055
transform 1 0 22368 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_218
timestamp 1621261055
transform 1 0 22080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_230
timestamp 1621261055
transform 1 0 22272 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_116
timestamp 1621261055
transform 1 0 22560 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output487
timestamp 1621261055
transform 1 0 22752 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_229
timestamp 1621261055
transform 1 0 23136 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input222
timestamp 1621261055
transform 1 0 25632 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output489
timestamp 1621261055
transform 1 0 23520 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output491
timestamp 1621261055
transform 1 0 24288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_120
timestamp 1621261055
transform 1 0 24096 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_237
timestamp 1621261055
transform 1 0 23904 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_245
timestamp 1621261055
transform 1 0 24672 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_253
timestamp 1621261055
transform 1 0 25440 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_259
timestamp 1621261055
transform 1 0 26016 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input225
timestamp 1621261055
transform 1 0 26784 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_271
timestamp 1621261055
transform 1 0 27168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_276
timestamp 1621261055
transform 1 0 27648 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_124
timestamp 1621261055
transform -1 0 28032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_231
timestamp 1621261055
transform 1 0 27552 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output501
timestamp 1621261055
transform -1 0 28416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_284
timestamp 1621261055
transform 1 0 28416 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_126
timestamp 1621261055
transform 1 0 28608 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output504
timestamp 1621261055
transform 1 0 28800 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_292
timestamp 1621261055
transform 1 0 29184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_296
timestamp 1621261055
transform 1 0 29568 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input234
timestamp 1621261055
transform 1 0 29664 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_232
timestamp 1621261055
transform 1 0 32832 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input238
timestamp 1621261055
transform 1 0 31200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output509
timestamp 1621261055
transform 1 0 30432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output513
timestamp 1621261055
transform 1 0 31968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_301
timestamp 1621261055
transform 1 0 30048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_309
timestamp 1621261055
transform 1 0 30816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_317
timestamp 1621261055
transform 1 0 31584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_325
timestamp 1621261055
transform 1 0 32352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_329
timestamp 1621261055
transform 1 0 32736 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output518
timestamp 1621261055
transform 1 0 33312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output520
timestamp 1621261055
transform 1 0 34080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output522
timestamp 1621261055
transform 1 0 34848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_140
timestamp 1621261055
transform 1 0 33120 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_331
timestamp 1621261055
transform 1 0 32928 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_339
timestamp 1621261055
transform 1 0 33696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_347
timestamp 1621261055
transform 1 0 34464 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_355
timestamp 1621261055
transform 1 0 35232 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_363
timestamp 1621261055
transform 1 0 36000 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_365
timestamp 1621261055
transform 1 0 36192 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input254
timestamp 1621261055
transform 1 0 36288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_370
timestamp 1621261055
transform 1 0 36672 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_143
timestamp 1621261055
transform -1 0 37056 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output529
timestamp 1621261055
transform -1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_382
timestamp 1621261055
transform 1 0 37824 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_378
timestamp 1621261055
transform 1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_386
timestamp 1621261055
transform 1 0 38208 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_384
timestamp 1621261055
transform 1 0 38016 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_233
timestamp 1621261055
transform 1 0 38112 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_390
timestamp 1621261055
transform 1 0 38592 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_392
timestamp 1621261055
transform 1 0 38784 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input262
timestamp 1621261055
transform 1 0 38880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input266
timestamp 1621261055
transform 1 0 40320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input269
timestamp 1621261055
transform 1 0 41472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input270
timestamp 1621261055
transform 1 0 42240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_397
timestamp 1621261055
transform 1 0 39264 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_405
timestamp 1621261055
transform 1 0 40032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_407
timestamp 1621261055
transform 1 0 40224 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_5_412
timestamp 1621261055
transform 1 0 40704 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_5_424
timestamp 1621261055
transform 1 0 41856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_234
timestamp 1621261055
transform 1 0 43392 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input275
timestamp 1621261055
transform 1 0 43872 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input279
timestamp 1621261055
transform 1 0 44736 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input281
timestamp 1621261055
transform 1 0 45504 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_432
timestamp 1621261055
transform 1 0 42624 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_5_441
timestamp 1621261055
transform 1 0 43488 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_449
timestamp 1621261055
transform 1 0 44256 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_453
timestamp 1621261055
transform 1 0 44640 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_458
timestamp 1621261055
transform 1 0 45120 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_235
timestamp 1621261055
transform 1 0 48672 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input286
timestamp 1621261055
transform 1 0 46944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input288
timestamp 1621261055
transform 1 0 47712 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_466
timestamp 1621261055
transform 1 0 45888 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_474
timestamp 1621261055
transform 1 0 46656 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_476
timestamp 1621261055
transform 1 0 46848 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_481
timestamp 1621261055
transform 1 0 47328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_489
timestamp 1621261055
transform 1 0 48096 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_493
timestamp 1621261055
transform 1 0 48480 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_496
timestamp 1621261055
transform 1 0 48768 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_504
timestamp 1621261055
transform 1 0 49536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input291
timestamp 1621261055
transform 1 0 49152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input293
timestamp 1621261055
transform 1 0 49920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_512
timestamp 1621261055
transform 1 0 50304 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_74
timestamp 1621261055
transform -1 0 50688 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output445
timestamp 1621261055
transform -1 0 51072 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_520
timestamp 1621261055
transform 1 0 51072 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_528
timestamp 1621261055
transform 1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output447
timestamp 1621261055
transform 1 0 51456 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_236
timestamp 1621261055
transform 1 0 53952 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input180
timestamp 1621261055
transform 1 0 54432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input192
timestamp 1621261055
transform 1 0 53184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output448
timestamp 1621261055
transform 1 0 52224 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_536
timestamp 1621261055
transform 1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_540
timestamp 1621261055
transform 1 0 52992 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_546
timestamp 1621261055
transform 1 0 53568 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_551
timestamp 1621261055
transform 1 0 54048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_559
timestamp 1621261055
transform 1 0 54816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input65
timestamp 1621261055
transform 1 0 57696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input67
timestamp 1621261055
transform 1 0 56928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input181
timestamp 1621261055
transform 1 0 55200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input183
timestamp 1621261055
transform 1 0 55968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_567
timestamp 1621261055
transform 1 0 55584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_575
timestamp 1621261055
transform 1 0 56352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_579
timestamp 1621261055
transform 1 0 56736 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_585
timestamp 1621261055
transform 1 0 57312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_593
timestamp 1621261055
transform 1 0 58080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_11
timestamp 1621261055
transform -1 0 58848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_8
timestamp 1621261055
transform 1 0 1920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input366
timestamp 1621261055
transform 1 0 1536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_12
timestamp 1621261055
transform 1 0 1152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_12
timestamp 1621261055
transform 1 0 2304 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input365
timestamp 1621261055
transform 1 0 2496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_26
timestamp 1621261055
transform 1 0 3648 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_18
timestamp 1621261055
transform 1 0 2880 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_29
timestamp 1621261055
transform 1 0 3936 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_223
timestamp 1621261055
transform 1 0 4128 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output598
timestamp 1621261055
transform 1 0 4320 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_237
timestamp 1621261055
transform 1 0 3840 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_37
timestamp 1621261055
transform 1 0 4704 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output601
timestamp 1621261055
transform 1 0 5088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_45
timestamp 1621261055
transform 1 0 5472 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_195
timestamp 1621261055
transform 1 0 5664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output576
timestamp 1621261055
transform 1 0 5856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_53
timestamp 1621261055
transform 1 0 6240 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_197
timestamp 1621261055
transform 1 0 6432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output578
timestamp 1621261055
transform 1 0 6624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_61
timestamp 1621261055
transform 1 0 7008 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_199
timestamp 1621261055
transform 1 0 7200 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output580
timestamp 1621261055
transform 1 0 7392 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_69
timestamp 1621261055
transform 1 0 7776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_203
timestamp 1621261055
transform 1 0 7968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output582
timestamp 1621261055
transform 1 0 8160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_77
timestamp 1621261055
transform 1 0 8544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_84
timestamp 1621261055
transform 1 0 9216 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_81
timestamp 1621261055
transform 1 0 8928 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_238
timestamp 1621261055
transform 1 0 9120 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output585
timestamp 1621261055
transform 1 0 9600 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_92
timestamp 1621261055
transform 1 0 9984 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_209
timestamp 1621261055
transform 1 0 10176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output587
timestamp 1621261055
transform 1 0 10368 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_104
timestamp 1621261055
transform 1 0 11136 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_100
timestamp 1621261055
transform 1 0 10752 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input349
timestamp 1621261055
transform 1 0 11232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_109
timestamp 1621261055
transform 1 0 11616 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_6_124
timestamp 1621261055
transform 1 0 13056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_119
timestamp 1621261055
transform 1 0 12576 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_117
timestamp 1621261055
transform 1 0 12384 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input354
timestamp 1621261055
transform 1 0 12672 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_132
timestamp 1621261055
transform 1 0 13824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output483
timestamp 1621261055
transform 1 0 13440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_239
timestamp 1621261055
transform 1 0 14400 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output516
timestamp 1621261055
transform 1 0 14880 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output527
timestamp 1621261055
transform 1 0 15648 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_136
timestamp 1621261055
transform 1 0 14208 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_139
timestamp 1621261055
transform 1 0 14496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_147
timestamp 1621261055
transform 1 0 15264 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_155
timestamp 1621261055
transform 1 0 16032 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_163
timestamp 1621261055
transform 1 0 16800 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_165
timestamp 1621261055
transform 1 0 16992 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output466
timestamp 1621261055
transform 1 0 17088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_170
timestamp 1621261055
transform 1 0 17472 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_102
timestamp 1621261055
transform 1 0 17664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output476
timestamp 1621261055
transform 1 0 17856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_178
timestamp 1621261055
transform 1 0 18240 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output478
timestamp 1621261055
transform 1 0 18624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_186
timestamp 1621261055
transform 1 0 19008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_192
timestamp 1621261055
transform 1 0 19584 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_190
timestamp 1621261055
transform 1 0 19392 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_240
timestamp 1621261055
transform 1 0 19680 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_194
timestamp 1621261055
transform 1 0 19776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_110
timestamp 1621261055
transform 1 0 19968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output481
timestamp 1621261055
transform 1 0 20160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output484
timestamp 1621261055
transform 1 0 20928 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output486
timestamp 1621261055
transform 1 0 21696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output488
timestamp 1621261055
transform -1 0 22848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output490
timestamp 1621261055
transform 1 0 23232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_118
timestamp 1621261055
transform -1 0 22464 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_202
timestamp 1621261055
transform 1 0 20544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_210
timestamp 1621261055
transform 1 0 21312 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_218
timestamp 1621261055
transform 1 0 22080 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_226
timestamp 1621261055
transform 1 0 22848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_241
timestamp 1621261055
transform 1 0 24960 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output492
timestamp 1621261055
transform 1 0 24000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output496
timestamp 1621261055
transform 1 0 25440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output498
timestamp 1621261055
transform 1 0 26208 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_234
timestamp 1621261055
transform 1 0 23616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_242
timestamp 1621261055
transform 1 0 24384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_246
timestamp 1621261055
transform 1 0 24768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_249
timestamp 1621261055
transform 1 0 25056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_257
timestamp 1621261055
transform 1 0 25824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_265
timestamp 1621261055
transform 1 0 26592 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_273
timestamp 1621261055
transform 1 0 27360 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output500
timestamp 1621261055
transform 1 0 26976 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output503
timestamp 1621261055
transform 1 0 27744 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_281
timestamp 1621261055
transform 1 0 28128 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_130
timestamp 1621261055
transform -1 0 28512 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output506
timestamp 1621261055
transform -1 0 28896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_289
timestamp 1621261055
transform 1 0 28896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_297
timestamp 1621261055
transform 1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output508
timestamp 1621261055
transform 1 0 29280 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_242
timestamp 1621261055
transform 1 0 30240 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output512
timestamp 1621261055
transform 1 0 30720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output514
timestamp 1621261055
transform 1 0 31488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output517
timestamp 1621261055
transform 1 0 32256 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_301
timestamp 1621261055
transform 1 0 30048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_304
timestamp 1621261055
transform 1 0 30336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_312
timestamp 1621261055
transform 1 0 31104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_320
timestamp 1621261055
transform 1 0 31872 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_328
timestamp 1621261055
transform 1 0 32640 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output519
timestamp 1621261055
transform 1 0 33024 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_336
timestamp 1621261055
transform 1 0 33408 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_344
timestamp 1621261055
transform 1 0 34176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output521
timestamp 1621261055
transform 1 0 33792 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output524
timestamp 1621261055
transform 1 0 34560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_352
timestamp 1621261055
transform 1 0 34944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_356
timestamp 1621261055
transform 1 0 35328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_243
timestamp 1621261055
transform 1 0 35520 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_359
timestamp 1621261055
transform 1 0 35616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output528
timestamp 1621261055
transform 1 0 36000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_367
timestamp 1621261055
transform 1 0 36384 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_147
timestamp 1621261055
transform -1 0 36768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output531
timestamp 1621261055
transform -1 0 37152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_151
timestamp 1621261055
transform -1 0 37536 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_148
timestamp 1621261055
transform -1 0 37344 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output533
timestamp 1621261055
transform -1 0 37920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_383
timestamp 1621261055
transform 1 0 37920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output534
timestamp 1621261055
transform 1 0 38304 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_391
timestamp 1621261055
transform 1 0 38688 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_153
timestamp 1621261055
transform 1 0 38880 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output535
timestamp 1621261055
transform 1 0 39072 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_244
timestamp 1621261055
transform 1 0 40800 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output537
timestamp 1621261055
transform 1 0 39840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output542
timestamp 1621261055
transform 1 0 41280 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output544
timestamp 1621261055
transform 1 0 42048 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_399
timestamp 1621261055
transform 1 0 39456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_407
timestamp 1621261055
transform 1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_411
timestamp 1621261055
transform 1 0 40608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_414
timestamp 1621261055
transform 1 0 40896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_422
timestamp 1621261055
transform 1 0 41664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_430
timestamp 1621261055
transform 1 0 42432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_163
timestamp 1621261055
transform -1 0 42816 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_438
timestamp 1621261055
transform 1 0 43200 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output546
timestamp 1621261055
transform -1 0 43200 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output548
timestamp 1621261055
transform 1 0 43584 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_446
timestamp 1621261055
transform 1 0 43968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_171
timestamp 1621261055
transform 1 0 44160 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output551
timestamp 1621261055
transform 1 0 44352 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_454
timestamp 1621261055
transform 1 0 44736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_462
timestamp 1621261055
transform 1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output553
timestamp 1621261055
transform 1 0 45120 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_466
timestamp 1621261055
transform 1 0 45888 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_469
timestamp 1621261055
transform 1 0 46176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_245
timestamp 1621261055
transform 1 0 46080 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output557
timestamp 1621261055
transform 1 0 46560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_477
timestamp 1621261055
transform 1 0 46944 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_179
timestamp 1621261055
transform -1 0 47328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output559
timestamp 1621261055
transform -1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_485
timestamp 1621261055
transform 1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output562
timestamp 1621261055
transform 1 0 48096 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_493
timestamp 1621261055
transform 1 0 48480 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_246
timestamp 1621261055
transform 1 0 51360 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output446
timestamp 1621261055
transform 1 0 50112 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output449
timestamp 1621261055
transform 1 0 51840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output564
timestamp 1621261055
transform 1 0 48864 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_501
timestamp 1621261055
transform 1 0 49248 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_6_509
timestamp 1621261055
transform 1 0 50016 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_6_514
timestamp 1621261055
transform 1 0 50496 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_6_522
timestamp 1621261055
transform 1 0 51264 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_524
timestamp 1621261055
transform 1 0 51456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input182
timestamp 1621261055
transform 1 0 54720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input196
timestamp 1621261055
transform 1 0 53952 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output451
timestamp 1621261055
transform -1 0 52992 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_76
timestamp 1621261055
transform -1 0 52608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_532
timestamp 1621261055
transform 1 0 52224 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_540
timestamp 1621261055
transform 1 0 52992 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_548
timestamp 1621261055
transform 1 0 53760 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_554
timestamp 1621261055
transform 1 0 54336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_247
timestamp 1621261055
transform 1 0 56640 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input66
timestamp 1621261055
transform 1 0 57696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input184
timestamp 1621261055
transform 1 0 55488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_562
timestamp 1621261055
transform 1 0 55104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_570
timestamp 1621261055
transform 1 0 55872 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_6_579
timestamp 1621261055
transform 1 0 56736 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_587
timestamp 1621261055
transform 1 0 57504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_593
timestamp 1621261055
transform 1 0 58080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_13
timestamp 1621261055
transform -1 0 58848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output572
timestamp 1621261055
transform 1 0 1536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input367
timestamp 1621261055
transform 1 0 1536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_16
timestamp 1621261055
transform 1 0 1152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_14
timestamp 1621261055
transform 1 0 1152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_8
timestamp 1621261055
transform 1 0 1920 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_191
timestamp 1621261055
transform 1 0 1920 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_207
timestamp 1621261055
transform 1 0 2112 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_193
timestamp 1621261055
transform 1 0 2112 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output584
timestamp 1621261055
transform 1 0 2304 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output573
timestamp 1621261055
transform 1 0 2304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_16
timestamp 1621261055
transform 1 0 2688 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_16
timestamp 1621261055
transform 1 0 2688 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_225
timestamp 1621261055
transform 1 0 2880 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_219
timestamp 1621261055
transform 1 0 2880 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_24
timestamp 1621261055
transform 1 0 3456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_24
timestamp 1621261055
transform 1 0 3456 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output599
timestamp 1621261055
transform 1 0 3072 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output595
timestamp 1621261055
transform 1 0 3072 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output600
timestamp 1621261055
transform 1 0 3840 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_258
timestamp 1621261055
transform 1 0 3840 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_29
timestamp 1621261055
transform 1 0 3936 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_32
timestamp 1621261055
transform 1 0 4224 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_229
timestamp 1621261055
transform 1 0 4128 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output603
timestamp 1621261055
transform 1 0 4320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_37
timestamp 1621261055
transform 1 0 4704 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_40
timestamp 1621261055
transform 1 0 4992 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_227
timestamp 1621261055
transform 1 0 4416 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output602
timestamp 1621261055
transform 1 0 4608 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_45
timestamp 1621261055
transform 1 0 5472 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_48
timestamp 1621261055
transform 1 0 5760 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output604
timestamp 1621261055
transform 1 0 5376 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_53
timestamp 1621261055
transform 1 0 6240 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_56
timestamp 1621261055
transform 1 0 6528 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_54
timestamp 1621261055
transform 1 0 6336 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_52
timestamp 1621261055
transform 1 0 6144 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_248
timestamp 1621261055
transform 1 0 6432 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_63
timestamp 1621261055
transform 1 0 7200 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_61
timestamp 1621261055
transform 1 0 7008 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_64
timestamp 1621261055
transform 1 0 7296 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _106_
timestamp 1621261055
transform 1 0 7296 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_67
timestamp 1621261055
transform 1 0 7584 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_72
timestamp 1621261055
transform 1 0 8064 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_75
timestamp 1621261055
transform 1 0 8352 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_82
timestamp 1621261055
transform 1 0 9024 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_80
timestamp 1621261055
transform 1 0 8832 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output586
timestamp 1621261055
transform 1 0 9120 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_259
timestamp 1621261055
transform 1 0 9120 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_92
timestamp 1621261055
transform 1 0 9984 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_84
timestamp 1621261055
transform 1 0 9216 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_87
timestamp 1621261055
transform 1 0 9504 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output588
timestamp 1621261055
transform 1 0 9888 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_96
timestamp 1621261055
transform 1 0 10368 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_95
timestamp 1621261055
transform 1 0 10272 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_211
timestamp 1621261055
transform 1 0 10464 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output590
timestamp 1621261055
transform 1 0 10560 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output589
timestamp 1621261055
transform 1 0 10656 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_102
timestamp 1621261055
transform 1 0 10944 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_103
timestamp 1621261055
transform 1 0 11040 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_107
timestamp 1621261055
transform 1 0 11424 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_213
timestamp 1621261055
transform 1 0 11136 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output591
timestamp 1621261055
transform 1 0 11328 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_110
timestamp 1621261055
transform 1 0 11712 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_111
timestamp 1621261055
transform 1 0 11808 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_7_109
timestamp 1621261055
transform 1 0 11616 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_215
timestamp 1621261055
transform 1 0 12000 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_249
timestamp 1621261055
transform 1 0 11712 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_118
timestamp 1621261055
transform 1 0 12480 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output593
timestamp 1621261055
transform 1 0 12096 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output592
timestamp 1621261055
transform 1 0 12192 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_119
timestamp 1621261055
transform 1 0 12576 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_217
timestamp 1621261055
transform -1 0 12960 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output596
timestamp 1621261055
transform 1 0 12864 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output594
timestamp 1621261055
transform -1 0 13344 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_126
timestamp 1621261055
transform 1 0 13248 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_127
timestamp 1621261055
transform 1 0 13344 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_221
timestamp 1621261055
transform 1 0 13536 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output597
timestamp 1621261055
transform 1 0 13728 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _063_
timestamp 1621261055
transform 1 0 13632 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_139
timestamp 1621261055
transform 1 0 14496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_137
timestamp 1621261055
transform 1 0 14304 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_133
timestamp 1621261055
transform 1 0 13920 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_135
timestamp 1621261055
transform 1 0 14112 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_260
timestamp 1621261055
transform 1 0 14400 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_147
timestamp 1621261055
transform 1 0 15264 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_143
timestamp 1621261055
transform 1 0 14880 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_155
timestamp 1621261055
transform -1 0 15264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output538
timestamp 1621261055
transform -1 0 15648 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_151
timestamp 1621261055
transform 1 0 15648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_167
timestamp 1621261055
transform 1 0 15840 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output560
timestamp 1621261055
transform 1 0 16032 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output549
timestamp 1621261055
transform 1 0 16032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_159
timestamp 1621261055
transform 1 0 16416 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_163
timestamp 1621261055
transform 1 0 16800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_159
timestamp 1621261055
transform 1 0 16416 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_189
timestamp 1621261055
transform 1 0 16608 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output571
timestamp 1621261055
transform 1 0 16800 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_250
timestamp 1621261055
transform 1 0 16992 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_167
timestamp 1621261055
transform 1 0 17184 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_170
timestamp 1621261055
transform 1 0 17472 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_166
timestamp 1621261055
transform 1 0 17088 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_18
timestamp 1621261055
transform 1 0 17568 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _032_
timestamp 1621261055
transform 1 0 17760 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_175
timestamp 1621261055
transform 1 0 17952 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_176
timestamp 1621261055
transform 1 0 18048 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _132_
timestamp 1621261055
transform 1 0 18432 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_191
timestamp 1621261055
transform 1 0 19488 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_183
timestamp 1621261055
transform 1 0 18720 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_191
timestamp 1621261055
transform 1 0 19488 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_183
timestamp 1621261055
transform 1 0 18720 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_194
timestamp 1621261055
transform 1 0 19776 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_261
timestamp 1621261055
transform 1 0 19680 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_202
timestamp 1621261055
transform 1 0 20544 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_201
timestamp 1621261055
transform 1 0 20448 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_199
timestamp 1621261055
transform 1 0 20256 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_114
timestamp 1621261055
transform 1 0 20544 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output485
timestamp 1621261055
transform 1 0 20736 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_210
timestamp 1621261055
transform 1 0 21312 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_215
timestamp 1621261055
transform 1 0 21792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_208
timestamp 1621261055
transform 1 0 21120 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _203_
timestamp 1621261055
transform 1 0 21504 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_218
timestamp 1621261055
transform 1 0 22080 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_221
timestamp 1621261055
transform 1 0 22368 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_219
timestamp 1621261055
transform 1 0 22176 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_251
timestamp 1621261055
transform 1 0 22272 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_226
timestamp 1621261055
transform 1 0 22848 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_229
timestamp 1621261055
transform 1 0 23136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_234
timestamp 1621261055
transform 1 0 23616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_239
timestamp 1621261055
transform 1 0 24096 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_233
timestamp 1621261055
transform 1 0 23520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output493
timestamp 1621261055
transform 1 0 23712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_246
timestamp 1621261055
transform 1 0 24768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_242
timestamp 1621261055
transform 1 0 24384 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_247
timestamp 1621261055
transform 1 0 24864 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_122
timestamp 1621261055
transform 1 0 24288 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output495
timestamp 1621261055
transform 1 0 24480 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_262
timestamp 1621261055
transform 1 0 24960 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_257
timestamp 1621261055
transform 1 0 25824 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_249
timestamp 1621261055
transform 1 0 25056 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_255
timestamp 1621261055
transform 1 0 25632 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output497
timestamp 1621261055
transform 1 0 25248 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_263
timestamp 1621261055
transform 1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output499
timestamp 1621261055
transform 1 0 26016 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_265
timestamp 1621261055
transform 1 0 26592 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_271
timestamp 1621261055
transform 1 0 27168 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output502
timestamp 1621261055
transform 1 0 26784 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_281
timestamp 1621261055
transform 1 0 28128 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_273
timestamp 1621261055
transform 1 0 27360 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_278
timestamp 1621261055
transform 1 0 27840 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_276
timestamp 1621261055
transform 1 0 27648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_132
timestamp 1621261055
transform 1 0 27936 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output507
timestamp 1621261055
transform 1 0 28128 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_252
timestamp 1621261055
transform 1 0 27552 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_289
timestamp 1621261055
transform 1 0 28896 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_289
timestamp 1621261055
transform 1 0 28896 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_285
timestamp 1621261055
transform 1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_134
timestamp 1621261055
transform 1 0 28992 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_297
timestamp 1621261055
transform 1 0 29664 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_296
timestamp 1621261055
transform 1 0 29568 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output510
timestamp 1621261055
transform 1 0 29184 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_304
timestamp 1621261055
transform 1 0 30336 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_301
timestamp 1621261055
transform 1 0 30048 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_304
timestamp 1621261055
transform 1 0 30336 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_136
timestamp 1621261055
transform 1 0 29760 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output511
timestamp 1621261055
transform 1 0 29952 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_263
timestamp 1621261055
transform 1 0 30240 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_312
timestamp 1621261055
transform 1 0 31104 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_308
timestamp 1621261055
transform 1 0 30720 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_138
timestamp 1621261055
transform -1 0 31008 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output515
timestamp 1621261055
transform -1 0 31392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_320
timestamp 1621261055
transform 1 0 31872 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_315
timestamp 1621261055
transform 1 0 31392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _216_
timestamp 1621261055
transform 1 0 32160 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_328
timestamp 1621261055
transform 1 0 32640 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_326
timestamp 1621261055
transform 1 0 32448 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_253
timestamp 1621261055
transform 1 0 32832 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_336
timestamp 1621261055
transform 1 0 33408 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_337
timestamp 1621261055
transform 1 0 33504 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_335
timestamp 1621261055
transform 1 0 33312 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_331
timestamp 1621261055
transform 1 0 32928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output523
timestamp 1621261055
transform 1 0 33600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_344
timestamp 1621261055
transform 1 0 34176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_342
timestamp 1621261055
transform 1 0 33984 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_142
timestamp 1621261055
transform 1 0 34176 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output525
timestamp 1621261055
transform 1 0 34368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_356
timestamp 1621261055
transform 1 0 35328 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_352
timestamp 1621261055
transform 1 0 34944 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_350
timestamp 1621261055
transform 1 0 34752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output526
timestamp 1621261055
transform 1 0 35136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_359
timestamp 1621261055
transform 1 0 35616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_358
timestamp 1621261055
transform 1 0 35520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_145
timestamp 1621261055
transform -1 0 35904 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output530
timestamp 1621261055
transform -1 0 36288 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_264
timestamp 1621261055
transform 1 0 35520 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_367
timestamp 1621261055
transform 1 0 36384 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_366
timestamp 1621261055
transform 1 0 36288 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_149
timestamp 1621261055
transform -1 0 36672 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output532
timestamp 1621261055
transform -1 0 37056 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_375
timestamp 1621261055
transform 1 0 37152 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_374
timestamp 1621261055
transform 1 0 37056 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_383
timestamp 1621261055
transform 1 0 37920 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_386
timestamp 1621261055
transform 1 0 38208 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_384
timestamp 1621261055
transform 1 0 38016 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_382
timestamp 1621261055
transform 1 0 37824 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_254
timestamp 1621261055
transform 1 0 38112 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_393
timestamp 1621261055
transform 1 0 38880 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_391
timestamp 1621261055
transform 1 0 38688 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_394
timestamp 1621261055
transform 1 0 38976 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_159
timestamp 1621261055
transform -1 0 39168 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_157
timestamp 1621261055
transform -1 0 39360 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output540
timestamp 1621261055
transform -1 0 39552 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output536
timestamp 1621261055
transform 1 0 38592 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_400
timestamp 1621261055
transform 1 0 39552 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_402
timestamp 1621261055
transform 1 0 39744 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_161
timestamp 1621261055
transform -1 0 40128 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output539
timestamp 1621261055
transform -1 0 39744 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _212_
timestamp 1621261055
transform 1 0 39936 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_411
timestamp 1621261055
transform 1 0 40608 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_407
timestamp 1621261055
transform 1 0 40224 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_410
timestamp 1621261055
transform 1 0 40512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output541
timestamp 1621261055
transform -1 0 40512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_265
timestamp 1621261055
transform 1 0 40800 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_422
timestamp 1621261055
transform 1 0 41664 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_414
timestamp 1621261055
transform 1 0 40896 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_418
timestamp 1621261055
transform 1 0 41280 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output545
timestamp 1621261055
transform 1 0 41664 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output543
timestamp 1621261055
transform 1 0 40896 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_426
timestamp 1621261055
transform 1 0 42048 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_426
timestamp 1621261055
transform 1 0 42048 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_169
timestamp 1621261055
transform -1 0 42432 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_165
timestamp 1621261055
transform 1 0 42240 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_434
timestamp 1621261055
transform 1 0 42816 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_434
timestamp 1621261055
transform 1 0 42816 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output550
timestamp 1621261055
transform -1 0 42816 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output547
timestamp 1621261055
transform 1 0 42432 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_445
timestamp 1621261055
transform 1 0 43872 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_441
timestamp 1621261055
transform 1 0 43488 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_441
timestamp 1621261055
transform 1 0 43488 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_438
timestamp 1621261055
transform 1 0 43200 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_173
timestamp 1621261055
transform 1 0 43680 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output552
timestamp 1621261055
transform 1 0 43872 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_255
timestamp 1621261055
transform 1 0 43392 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _179_
timestamp 1621261055
transform 1 0 43200 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_453
timestamp 1621261055
transform 1 0 44640 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_449
timestamp 1621261055
transform 1 0 44256 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_176
timestamp 1621261055
transform -1 0 44256 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_175
timestamp 1621261055
transform -1 0 44640 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output555
timestamp 1621261055
transform -1 0 44640 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output554
timestamp 1621261055
transform -1 0 45024 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_461
timestamp 1621261055
transform 1 0 45408 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_457
timestamp 1621261055
transform 1 0 45024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_177
timestamp 1621261055
transform -1 0 45408 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output556
timestamp 1621261055
transform -1 0 45792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_469
timestamp 1621261055
transform 1 0 46176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_467
timestamp 1621261055
transform 1 0 45984 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_465
timestamp 1621261055
transform 1 0 45792 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_465
timestamp 1621261055
transform 1 0 45792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output558
timestamp 1621261055
transform 1 0 46176 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_266
timestamp 1621261055
transform 1 0 46080 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_477
timestamp 1621261055
transform 1 0 46944 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_473
timestamp 1621261055
transform 1 0 46560 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_180
timestamp 1621261055
transform -1 0 46944 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output561
timestamp 1621261055
transform -1 0 47328 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_488
timestamp 1621261055
transform 1 0 48000 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_481
timestamp 1621261055
transform 1 0 47328 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_481
timestamp 1621261055
transform 1 0 47328 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_182
timestamp 1621261055
transform 1 0 47424 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output565
timestamp 1621261055
transform 1 0 47616 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output563
timestamp 1621261055
transform 1 0 47712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_493
timestamp 1621261055
transform 1 0 48480 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_489
timestamp 1621261055
transform 1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_183
timestamp 1621261055
transform -1 0 48384 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output566
timestamp 1621261055
transform -1 0 48768 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_256
timestamp 1621261055
transform 1 0 48672 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_496
timestamp 1621261055
transform 1 0 48768 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_496
timestamp 1621261055
transform 1 0 48768 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_185
timestamp 1621261055
transform -1 0 49152 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output568
timestamp 1621261055
transform 1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output567
timestamp 1621261055
transform -1 0 49536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_512
timestamp 1621261055
transform 1 0 50304 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_8_504
timestamp 1621261055
transform 1 0 49536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_512
timestamp 1621261055
transform 1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_504
timestamp 1621261055
transform 1 0 49536 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_187
timestamp 1621261055
transform -1 0 49920 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output570
timestamp 1621261055
transform 1 0 49920 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output569
timestamp 1621261055
transform -1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_520
timestamp 1621261055
transform 1 0 51072 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_516
timestamp 1621261055
transform 1 0 50688 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output473
timestamp 1621261055
transform 1 0 50880 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_528
timestamp 1621261055
transform 1 0 51840 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_524
timestamp 1621261055
transform 1 0 51456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_522
timestamp 1621261055
transform 1 0 51264 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_522
timestamp 1621261055
transform 1 0 51264 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output450
timestamp 1621261055
transform 1 0 51648 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_267
timestamp 1621261055
transform 1 0 51360 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_530
timestamp 1621261055
transform 1 0 52032 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_530
timestamp 1621261055
transform 1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_99
timestamp 1621261055
transform -1 0 52320 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output472
timestamp 1621261055
transform -1 0 52704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output452
timestamp 1621261055
transform 1 0 52416 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_545
timestamp 1621261055
transform 1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_537
timestamp 1621261055
transform 1 0 52704 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_538
timestamp 1621261055
transform 1 0 52800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_79
timestamp 1621261055
transform -1 0 53088 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_78
timestamp 1621261055
transform -1 0 53184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output454
timestamp 1621261055
transform -1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output453
timestamp 1621261055
transform -1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_553
timestamp 1621261055
transform 1 0 54240 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_551
timestamp 1621261055
transform 1 0 54048 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_546
timestamp 1621261055
transform 1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output456
timestamp 1621261055
transform 1 0 53856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_257
timestamp 1621261055
transform 1 0 53952 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_561
timestamp 1621261055
transform 1 0 55008 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_559
timestamp 1621261055
transform 1 0 54816 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input194
timestamp 1621261055
transform 1 0 55008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_566
timestamp 1621261055
transform 1 0 55488 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_565
timestamp 1621261055
transform 1 0 55392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input197
timestamp 1621261055
transform 1 0 55104 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input185
timestamp 1621261055
transform 1 0 55776 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_574
timestamp 1621261055
transform 1 0 56256 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_573
timestamp 1621261055
transform 1 0 56160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input193
timestamp 1621261055
transform 1 0 55872 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input186
timestamp 1621261055
transform 1 0 56544 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_268
timestamp 1621261055
transform 1 0 56640 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_587
timestamp 1621261055
transform 1 0 57504 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_8_579
timestamp 1621261055
transform 1 0 56736 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_581
timestamp 1621261055
transform 1 0 56928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input188
timestamp 1621261055
transform 1 0 57120 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input187
timestamp 1621261055
transform 1 0 57312 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_589
timestamp 1621261055
transform 1 0 57696 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_15
timestamp 1621261055
transform -1 0 58848 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_17
timestamp 1621261055
transform -1 0 58848 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_595
timestamp 1621261055
transform 1 0 58272 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _061_
timestamp 1621261055
transform 1 0 3264 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _114_
timestamp 1621261055
transform 1 0 1536 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_18
timestamp 1621261055
transform 1 0 1152 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_7
timestamp 1621261055
transform 1 0 1824 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_15
timestamp 1621261055
transform 1 0 2592 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_19
timestamp 1621261055
transform 1 0 2976 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_21
timestamp 1621261055
transform 1 0 3168 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_25
timestamp 1621261055
transform 1 0 3552 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_33
timestamp 1621261055
transform 1 0 4320 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_269
timestamp 1621261055
transform 1 0 6432 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_41
timestamp 1621261055
transform 1 0 5088 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_49
timestamp 1621261055
transform 1 0 5856 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_53
timestamp 1621261055
transform 1 0 6240 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_56
timestamp 1621261055
transform 1 0 6528 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_64
timestamp 1621261055
transform 1 0 7296 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_72
timestamp 1621261055
transform 1 0 8064 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_80
timestamp 1621261055
transform 1 0 8832 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_88
timestamp 1621261055
transform 1 0 9600 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_96
timestamp 1621261055
transform 1 0 10368 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _011_
timestamp 1621261055
transform -1 0 11328 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_270
timestamp 1621261055
transform 1 0 11712 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_21
timestamp 1621261055
transform -1 0 11040 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_100
timestamp 1621261055
transform 1 0 10752 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_106
timestamp 1621261055
transform 1 0 11328 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_111
timestamp 1621261055
transform 1 0 11808 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_119
timestamp 1621261055
transform 1 0 12576 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_127
timestamp 1621261055
transform 1 0 13344 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_271
timestamp 1621261055
transform 1 0 16992 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_135
timestamp 1621261055
transform 1 0 14112 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_143
timestamp 1621261055
transform 1 0 14880 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_151
timestamp 1621261055
transform 1 0 15648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_159
timestamp 1621261055
transform 1 0 16416 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_163
timestamp 1621261055
transform 1 0 16800 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_166
timestamp 1621261055
transform 1 0 17088 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_174
timestamp 1621261055
transform 1 0 17856 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_182
timestamp 1621261055
transform 1 0 18624 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_190
timestamp 1621261055
transform 1 0 19392 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_198
timestamp 1621261055
transform 1 0 20160 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_272
timestamp 1621261055
transform 1 0 22272 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_206
timestamp 1621261055
transform 1 0 20928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_214
timestamp 1621261055
transform 1 0 21696 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_218
timestamp 1621261055
transform 1 0 22080 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_221
timestamp 1621261055
transform 1 0 22368 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_229
timestamp 1621261055
transform 1 0 23136 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_237
timestamp 1621261055
transform 1 0 23904 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_245
timestamp 1621261055
transform 1 0 24672 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_253
timestamp 1621261055
transform 1 0 25440 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_261
timestamp 1621261055
transform 1 0 26208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_273
timestamp 1621261055
transform 1 0 27552 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_269
timestamp 1621261055
transform 1 0 26976 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_273
timestamp 1621261055
transform 1 0 27360 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_276
timestamp 1621261055
transform 1 0 27648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_284
timestamp 1621261055
transform 1 0 28416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_292
timestamp 1621261055
transform 1 0 29184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_274
timestamp 1621261055
transform 1 0 32832 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_300
timestamp 1621261055
transform 1 0 29952 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_308
timestamp 1621261055
transform 1 0 30720 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_316
timestamp 1621261055
transform 1 0 31488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_324
timestamp 1621261055
transform 1 0 32256 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_328
timestamp 1621261055
transform 1 0 32640 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_331
timestamp 1621261055
transform 1 0 32928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_339
timestamp 1621261055
transform 1 0 33696 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_347
timestamp 1621261055
transform 1 0 34464 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_355
timestamp 1621261055
transform 1 0 35232 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_363
timestamp 1621261055
transform 1 0 36000 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _210_
timestamp 1621261055
transform 1 0 38592 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_275
timestamp 1621261055
transform 1 0 38112 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_371
timestamp 1621261055
transform 1 0 36768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_379
timestamp 1621261055
transform 1 0 37536 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_383
timestamp 1621261055
transform 1 0 37920 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_9_386
timestamp 1621261055
transform 1 0 38208 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_393
timestamp 1621261055
transform 1 0 38880 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_401
timestamp 1621261055
transform 1 0 39648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_409
timestamp 1621261055
transform 1 0 40416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_417
timestamp 1621261055
transform 1 0 41184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_425
timestamp 1621261055
transform 1 0 41952 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_276
timestamp 1621261055
transform 1 0 43392 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_433
timestamp 1621261055
transform 1 0 42720 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_437
timestamp 1621261055
transform 1 0 43104 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_439
timestamp 1621261055
transform 1 0 43296 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_441
timestamp 1621261055
transform 1 0 43488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_449
timestamp 1621261055
transform 1 0 44256 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_457
timestamp 1621261055
transform 1 0 45024 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_277
timestamp 1621261055
transform 1 0 48672 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_465
timestamp 1621261055
transform 1 0 45792 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_473
timestamp 1621261055
transform 1 0 46560 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_481
timestamp 1621261055
transform 1 0 47328 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_489
timestamp 1621261055
transform 1 0 48096 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_493
timestamp 1621261055
transform 1 0 48480 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_496
timestamp 1621261055
transform 1 0 48768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_504
timestamp 1621261055
transform 1 0 49536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_512
timestamp 1621261055
transform 1 0 50304 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_520
timestamp 1621261055
transform 1 0 51072 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_528
timestamp 1621261055
transform 1 0 51840 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_532
timestamp 1621261055
transform 1 0 52224 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_534
timestamp 1621261055
transform 1 0 52416 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _136_
timestamp 1621261055
transform 1 0 52512 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_538
timestamp 1621261055
transform 1 0 52800 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_94
timestamp 1621261055
transform -1 0 53184 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output469
timestamp 1621261055
transform -1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_546
timestamp 1621261055
transform 1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_551
timestamp 1621261055
transform 1 0 54048 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_278
timestamp 1621261055
transform 1 0 53952 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_80
timestamp 1621261055
transform -1 0 54432 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output457
timestamp 1621261055
transform -1 0 54816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_559
timestamp 1621261055
transform 1 0 54816 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_81
timestamp 1621261055
transform -1 0 55200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input190
timestamp 1621261055
transform 1 0 57216 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input195
timestamp 1621261055
transform 1 0 56448 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output459
timestamp 1621261055
transform -1 0 55584 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_567
timestamp 1621261055
transform 1 0 55584 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_9_575
timestamp 1621261055
transform 1 0 56352 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_580
timestamp 1621261055
transform 1 0 56832 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_588
timestamp 1621261055
transform 1 0 57600 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_19
timestamp 1621261055
transform -1 0 58848 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_596
timestamp 1621261055
transform 1 0 58368 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_20
timestamp 1621261055
transform 1 0 1152 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_279
timestamp 1621261055
transform 1 0 3840 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_60
timestamp 1621261055
transform -1 0 4512 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_4
timestamp 1621261055
transform 1 0 1536 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_12
timestamp 1621261055
transform 1 0 2304 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_20
timestamp 1621261055
transform 1 0 3072 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_29
timestamp 1621261055
transform 1 0 3936 0 -1 9990
box -38 -49 422 715
use INVX8  INVX8
timestamp 1623610208
transform -1 0 5952 0 -1 9990
box 0 -48 1440 714
use sky130_fd_sc_ls__decap_8  FILLER_10_50
timestamp 1621261055
transform 1 0 5952 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_58
timestamp 1621261055
transform 1 0 6720 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_66
timestamp 1621261055
transform 1 0 7488 0 -1 9990
box -38 -49 806 715
use INVX2  INVX2
timestamp 1623610208
transform 1 0 9600 0 -1 9990
box 0 -48 576 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_280
timestamp 1621261055
transform 1 0 9120 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_74
timestamp 1621261055
transform 1 0 8256 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_10_82
timestamp 1621261055
transform 1 0 9024 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_84
timestamp 1621261055
transform 1 0 9216 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_94
timestamp 1621261055
transform 1 0 10176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_102
timestamp 1621261055
transform 1 0 10944 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_110
timestamp 1621261055
transform 1 0 11712 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_118
timestamp 1621261055
transform 1 0 12480 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_126
timestamp 1621261055
transform 1 0 13248 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_281
timestamp 1621261055
transform 1 0 14400 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_134
timestamp 1621261055
transform 1 0 14016 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_139
timestamp 1621261055
transform 1 0 14496 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_147
timestamp 1621261055
transform 1 0 15264 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_155
timestamp 1621261055
transform 1 0 16032 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_163
timestamp 1621261055
transform 1 0 16800 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_282
timestamp 1621261055
transform 1 0 19680 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_171
timestamp 1621261055
transform 1 0 17568 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_179
timestamp 1621261055
transform 1 0 18336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_187
timestamp 1621261055
transform 1 0 19104 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_191
timestamp 1621261055
transform 1 0 19488 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_194
timestamp 1621261055
transform 1 0 19776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_202
timestamp 1621261055
transform 1 0 20544 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_210
timestamp 1621261055
transform 1 0 21312 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_218
timestamp 1621261055
transform 1 0 22080 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_226
timestamp 1621261055
transform 1 0 22848 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _042_
timestamp 1621261055
transform -1 0 26688 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_283
timestamp 1621261055
transform 1 0 24960 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_34
timestamp 1621261055
transform -1 0 26400 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_234
timestamp 1621261055
transform 1 0 23616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_242
timestamp 1621261055
transform 1 0 24384 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_246
timestamp 1621261055
transform 1 0 24768 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_249
timestamp 1621261055
transform 1 0 25056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_257
timestamp 1621261055
transform 1 0 25824 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_266
timestamp 1621261055
transform 1 0 26688 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_274
timestamp 1621261055
transform 1 0 27456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_282
timestamp 1621261055
transform 1 0 28224 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_290
timestamp 1621261055
transform 1 0 28992 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_284
timestamp 1621261055
transform 1 0 30240 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_298
timestamp 1621261055
transform 1 0 29760 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_302
timestamp 1621261055
transform 1 0 30144 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_304
timestamp 1621261055
transform 1 0 30336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_312
timestamp 1621261055
transform 1 0 31104 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_320
timestamp 1621261055
transform 1 0 31872 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_328
timestamp 1621261055
transform 1 0 32640 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_285
timestamp 1621261055
transform 1 0 35520 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_336
timestamp 1621261055
transform 1 0 33408 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_344
timestamp 1621261055
transform 1 0 34176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_352
timestamp 1621261055
transform 1 0 34944 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_356
timestamp 1621261055
transform 1 0 35328 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_359
timestamp 1621261055
transform 1 0 35616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_367
timestamp 1621261055
transform 1 0 36384 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_375
timestamp 1621261055
transform 1 0 37152 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_383
timestamp 1621261055
transform 1 0 37920 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_391
timestamp 1621261055
transform 1 0 38688 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_286
timestamp 1621261055
transform 1 0 40800 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_399
timestamp 1621261055
transform 1 0 39456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_407
timestamp 1621261055
transform 1 0 40224 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_411
timestamp 1621261055
transform 1 0 40608 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_414
timestamp 1621261055
transform 1 0 40896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_422
timestamp 1621261055
transform 1 0 41664 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _113_
timestamp 1621261055
transform 1 0 45408 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_10_430
timestamp 1621261055
transform 1 0 42432 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_438
timestamp 1621261055
transform 1 0 43200 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_446
timestamp 1621261055
transform 1 0 43968 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_454
timestamp 1621261055
transform 1 0 44736 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_458
timestamp 1621261055
transform 1 0 45120 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_460
timestamp 1621261055
transform 1 0 45312 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _091_
timestamp 1621261055
transform 1 0 46560 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_287
timestamp 1621261055
transform 1 0 46080 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_464
timestamp 1621261055
transform 1 0 45696 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_469
timestamp 1621261055
transform 1 0 46176 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_476
timestamp 1621261055
transform 1 0 46848 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_484
timestamp 1621261055
transform 1 0 47616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_492
timestamp 1621261055
transform 1 0 48384 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_288
timestamp 1621261055
transform 1 0 51360 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_500
timestamp 1621261055
transform 1 0 49152 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_508
timestamp 1621261055
transform 1 0 49920 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_516
timestamp 1621261055
transform 1 0 50688 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_520
timestamp 1621261055
transform 1 0 51072 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_522
timestamp 1621261055
transform 1 0 51264 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_524
timestamp 1621261055
transform 1 0 51456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _040_
timestamp 1621261055
transform -1 0 53856 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output458
timestamp 1621261055
transform 1 0 54240 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output460
timestamp 1621261055
transform -1 0 55392 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_69
timestamp 1621261055
transform -1 0 53568 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_83
timestamp 1621261055
transform -1 0 55008 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_532
timestamp 1621261055
transform 1 0 52224 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_540
timestamp 1621261055
transform 1 0 52992 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_549
timestamp 1621261055
transform 1 0 53856 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_557
timestamp 1621261055
transform 1 0 54624 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_565
timestamp 1621261055
transform 1 0 55392 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_85
timestamp 1621261055
transform -1 0 55776 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output461
timestamp 1621261055
transform -1 0 56160 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_577
timestamp 1621261055
transform 1 0 56544 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_575
timestamp 1621261055
transform 1 0 56352 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_86
timestamp 1621261055
transform -1 0 56352 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_289
timestamp 1621261055
transform 1 0 56640 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_10_587
timestamp 1621261055
transform 1 0 57504 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_579
timestamp 1621261055
transform 1 0 56736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_592
timestamp 1621261055
transform 1 0 57984 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input191
timestamp 1621261055
transform 1 0 57600 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_21
timestamp 1621261055
transform -1 0 58848 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_596
timestamp 1621261055
transform 1 0 58368 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_22
timestamp 1621261055
transform 1 0 1152 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_4
timestamp 1621261055
transform 1 0 1536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_12
timestamp 1621261055
transform 1 0 2304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_20
timestamp 1621261055
transform 1 0 3072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_28
timestamp 1621261055
transform 1 0 3840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_290
timestamp 1621261055
transform 1 0 6432 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_36
timestamp 1621261055
transform 1 0 4608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_44
timestamp 1621261055
transform 1 0 5376 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_52
timestamp 1621261055
transform 1 0 6144 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_54
timestamp 1621261055
transform 1 0 6336 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_56
timestamp 1621261055
transform 1 0 6528 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_64
timestamp 1621261055
transform 1 0 7296 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_72
timestamp 1621261055
transform 1 0 8064 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_80
timestamp 1621261055
transform 1 0 8832 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_88
timestamp 1621261055
transform 1 0 9600 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_96
timestamp 1621261055
transform 1 0 10368 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _162_
timestamp 1621261055
transform 1 0 12384 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_291
timestamp 1621261055
transform 1 0 11712 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_104
timestamp 1621261055
transform 1 0 11136 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_108
timestamp 1621261055
transform 1 0 11520 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_111
timestamp 1621261055
transform 1 0 11808 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_115
timestamp 1621261055
transform 1 0 12192 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_120
timestamp 1621261055
transform 1 0 12672 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_128
timestamp 1621261055
transform 1 0 13440 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_292
timestamp 1621261055
transform 1 0 16992 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_136
timestamp 1621261055
transform 1 0 14208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_144
timestamp 1621261055
transform 1 0 14976 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_152
timestamp 1621261055
transform 1 0 15744 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_160
timestamp 1621261055
transform 1 0 16512 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_164
timestamp 1621261055
transform 1 0 16896 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_166
timestamp 1621261055
transform 1 0 17088 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_174
timestamp 1621261055
transform 1 0 17856 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_182
timestamp 1621261055
transform 1 0 18624 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_190
timestamp 1621261055
transform 1 0 19392 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_198
timestamp 1621261055
transform 1 0 20160 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_293
timestamp 1621261055
transform 1 0 22272 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_206
timestamp 1621261055
transform 1 0 20928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_214
timestamp 1621261055
transform 1 0 21696 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_218
timestamp 1621261055
transform 1 0 22080 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_221
timestamp 1621261055
transform 1 0 22368 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_229
timestamp 1621261055
transform 1 0 23136 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_237
timestamp 1621261055
transform 1 0 23904 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_245
timestamp 1621261055
transform 1 0 24672 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_253
timestamp 1621261055
transform 1 0 25440 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_261
timestamp 1621261055
transform 1 0 26208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_294
timestamp 1621261055
transform 1 0 27552 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_269
timestamp 1621261055
transform 1 0 26976 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_273
timestamp 1621261055
transform 1 0 27360 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_276
timestamp 1621261055
transform 1 0 27648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_284
timestamp 1621261055
transform 1 0 28416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_292
timestamp 1621261055
transform 1 0 29184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_295
timestamp 1621261055
transform 1 0 32832 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_300
timestamp 1621261055
transform 1 0 29952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_308
timestamp 1621261055
transform 1 0 30720 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_316
timestamp 1621261055
transform 1 0 31488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_324
timestamp 1621261055
transform 1 0 32256 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_328
timestamp 1621261055
transform 1 0 32640 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_331
timestamp 1621261055
transform 1 0 32928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_339
timestamp 1621261055
transform 1 0 33696 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_347
timestamp 1621261055
transform 1 0 34464 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_355
timestamp 1621261055
transform 1 0 35232 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_363
timestamp 1621261055
transform 1 0 36000 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _145_
timestamp 1621261055
transform 1 0 38592 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_296
timestamp 1621261055
transform 1 0 38112 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_371
timestamp 1621261055
transform 1 0 36768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_379
timestamp 1621261055
transform 1 0 37536 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_383
timestamp 1621261055
transform 1 0 37920 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_386
timestamp 1621261055
transform 1 0 38208 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_393
timestamp 1621261055
transform 1 0 38880 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_401
timestamp 1621261055
transform 1 0 39648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_409
timestamp 1621261055
transform 1 0 40416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_417
timestamp 1621261055
transform 1 0 41184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_425
timestamp 1621261055
transform 1 0 41952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_297
timestamp 1621261055
transform 1 0 43392 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_433
timestamp 1621261055
transform 1 0 42720 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_437
timestamp 1621261055
transform 1 0 43104 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_439
timestamp 1621261055
transform 1 0 43296 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_441
timestamp 1621261055
transform 1 0 43488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_449
timestamp 1621261055
transform 1 0 44256 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_457
timestamp 1621261055
transform 1 0 45024 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_298
timestamp 1621261055
transform 1 0 48672 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_465
timestamp 1621261055
transform 1 0 45792 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_473
timestamp 1621261055
transform 1 0 46560 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_481
timestamp 1621261055
transform 1 0 47328 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_489
timestamp 1621261055
transform 1 0 48096 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_493
timestamp 1621261055
transform 1 0 48480 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_496
timestamp 1621261055
transform 1 0 48768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_504
timestamp 1621261055
transform 1 0 49536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_512
timestamp 1621261055
transform 1 0 50304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_520
timestamp 1621261055
transform 1 0 51072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_528
timestamp 1621261055
transform 1 0 51840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_299
timestamp 1621261055
transform 1 0 53952 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output471
timestamp 1621261055
transform -1 0 55296 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_96
timestamp 1621261055
transform -1 0 54912 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_536
timestamp 1621261055
transform 1 0 52608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_544
timestamp 1621261055
transform 1 0 53376 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_548
timestamp 1621261055
transform 1 0 53760 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_551
timestamp 1621261055
transform 1 0 54048 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_555
timestamp 1621261055
transform 1 0 54432 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_557
timestamp 1621261055
transform 1 0 54624 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output462
timestamp 1621261055
transform 1 0 55680 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output463
timestamp 1621261055
transform -1 0 56832 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output464
timestamp 1621261055
transform 1 0 57216 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_88
timestamp 1621261055
transform -1 0 56448 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_97
timestamp 1621261055
transform -1 0 55488 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_566
timestamp 1621261055
transform 1 0 55488 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_572
timestamp 1621261055
transform 1 0 56064 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_580
timestamp 1621261055
transform 1 0 56832 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_588
timestamp 1621261055
transform 1 0 57600 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_23
timestamp 1621261055
transform -1 0 58848 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_596
timestamp 1621261055
transform 1 0 58368 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_24
timestamp 1621261055
transform 1 0 1152 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_300
timestamp 1621261055
transform 1 0 3840 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_4
timestamp 1621261055
transform 1 0 1536 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_12
timestamp 1621261055
transform 1 0 2304 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_20
timestamp 1621261055
transform 1 0 3072 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_29
timestamp 1621261055
transform 1 0 3936 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _065_
timestamp 1621261055
transform 1 0 6720 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_37
timestamp 1621261055
transform 1 0 4704 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_45
timestamp 1621261055
transform 1 0 5472 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_53
timestamp 1621261055
transform 1 0 6240 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_12_57
timestamp 1621261055
transform 1 0 6624 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_61
timestamp 1621261055
transform 1 0 7008 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_301
timestamp 1621261055
transform 1 0 9120 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_69
timestamp 1621261055
transform 1 0 7776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_77
timestamp 1621261055
transform 1 0 8544 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_81
timestamp 1621261055
transform 1 0 8928 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_84
timestamp 1621261055
transform 1 0 9216 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_92
timestamp 1621261055
transform 1 0 9984 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_100
timestamp 1621261055
transform 1 0 10752 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_108
timestamp 1621261055
transform 1 0 11520 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_116
timestamp 1621261055
transform 1 0 12288 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_124
timestamp 1621261055
transform 1 0 13056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_132
timestamp 1621261055
transform 1 0 13824 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _100_
timestamp 1621261055
transform 1 0 15456 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_302
timestamp 1621261055
transform 1 0 14400 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_136
timestamp 1621261055
transform 1 0 14208 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_139
timestamp 1621261055
transform 1 0 14496 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_147
timestamp 1621261055
transform 1 0 15264 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_152
timestamp 1621261055
transform 1 0 15744 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_160
timestamp 1621261055
transform 1 0 16512 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_303
timestamp 1621261055
transform 1 0 19680 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_168
timestamp 1621261055
transform 1 0 17280 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_176
timestamp 1621261055
transform 1 0 18048 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_184
timestamp 1621261055
transform 1 0 18816 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_12_192
timestamp 1621261055
transform 1 0 19584 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_194
timestamp 1621261055
transform 1 0 19776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_202
timestamp 1621261055
transform 1 0 20544 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_210
timestamp 1621261055
transform 1 0 21312 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_218
timestamp 1621261055
transform 1 0 22080 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_226
timestamp 1621261055
transform 1 0 22848 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_304
timestamp 1621261055
transform 1 0 24960 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_234
timestamp 1621261055
transform 1 0 23616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_242
timestamp 1621261055
transform 1 0 24384 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_246
timestamp 1621261055
transform 1 0 24768 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_249
timestamp 1621261055
transform 1 0 25056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_257
timestamp 1621261055
transform 1 0 25824 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_265
timestamp 1621261055
transform 1 0 26592 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_273
timestamp 1621261055
transform 1 0 27360 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_281
timestamp 1621261055
transform 1 0 28128 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_289
timestamp 1621261055
transform 1 0 28896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_297
timestamp 1621261055
transform 1 0 29664 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _008_
timestamp 1621261055
transform -1 0 31488 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_305
timestamp 1621261055
transform 1 0 30240 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_12
timestamp 1621261055
transform -1 0 31200 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_301
timestamp 1621261055
transform 1 0 30048 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_12_304
timestamp 1621261055
transform 1 0 30336 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_308
timestamp 1621261055
transform 1 0 30720 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_310
timestamp 1621261055
transform 1 0 30912 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_316
timestamp 1621261055
transform 1 0 31488 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_324
timestamp 1621261055
transform 1 0 32256 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_306
timestamp 1621261055
transform 1 0 35520 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_332
timestamp 1621261055
transform 1 0 33024 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_340
timestamp 1621261055
transform 1 0 33792 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_348
timestamp 1621261055
transform 1 0 34560 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_356
timestamp 1621261055
transform 1 0 35328 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_359
timestamp 1621261055
transform 1 0 35616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_367
timestamp 1621261055
transform 1 0 36384 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_375
timestamp 1621261055
transform 1 0 37152 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_383
timestamp 1621261055
transform 1 0 37920 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_391
timestamp 1621261055
transform 1 0 38688 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_307
timestamp 1621261055
transform 1 0 40800 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_399
timestamp 1621261055
transform 1 0 39456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_407
timestamp 1621261055
transform 1 0 40224 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_411
timestamp 1621261055
transform 1 0 40608 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_414
timestamp 1621261055
transform 1 0 40896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_422
timestamp 1621261055
transform 1 0 41664 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _127_
timestamp 1621261055
transform 1 0 42432 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_433
timestamp 1621261055
transform 1 0 42720 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_441
timestamp 1621261055
transform 1 0 43488 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_449
timestamp 1621261055
transform 1 0 44256 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_457
timestamp 1621261055
transform 1 0 45024 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_308
timestamp 1621261055
transform 1 0 46080 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_465
timestamp 1621261055
transform 1 0 45792 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_467
timestamp 1621261055
transform 1 0 45984 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_469
timestamp 1621261055
transform 1 0 46176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_477
timestamp 1621261055
transform 1 0 46944 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_485
timestamp 1621261055
transform 1 0 47712 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_493
timestamp 1621261055
transform 1 0 48480 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_309
timestamp 1621261055
transform 1 0 51360 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_501
timestamp 1621261055
transform 1 0 49248 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_509
timestamp 1621261055
transform 1 0 50016 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_517
timestamp 1621261055
transform 1 0 50784 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_521
timestamp 1621261055
transform 1 0 51168 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_524
timestamp 1621261055
transform 1 0 51456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _163_
timestamp 1621261055
transform 1 0 54144 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_532
timestamp 1621261055
transform 1 0 52224 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_540
timestamp 1621261055
transform 1 0 52992 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_548
timestamp 1621261055
transform 1 0 53760 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_555
timestamp 1621261055
transform 1 0 54432 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_310
timestamp 1621261055
transform 1 0 56640 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output465
timestamp 1621261055
transform 1 0 57120 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output470
timestamp 1621261055
transform 1 0 55872 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_12_563
timestamp 1621261055
transform 1 0 55200 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_567
timestamp 1621261055
transform 1 0 55584 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_569
timestamp 1621261055
transform 1 0 55776 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_574
timestamp 1621261055
transform 1 0 56256 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_12_579
timestamp 1621261055
transform 1 0 56736 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_587
timestamp 1621261055
transform 1 0 57504 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_25
timestamp 1621261055
transform -1 0 58848 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_595
timestamp 1621261055
transform 1 0 58272 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_26
timestamp 1621261055
transform 1 0 1152 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_4
timestamp 1621261055
transform 1 0 1536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_12
timestamp 1621261055
transform 1 0 2304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_20
timestamp 1621261055
transform 1 0 3072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_28
timestamp 1621261055
transform 1 0 3840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_311
timestamp 1621261055
transform 1 0 6432 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_36
timestamp 1621261055
transform 1 0 4608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_44
timestamp 1621261055
transform 1 0 5376 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_52
timestamp 1621261055
transform 1 0 6144 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_54
timestamp 1621261055
transform 1 0 6336 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_56
timestamp 1621261055
transform 1 0 6528 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_64
timestamp 1621261055
transform 1 0 7296 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_72
timestamp 1621261055
transform 1 0 8064 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_80
timestamp 1621261055
transform 1 0 8832 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_88
timestamp 1621261055
transform 1 0 9600 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_96
timestamp 1621261055
transform 1 0 10368 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_312
timestamp 1621261055
transform 1 0 11712 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_104
timestamp 1621261055
transform 1 0 11136 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_108
timestamp 1621261055
transform 1 0 11520 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_111
timestamp 1621261055
transform 1 0 11808 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_119
timestamp 1621261055
transform 1 0 12576 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_127
timestamp 1621261055
transform 1 0 13344 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _164_
timestamp 1621261055
transform 1 0 14400 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_313
timestamp 1621261055
transform 1 0 16992 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_135
timestamp 1621261055
transform 1 0 14112 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_137
timestamp 1621261055
transform 1 0 14304 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_141
timestamp 1621261055
transform 1 0 14688 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_149
timestamp 1621261055
transform 1 0 15456 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_157
timestamp 1621261055
transform 1 0 16224 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_166
timestamp 1621261055
transform 1 0 17088 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_174
timestamp 1621261055
transform 1 0 17856 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_182
timestamp 1621261055
transform 1 0 18624 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_190
timestamp 1621261055
transform 1 0 19392 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_198
timestamp 1621261055
transform 1 0 20160 0 1 11322
box -38 -49 806 715
use INVX4  INVX4
timestamp 1623610208
transform -1 0 23616 0 1 11322
box 0 -48 864 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_314
timestamp 1621261055
transform 1 0 22272 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_55
timestamp 1621261055
transform -1 0 22752 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_206
timestamp 1621261055
transform 1 0 20928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_214
timestamp 1621261055
transform 1 0 21696 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_218
timestamp 1621261055
transform 1 0 22080 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_221
timestamp 1621261055
transform 1 0 22368 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_234
timestamp 1621261055
transform 1 0 23616 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_242
timestamp 1621261055
transform 1 0 24384 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_250
timestamp 1621261055
transform 1 0 25152 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_258
timestamp 1621261055
transform 1 0 25920 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _192_
timestamp 1621261055
transform 1 0 29088 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_315
timestamp 1621261055
transform 1 0 27552 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_266
timestamp 1621261055
transform 1 0 26688 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_13_274
timestamp 1621261055
transform 1 0 27456 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_276
timestamp 1621261055
transform 1 0 27648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_284
timestamp 1621261055
transform 1 0 28416 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_288
timestamp 1621261055
transform 1 0 28800 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_290
timestamp 1621261055
transform 1 0 28992 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_294
timestamp 1621261055
transform 1 0 29376 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_316
timestamp 1621261055
transform 1 0 32832 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_302
timestamp 1621261055
transform 1 0 30144 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_310
timestamp 1621261055
transform 1 0 30912 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_318
timestamp 1621261055
transform 1 0 31680 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_326
timestamp 1621261055
transform 1 0 32448 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_331
timestamp 1621261055
transform 1 0 32928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_339
timestamp 1621261055
transform 1 0 33696 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_347
timestamp 1621261055
transform 1 0 34464 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_355
timestamp 1621261055
transform 1 0 35232 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_363
timestamp 1621261055
transform 1 0 36000 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_317
timestamp 1621261055
transform 1 0 38112 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_371
timestamp 1621261055
transform 1 0 36768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_379
timestamp 1621261055
transform 1 0 37536 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_383
timestamp 1621261055
transform 1 0 37920 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_386
timestamp 1621261055
transform 1 0 38208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_394
timestamp 1621261055
transform 1 0 38976 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_396
timestamp 1621261055
transform 1 0 39168 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _038_
timestamp 1621261055
transform -1 0 40320 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _144_
timestamp 1621261055
transform 1 0 39264 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_67
timestamp 1621261055
transform -1 0 40032 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_400
timestamp 1621261055
transform 1 0 39552 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_402
timestamp 1621261055
transform 1 0 39744 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_408
timestamp 1621261055
transform 1 0 40320 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_416
timestamp 1621261055
transform 1 0 41088 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_424
timestamp 1621261055
transform 1 0 41856 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_318
timestamp 1621261055
transform 1 0 43392 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_432
timestamp 1621261055
transform 1 0 42624 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_441
timestamp 1621261055
transform 1 0 43488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_449
timestamp 1621261055
transform 1 0 44256 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_457
timestamp 1621261055
transform 1 0 45024 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_319
timestamp 1621261055
transform 1 0 48672 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_465
timestamp 1621261055
transform 1 0 45792 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_473
timestamp 1621261055
transform 1 0 46560 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_481
timestamp 1621261055
transform 1 0 47328 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_489
timestamp 1621261055
transform 1 0 48096 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_493
timestamp 1621261055
transform 1 0 48480 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_496
timestamp 1621261055
transform 1 0 48768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_504
timestamp 1621261055
transform 1 0 49536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_512
timestamp 1621261055
transform 1 0 50304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_520
timestamp 1621261055
transform 1 0 51072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_528
timestamp 1621261055
transform 1 0 51840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_320
timestamp 1621261055
transform 1 0 53952 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_536
timestamp 1621261055
transform 1 0 52608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_544
timestamp 1621261055
transform 1 0 53376 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_548
timestamp 1621261055
transform 1 0 53760 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_551
timestamp 1621261055
transform 1 0 54048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_559
timestamp 1621261055
transform 1 0 54816 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output467
timestamp 1621261055
transform -1 0 57504 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output474
timestamp 1621261055
transform -1 0 56736 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_90
timestamp 1621261055
transform -1 0 57120 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_100
timestamp 1621261055
transform -1 0 56352 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_567
timestamp 1621261055
transform 1 0 55584 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_571
timestamp 1621261055
transform 1 0 55968 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_579
timestamp 1621261055
transform 1 0 56736 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_587
timestamp 1621261055
transform 1 0 57504 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_27
timestamp 1621261055
transform -1 0 58848 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_595
timestamp 1621261055
transform 1 0 58272 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_28
timestamp 1621261055
transform 1 0 1152 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_321
timestamp 1621261055
transform 1 0 3840 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_4
timestamp 1621261055
transform 1 0 1536 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_12
timestamp 1621261055
transform 1 0 2304 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_20
timestamp 1621261055
transform 1 0 3072 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_29
timestamp 1621261055
transform 1 0 3936 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_37
timestamp 1621261055
transform 1 0 4704 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_45
timestamp 1621261055
transform 1 0 5472 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_53
timestamp 1621261055
transform 1 0 6240 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_61
timestamp 1621261055
transform 1 0 7008 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _048_
timestamp 1621261055
transform 1 0 9696 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_322
timestamp 1621261055
transform 1 0 9120 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_44
timestamp 1621261055
transform 1 0 9504 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_69
timestamp 1621261055
transform 1 0 7776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_77
timestamp 1621261055
transform 1 0 8544 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_81
timestamp 1621261055
transform 1 0 8928 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_84
timestamp 1621261055
transform 1 0 9216 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_86
timestamp 1621261055
transform 1 0 9408 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_92
timestamp 1621261055
transform 1 0 9984 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_100
timestamp 1621261055
transform 1 0 10752 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_108
timestamp 1621261055
transform 1 0 11520 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_116
timestamp 1621261055
transform 1 0 12288 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_124
timestamp 1621261055
transform 1 0 13056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_132
timestamp 1621261055
transform 1 0 13824 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_323
timestamp 1621261055
transform 1 0 14400 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_136
timestamp 1621261055
transform 1 0 14208 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_139
timestamp 1621261055
transform 1 0 14496 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_147
timestamp 1621261055
transform 1 0 15264 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_155
timestamp 1621261055
transform 1 0 16032 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_163
timestamp 1621261055
transform 1 0 16800 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_324
timestamp 1621261055
transform 1 0 19680 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_171
timestamp 1621261055
transform 1 0 17568 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_179
timestamp 1621261055
transform 1 0 18336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_187
timestamp 1621261055
transform 1 0 19104 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_191
timestamp 1621261055
transform 1 0 19488 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_194
timestamp 1621261055
transform 1 0 19776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _054_
timestamp 1621261055
transform 1 0 20832 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_62
timestamp 1621261055
transform 1 0 20640 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_202
timestamp 1621261055
transform 1 0 20544 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_208
timestamp 1621261055
transform 1 0 21120 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_216
timestamp 1621261055
transform 1 0 21888 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_224
timestamp 1621261055
transform 1 0 22656 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_325
timestamp 1621261055
transform 1 0 24960 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_232
timestamp 1621261055
transform 1 0 23424 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_240
timestamp 1621261055
transform 1 0 24192 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_249
timestamp 1621261055
transform 1 0 25056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_257
timestamp 1621261055
transform 1 0 25824 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _059_
timestamp 1621261055
transform 1 0 29568 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_14_265
timestamp 1621261055
transform 1 0 26592 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_273
timestamp 1621261055
transform 1 0 27360 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_281
timestamp 1621261055
transform 1 0 28128 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_289
timestamp 1621261055
transform 1 0 28896 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_293
timestamp 1621261055
transform 1 0 29280 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_295
timestamp 1621261055
transform 1 0 29472 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_326
timestamp 1621261055
transform 1 0 30240 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_299
timestamp 1621261055
transform 1 0 29856 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_304
timestamp 1621261055
transform 1 0 30336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_312
timestamp 1621261055
transform 1 0 31104 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_320
timestamp 1621261055
transform 1 0 31872 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_328
timestamp 1621261055
transform 1 0 32640 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_327
timestamp 1621261055
transform 1 0 35520 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_336
timestamp 1621261055
transform 1 0 33408 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_344
timestamp 1621261055
transform 1 0 34176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_352
timestamp 1621261055
transform 1 0 34944 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_356
timestamp 1621261055
transform 1 0 35328 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_359
timestamp 1621261055
transform 1 0 35616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_367
timestamp 1621261055
transform 1 0 36384 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_375
timestamp 1621261055
transform 1 0 37152 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_383
timestamp 1621261055
transform 1 0 37920 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_391
timestamp 1621261055
transform 1 0 38688 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_328
timestamp 1621261055
transform 1 0 40800 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_399
timestamp 1621261055
transform 1 0 39456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_407
timestamp 1621261055
transform 1 0 40224 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_411
timestamp 1621261055
transform 1 0 40608 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_414
timestamp 1621261055
transform 1 0 40896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_422
timestamp 1621261055
transform 1 0 41664 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_430
timestamp 1621261055
transform 1 0 42432 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_438
timestamp 1621261055
transform 1 0 43200 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_446
timestamp 1621261055
transform 1 0 43968 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_454
timestamp 1621261055
transform 1 0 44736 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_462
timestamp 1621261055
transform 1 0 45504 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_329
timestamp 1621261055
transform 1 0 46080 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_466
timestamp 1621261055
transform 1 0 45888 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_469
timestamp 1621261055
transform 1 0 46176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_477
timestamp 1621261055
transform 1 0 46944 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_485
timestamp 1621261055
transform 1 0 47712 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_493
timestamp 1621261055
transform 1 0 48480 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_330
timestamp 1621261055
transform 1 0 51360 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_501
timestamp 1621261055
transform 1 0 49248 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_509
timestamp 1621261055
transform 1 0 50016 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_517
timestamp 1621261055
transform 1 0 50784 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_521
timestamp 1621261055
transform 1 0 51168 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_524
timestamp 1621261055
transform 1 0 51456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_532
timestamp 1621261055
transform 1 0 52224 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_540
timestamp 1621261055
transform 1 0 52992 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_548
timestamp 1621261055
transform 1 0 53760 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_556
timestamp 1621261055
transform 1 0 54528 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_331
timestamp 1621261055
transform 1 0 56640 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output468
timestamp 1621261055
transform -1 0 57888 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_92
timestamp 1621261055
transform -1 0 57504 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_564
timestamp 1621261055
transform 1 0 55296 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_572
timestamp 1621261055
transform 1 0 56064 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_576
timestamp 1621261055
transform 1 0 56448 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_579
timestamp 1621261055
transform 1 0 56736 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_583
timestamp 1621261055
transform 1 0 57120 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_591
timestamp 1621261055
transform 1 0 57888 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_29
timestamp 1621261055
transform -1 0 58848 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_595
timestamp 1621261055
transform 1 0 58272 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_4
timestamp 1621261055
transform 1 0 1536 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_4
timestamp 1621261055
transform 1 0 1536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_32
timestamp 1621261055
transform 1 0 1152 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_30
timestamp 1621261055
transform 1 0 1152 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_12
timestamp 1621261055
transform 1 0 2304 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_12
timestamp 1621261055
transform 1 0 2304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_20
timestamp 1621261055
transform 1 0 3072 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_20
timestamp 1621261055
transform 1 0 3072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_29
timestamp 1621261055
transform 1 0 3936 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_28
timestamp 1621261055
transform 1 0 3840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_342
timestamp 1621261055
transform 1 0 3840 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_16_37
timestamp 1621261055
transform 1 0 4704 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_36
timestamp 1621261055
transform 1 0 4608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _187_
timestamp 1621261055
transform 1 0 5088 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_44
timestamp 1621261055
transform 1 0 5376 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_44
timestamp 1621261055
transform 1 0 5376 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_52
timestamp 1621261055
transform 1 0 6144 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_56
timestamp 1621261055
transform 1 0 6528 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_54
timestamp 1621261055
transform 1 0 6336 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_52
timestamp 1621261055
transform 1 0 6144 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_332
timestamp 1621261055
transform 1 0 6432 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_60
timestamp 1621261055
transform 1 0 6912 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_64
timestamp 1621261055
transform 1 0 7296 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_68
timestamp 1621261055
transform 1 0 7680 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_72
timestamp 1621261055
transform 1 0 8064 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_82
timestamp 1621261055
transform 1 0 9024 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_80
timestamp 1621261055
transform 1 0 8832 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_76
timestamp 1621261055
transform 1 0 8448 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_15_80
timestamp 1621261055
transform 1 0 8832 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_343
timestamp 1621261055
transform 1 0 9120 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_92
timestamp 1621261055
transform 1 0 9984 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_84
timestamp 1621261055
transform 1 0 9216 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_90
timestamp 1621261055
transform 1 0 9792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_86
timestamp 1621261055
transform 1 0 9408 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_84
timestamp 1621261055
transform 1 0 9216 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _138_
timestamp 1621261055
transform 1 0 9504 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_15_98
timestamp 1621261055
transform 1 0 10560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_100
timestamp 1621261055
transform 1 0 10752 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_106
timestamp 1621261055
transform 1 0 11328 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_108
timestamp 1621261055
transform 1 0 11520 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_111
timestamp 1621261055
transform 1 0 11808 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_49
timestamp 1621261055
transform -1 0 12480 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_333
timestamp 1621261055
transform 1 0 11712 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_124
timestamp 1621261055
transform 1 0 13056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_119
timestamp 1621261055
transform 1 0 12576 0 1 12654
box -38 -49 806 715
use INV  INV
timestamp 1623610208
transform -1 0 13056 0 -1 13986
box 0 -48 576 714
use sky130_fd_sc_ls__decap_4  FILLER_16_132
timestamp 1621261055
transform 1 0 13824 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_127
timestamp 1621261055
transform 1 0 13344 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_139
timestamp 1621261055
transform 1 0 14496 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_136
timestamp 1621261055
transform 1 0 14208 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_135
timestamp 1621261055
transform 1 0 14112 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_344
timestamp 1621261055
transform 1 0 14400 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_147
timestamp 1621261055
transform 1 0 15264 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_143
timestamp 1621261055
transform 1 0 14880 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_155
timestamp 1621261055
transform 1 0 16032 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_151
timestamp 1621261055
transform 1 0 15648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_163
timestamp 1621261055
transform 1 0 16800 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_163
timestamp 1621261055
transform 1 0 16800 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_159
timestamp 1621261055
transform 1 0 16416 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_334
timestamp 1621261055
transform 1 0 16992 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_171
timestamp 1621261055
transform 1 0 17568 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_166
timestamp 1621261055
transform 1 0 17088 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_179
timestamp 1621261055
transform 1 0 18336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_182
timestamp 1621261055
transform 1 0 18624 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_174
timestamp 1621261055
transform 1 0 17856 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_191
timestamp 1621261055
transform 1 0 19488 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_187
timestamp 1621261055
transform 1 0 19104 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_190
timestamp 1621261055
transform 1 0 19392 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_194
timestamp 1621261055
transform 1 0 19776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_198
timestamp 1621261055
transform 1 0 20160 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_345
timestamp 1621261055
transform 1 0 19680 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_202
timestamp 1621261055
transform 1 0 20544 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_206
timestamp 1621261055
transform 1 0 20928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_210
timestamp 1621261055
transform 1 0 21312 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_214
timestamp 1621261055
transform 1 0 21696 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_218
timestamp 1621261055
transform 1 0 22080 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_221
timestamp 1621261055
transform 1 0 22368 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_218
timestamp 1621261055
transform 1 0 22080 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_335
timestamp 1621261055
transform 1 0 22272 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_226
timestamp 1621261055
transform 1 0 22848 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_229
timestamp 1621261055
transform 1 0 23136 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_234
timestamp 1621261055
transform 1 0 23616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_237
timestamp 1621261055
transform 1 0 23904 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_246
timestamp 1621261055
transform 1 0 24768 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_242
timestamp 1621261055
transform 1 0 24384 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_245
timestamp 1621261055
transform 1 0 24672 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_346
timestamp 1621261055
transform 1 0 24960 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_257
timestamp 1621261055
transform 1 0 25824 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_249
timestamp 1621261055
transform 1 0 25056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_253
timestamp 1621261055
transform 1 0 25440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_261
timestamp 1621261055
transform 1 0 26208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_265
timestamp 1621261055
transform 1 0 26592 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_269
timestamp 1621261055
transform 1 0 26976 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_281
timestamp 1621261055
transform 1 0 28128 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_273
timestamp 1621261055
transform 1 0 27360 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_276
timestamp 1621261055
transform 1 0 27648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_273
timestamp 1621261055
transform 1 0 27360 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_336
timestamp 1621261055
transform 1 0 27552 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_289
timestamp 1621261055
transform 1 0 28896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_284
timestamp 1621261055
transform 1 0 28416 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_297
timestamp 1621261055
transform 1 0 29664 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_15_296
timestamp 1621261055
transform 1 0 29568 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_292
timestamp 1621261055
transform 1 0 29184 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _085_
timestamp 1621261055
transform 1 0 29664 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_304
timestamp 1621261055
transform 1 0 30336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_301
timestamp 1621261055
transform 1 0 30048 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_300
timestamp 1621261055
transform 1 0 29952 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_347
timestamp 1621261055
transform 1 0 30240 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_312
timestamp 1621261055
transform 1 0 31104 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_308
timestamp 1621261055
transform 1 0 30720 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_320
timestamp 1621261055
transform 1 0 31872 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_316
timestamp 1621261055
transform 1 0 31488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_328
timestamp 1621261055
transform 1 0 32640 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_328
timestamp 1621261055
transform 1 0 32640 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_324
timestamp 1621261055
transform 1 0 32256 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_337
timestamp 1621261055
transform 1 0 32832 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_336
timestamp 1621261055
transform 1 0 33408 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_331
timestamp 1621261055
transform 1 0 32928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_344
timestamp 1621261055
transform 1 0 34176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_347
timestamp 1621261055
transform 1 0 34464 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_339
timestamp 1621261055
transform 1 0 33696 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_356
timestamp 1621261055
transform 1 0 35328 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_352
timestamp 1621261055
transform 1 0 34944 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_355
timestamp 1621261055
transform 1 0 35232 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_359
timestamp 1621261055
transform 1 0 35616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_363
timestamp 1621261055
transform 1 0 36000 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_348
timestamp 1621261055
transform 1 0 35520 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_367
timestamp 1621261055
transform 1 0 36384 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_371
timestamp 1621261055
transform 1 0 36768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_375
timestamp 1621261055
transform 1 0 37152 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_379
timestamp 1621261055
transform 1 0 37536 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_383
timestamp 1621261055
transform 1 0 37920 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_386
timestamp 1621261055
transform 1 0 38208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_383
timestamp 1621261055
transform 1 0 37920 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_338
timestamp 1621261055
transform 1 0 38112 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_391
timestamp 1621261055
transform 1 0 38688 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_394
timestamp 1621261055
transform 1 0 38976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_399
timestamp 1621261055
transform 1 0 39456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_402
timestamp 1621261055
transform 1 0 39744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_411
timestamp 1621261055
transform 1 0 40608 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_407
timestamp 1621261055
transform 1 0 40224 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_410
timestamp 1621261055
transform 1 0 40512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_349
timestamp 1621261055
transform 1 0 40800 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_422
timestamp 1621261055
transform 1 0 41664 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_414
timestamp 1621261055
transform 1 0 40896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_418
timestamp 1621261055
transform 1 0 41280 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_426
timestamp 1621261055
transform 1 0 42048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_430
timestamp 1621261055
transform 1 0 42432 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_434
timestamp 1621261055
transform 1 0 42816 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_446
timestamp 1621261055
transform 1 0 43968 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_438
timestamp 1621261055
transform 1 0 43200 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_441
timestamp 1621261055
transform 1 0 43488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_438
timestamp 1621261055
transform 1 0 43200 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_339
timestamp 1621261055
transform 1 0 43392 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_454
timestamp 1621261055
transform 1 0 44736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_449
timestamp 1621261055
transform 1 0 44256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_462
timestamp 1621261055
transform 1 0 45504 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_457
timestamp 1621261055
transform 1 0 45024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_469
timestamp 1621261055
transform 1 0 46176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_466
timestamp 1621261055
transform 1 0 45888 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_465
timestamp 1621261055
transform 1 0 45792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_350
timestamp 1621261055
transform 1 0 46080 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_477
timestamp 1621261055
transform 1 0 46944 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_473
timestamp 1621261055
transform 1 0 46560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_485
timestamp 1621261055
transform 1 0 47712 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_481
timestamp 1621261055
transform 1 0 47328 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_493
timestamp 1621261055
transform 1 0 48480 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_493
timestamp 1621261055
transform 1 0 48480 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_489
timestamp 1621261055
transform 1 0 48096 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_340
timestamp 1621261055
transform 1 0 48672 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_501
timestamp 1621261055
transform 1 0 49248 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_503
timestamp 1621261055
transform 1 0 49440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_496
timestamp 1621261055
transform 1 0 48768 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _152_
timestamp 1621261055
transform 1 0 49152 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_509
timestamp 1621261055
transform 1 0 50016 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_511
timestamp 1621261055
transform 1 0 50208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_521
timestamp 1621261055
transform 1 0 51168 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_517
timestamp 1621261055
transform 1 0 50784 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_519
timestamp 1621261055
transform 1 0 50976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_524
timestamp 1621261055
transform 1 0 51456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_527
timestamp 1621261055
transform 1 0 51744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_351
timestamp 1621261055
transform 1 0 51360 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_532
timestamp 1621261055
transform 1 0 52224 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_535
timestamp 1621261055
transform 1 0 52512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_540
timestamp 1621261055
transform 1 0 52992 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_543
timestamp 1621261055
transform 1 0 53280 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_548
timestamp 1621261055
transform 1 0 53760 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_551
timestamp 1621261055
transform 1 0 54048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_549
timestamp 1621261055
transform 1 0 53856 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_547
timestamp 1621261055
transform 1 0 53664 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_341
timestamp 1621261055
transform 1 0 53952 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_556
timestamp 1621261055
transform 1 0 54528 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_559
timestamp 1621261055
transform 1 0 54816 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_564
timestamp 1621261055
transform 1 0 55296 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_567
timestamp 1621261055
transform 1 0 55584 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_576
timestamp 1621261055
transform 1 0 56448 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_572
timestamp 1621261055
transform 1 0 56064 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_575
timestamp 1621261055
transform 1 0 56352 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_352
timestamp 1621261055
transform 1 0 56640 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_587
timestamp 1621261055
transform 1 0 57504 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_579
timestamp 1621261055
transform 1 0 56736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_587
timestamp 1621261055
transform 1 0 57504 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_583
timestamp 1621261055
transform 1 0 57120 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_15_593
timestamp 1621261055
transform 1 0 58080 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_23
timestamp 1621261055
transform -1 0 57792 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _033_
timestamp 1621261055
transform -1 0 58080 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_31
timestamp 1621261055
transform -1 0 58848 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_33
timestamp 1621261055
transform -1 0 58848 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_595
timestamp 1621261055
transform 1 0 58272 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_34
timestamp 1621261055
transform 1 0 1152 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_4
timestamp 1621261055
transform 1 0 1536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_12
timestamp 1621261055
transform 1 0 2304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_20
timestamp 1621261055
transform 1 0 3072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_28
timestamp 1621261055
transform 1 0 3840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_353
timestamp 1621261055
transform 1 0 6432 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_36
timestamp 1621261055
transform 1 0 4608 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_44
timestamp 1621261055
transform 1 0 5376 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_52
timestamp 1621261055
transform 1 0 6144 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_54
timestamp 1621261055
transform 1 0 6336 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_56
timestamp 1621261055
transform 1 0 6528 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_64
timestamp 1621261055
transform 1 0 7296 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_72
timestamp 1621261055
transform 1 0 8064 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_80
timestamp 1621261055
transform 1 0 8832 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_88
timestamp 1621261055
transform 1 0 9600 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_96
timestamp 1621261055
transform 1 0 10368 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_354
timestamp 1621261055
transform 1 0 11712 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_104
timestamp 1621261055
transform 1 0 11136 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_108
timestamp 1621261055
transform 1 0 11520 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_111
timestamp 1621261055
transform 1 0 11808 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_119
timestamp 1621261055
transform 1 0 12576 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_127
timestamp 1621261055
transform 1 0 13344 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_355
timestamp 1621261055
transform 1 0 16992 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_135
timestamp 1621261055
transform 1 0 14112 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_143
timestamp 1621261055
transform 1 0 14880 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_151
timestamp 1621261055
transform 1 0 15648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_159
timestamp 1621261055
transform 1 0 16416 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_163
timestamp 1621261055
transform 1 0 16800 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_166
timestamp 1621261055
transform 1 0 17088 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_174
timestamp 1621261055
transform 1 0 17856 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_182
timestamp 1621261055
transform 1 0 18624 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_190
timestamp 1621261055
transform 1 0 19392 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_198
timestamp 1621261055
transform 1 0 20160 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_356
timestamp 1621261055
transform 1 0 22272 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_206
timestamp 1621261055
transform 1 0 20928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_214
timestamp 1621261055
transform 1 0 21696 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_218
timestamp 1621261055
transform 1 0 22080 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_221
timestamp 1621261055
transform 1 0 22368 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_229
timestamp 1621261055
transform 1 0 23136 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_237
timestamp 1621261055
transform 1 0 23904 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_245
timestamp 1621261055
transform 1 0 24672 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_253
timestamp 1621261055
transform 1 0 25440 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_261
timestamp 1621261055
transform 1 0 26208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_357
timestamp 1621261055
transform 1 0 27552 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_269
timestamp 1621261055
transform 1 0 26976 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_273
timestamp 1621261055
transform 1 0 27360 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_276
timestamp 1621261055
transform 1 0 27648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_284
timestamp 1621261055
transform 1 0 28416 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_292
timestamp 1621261055
transform 1 0 29184 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_358
timestamp 1621261055
transform 1 0 32832 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_300
timestamp 1621261055
transform 1 0 29952 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_308
timestamp 1621261055
transform 1 0 30720 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_316
timestamp 1621261055
transform 1 0 31488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_324
timestamp 1621261055
transform 1 0 32256 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_328
timestamp 1621261055
transform 1 0 32640 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_331
timestamp 1621261055
transform 1 0 32928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_339
timestamp 1621261055
transform 1 0 33696 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_347
timestamp 1621261055
transform 1 0 34464 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_355
timestamp 1621261055
transform 1 0 35232 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_363
timestamp 1621261055
transform 1 0 36000 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_359
timestamp 1621261055
transform 1 0 38112 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_371
timestamp 1621261055
transform 1 0 36768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_379
timestamp 1621261055
transform 1 0 37536 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_383
timestamp 1621261055
transform 1 0 37920 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_386
timestamp 1621261055
transform 1 0 38208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_394
timestamp 1621261055
transform 1 0 38976 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_402
timestamp 1621261055
transform 1 0 39744 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_410
timestamp 1621261055
transform 1 0 40512 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_418
timestamp 1621261055
transform 1 0 41280 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_426
timestamp 1621261055
transform 1 0 42048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _019_
timestamp 1621261055
transform 1 0 44832 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_360
timestamp 1621261055
transform 1 0 43392 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_28
timestamp 1621261055
transform 1 0 44640 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_17_434
timestamp 1621261055
transform 1 0 42816 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_438
timestamp 1621261055
transform 1 0 43200 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_441
timestamp 1621261055
transform 1 0 43488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_449
timestamp 1621261055
transform 1 0 44256 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_458
timestamp 1621261055
transform 1 0 45120 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _207_
timestamp 1621261055
transform 1 0 46368 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_361
timestamp 1621261055
transform 1 0 48672 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_466
timestamp 1621261055
transform 1 0 45888 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_17_470
timestamp 1621261055
transform 1 0 46272 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_474
timestamp 1621261055
transform 1 0 46656 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_482
timestamp 1621261055
transform 1 0 47424 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_490
timestamp 1621261055
transform 1 0 48192 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_17_494
timestamp 1621261055
transform 1 0 48576 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _031_
timestamp 1621261055
transform -1 0 49440 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_14
timestamp 1621261055
transform -1 0 49152 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_496
timestamp 1621261055
transform 1 0 48768 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_503
timestamp 1621261055
transform 1 0 49440 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_511
timestamp 1621261055
transform 1 0 50208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_519
timestamp 1621261055
transform 1 0 50976 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_527
timestamp 1621261055
transform 1 0 51744 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_362
timestamp 1621261055
transform 1 0 53952 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_535
timestamp 1621261055
transform 1 0 52512 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_543
timestamp 1621261055
transform 1 0 53280 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_547
timestamp 1621261055
transform 1 0 53664 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_549
timestamp 1621261055
transform 1 0 53856 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_551
timestamp 1621261055
transform 1 0 54048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_559
timestamp 1621261055
transform 1 0 54816 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_567
timestamp 1621261055
transform 1 0 55584 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_575
timestamp 1621261055
transform 1 0 56352 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_583
timestamp 1621261055
transform 1 0 57120 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_591
timestamp 1621261055
transform 1 0 57888 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_35
timestamp 1621261055
transform -1 0 58848 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_595
timestamp 1621261055
transform 1 0 58272 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_36
timestamp 1621261055
transform 1 0 1152 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_363
timestamp 1621261055
transform 1 0 3840 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_4
timestamp 1621261055
transform 1 0 1536 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_12
timestamp 1621261055
transform 1 0 2304 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_20
timestamp 1621261055
transform 1 0 3072 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_29
timestamp 1621261055
transform 1 0 3936 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_37
timestamp 1621261055
transform 1 0 4704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_45
timestamp 1621261055
transform 1 0 5472 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_53
timestamp 1621261055
transform 1 0 6240 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_61
timestamp 1621261055
transform 1 0 7008 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_364
timestamp 1621261055
transform 1 0 9120 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_69
timestamp 1621261055
transform 1 0 7776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_77
timestamp 1621261055
transform 1 0 8544 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_81
timestamp 1621261055
transform 1 0 8928 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_84
timestamp 1621261055
transform 1 0 9216 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_92
timestamp 1621261055
transform 1 0 9984 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_100
timestamp 1621261055
transform 1 0 10752 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_108
timestamp 1621261055
transform 1 0 11520 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_116
timestamp 1621261055
transform 1 0 12288 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_124
timestamp 1621261055
transform 1 0 13056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_132
timestamp 1621261055
transform 1 0 13824 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_365
timestamp 1621261055
transform 1 0 14400 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_136
timestamp 1621261055
transform 1 0 14208 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_139
timestamp 1621261055
transform 1 0 14496 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_147
timestamp 1621261055
transform 1 0 15264 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_155
timestamp 1621261055
transform 1 0 16032 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_163
timestamp 1621261055
transform 1 0 16800 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_366
timestamp 1621261055
transform 1 0 19680 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_171
timestamp 1621261055
transform 1 0 17568 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_179
timestamp 1621261055
transform 1 0 18336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_187
timestamp 1621261055
transform 1 0 19104 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_191
timestamp 1621261055
transform 1 0 19488 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_194
timestamp 1621261055
transform 1 0 19776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_202
timestamp 1621261055
transform 1 0 20544 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_210
timestamp 1621261055
transform 1 0 21312 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_218
timestamp 1621261055
transform 1 0 22080 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_226
timestamp 1621261055
transform 1 0 22848 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_367
timestamp 1621261055
transform 1 0 24960 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_234
timestamp 1621261055
transform 1 0 23616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_242
timestamp 1621261055
transform 1 0 24384 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_246
timestamp 1621261055
transform 1 0 24768 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_249
timestamp 1621261055
transform 1 0 25056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_257
timestamp 1621261055
transform 1 0 25824 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_265
timestamp 1621261055
transform 1 0 26592 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_273
timestamp 1621261055
transform 1 0 27360 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_281
timestamp 1621261055
transform 1 0 28128 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_289
timestamp 1621261055
transform 1 0 28896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_297
timestamp 1621261055
transform 1 0 29664 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _099_
timestamp 1621261055
transform 1 0 32064 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_368
timestamp 1621261055
transform 1 0 30240 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_301
timestamp 1621261055
transform 1 0 30048 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_304
timestamp 1621261055
transform 1 0 30336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_312
timestamp 1621261055
transform 1 0 31104 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_320
timestamp 1621261055
transform 1 0 31872 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_325
timestamp 1621261055
transform 1 0 32352 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_369
timestamp 1621261055
transform 1 0 35520 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_333
timestamp 1621261055
transform 1 0 33120 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_341
timestamp 1621261055
transform 1 0 33888 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_349
timestamp 1621261055
transform 1 0 34656 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_18_357
timestamp 1621261055
transform 1 0 35424 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_359
timestamp 1621261055
transform 1 0 35616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_367
timestamp 1621261055
transform 1 0 36384 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_375
timestamp 1621261055
transform 1 0 37152 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_383
timestamp 1621261055
transform 1 0 37920 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_391
timestamp 1621261055
transform 1 0 38688 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_370
timestamp 1621261055
transform 1 0 40800 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_399
timestamp 1621261055
transform 1 0 39456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_407
timestamp 1621261055
transform 1 0 40224 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_411
timestamp 1621261055
transform 1 0 40608 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_414
timestamp 1621261055
transform 1 0 40896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_422
timestamp 1621261055
transform 1 0 41664 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_430
timestamp 1621261055
transform 1 0 42432 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_438
timestamp 1621261055
transform 1 0 43200 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_446
timestamp 1621261055
transform 1 0 43968 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_454
timestamp 1621261055
transform 1 0 44736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_462
timestamp 1621261055
transform 1 0 45504 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_371
timestamp 1621261055
transform 1 0 46080 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_466
timestamp 1621261055
transform 1 0 45888 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_469
timestamp 1621261055
transform 1 0 46176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_477
timestamp 1621261055
transform 1 0 46944 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_485
timestamp 1621261055
transform 1 0 47712 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_493
timestamp 1621261055
transform 1 0 48480 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_372
timestamp 1621261055
transform 1 0 51360 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_501
timestamp 1621261055
transform 1 0 49248 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_509
timestamp 1621261055
transform 1 0 50016 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_517
timestamp 1621261055
transform 1 0 50784 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_521
timestamp 1621261055
transform 1 0 51168 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_524
timestamp 1621261055
transform 1 0 51456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_532
timestamp 1621261055
transform 1 0 52224 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_540
timestamp 1621261055
transform 1 0 52992 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_548
timestamp 1621261055
transform 1 0 53760 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_556
timestamp 1621261055
transform 1 0 54528 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_373
timestamp 1621261055
transform 1 0 56640 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_564
timestamp 1621261055
transform 1 0 55296 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_572
timestamp 1621261055
transform 1 0 56064 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_576
timestamp 1621261055
transform 1 0 56448 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_579
timestamp 1621261055
transform 1 0 56736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_587
timestamp 1621261055
transform 1 0 57504 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_37
timestamp 1621261055
transform -1 0 58848 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_595
timestamp 1621261055
transform 1 0 58272 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_38
timestamp 1621261055
transform 1 0 1152 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_4
timestamp 1621261055
transform 1 0 1536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_12
timestamp 1621261055
transform 1 0 2304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_20
timestamp 1621261055
transform 1 0 3072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_28
timestamp 1621261055
transform 1 0 3840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_374
timestamp 1621261055
transform 1 0 6432 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_36
timestamp 1621261055
transform 1 0 4608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_44
timestamp 1621261055
transform 1 0 5376 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_52
timestamp 1621261055
transform 1 0 6144 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_54
timestamp 1621261055
transform 1 0 6336 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_56
timestamp 1621261055
transform 1 0 6528 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_64
timestamp 1621261055
transform 1 0 7296 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _160_
timestamp 1621261055
transform 1 0 9600 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_19_72
timestamp 1621261055
transform 1 0 8064 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_80
timestamp 1621261055
transform 1 0 8832 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_91
timestamp 1621261055
transform 1 0 9888 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_99
timestamp 1621261055
transform 1 0 10656 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_375
timestamp 1621261055
transform 1 0 11712 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_107
timestamp 1621261055
transform 1 0 11424 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_109
timestamp 1621261055
transform 1 0 11616 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_111
timestamp 1621261055
transform 1 0 11808 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_119
timestamp 1621261055
transform 1 0 12576 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_127
timestamp 1621261055
transform 1 0 13344 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_376
timestamp 1621261055
transform 1 0 16992 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_135
timestamp 1621261055
transform 1 0 14112 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_143
timestamp 1621261055
transform 1 0 14880 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_151
timestamp 1621261055
transform 1 0 15648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_159
timestamp 1621261055
transform 1 0 16416 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_163
timestamp 1621261055
transform 1 0 16800 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_166
timestamp 1621261055
transform 1 0 17088 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_174
timestamp 1621261055
transform 1 0 17856 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_182
timestamp 1621261055
transform 1 0 18624 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_190
timestamp 1621261055
transform 1 0 19392 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_198
timestamp 1621261055
transform 1 0 20160 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_377
timestamp 1621261055
transform 1 0 22272 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_206
timestamp 1621261055
transform 1 0 20928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_214
timestamp 1621261055
transform 1 0 21696 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_218
timestamp 1621261055
transform 1 0 22080 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_221
timestamp 1621261055
transform 1 0 22368 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_229
timestamp 1621261055
transform 1 0 23136 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_237
timestamp 1621261055
transform 1 0 23904 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_245
timestamp 1621261055
transform 1 0 24672 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_253
timestamp 1621261055
transform 1 0 25440 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_261
timestamp 1621261055
transform 1 0 26208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_378
timestamp 1621261055
transform 1 0 27552 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_269
timestamp 1621261055
transform 1 0 26976 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_273
timestamp 1621261055
transform 1 0 27360 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_276
timestamp 1621261055
transform 1 0 27648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_284
timestamp 1621261055
transform 1 0 28416 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_292
timestamp 1621261055
transform 1 0 29184 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_379
timestamp 1621261055
transform 1 0 32832 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_300
timestamp 1621261055
transform 1 0 29952 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_308
timestamp 1621261055
transform 1 0 30720 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_316
timestamp 1621261055
transform 1 0 31488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_324
timestamp 1621261055
transform 1 0 32256 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_328
timestamp 1621261055
transform 1 0 32640 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_331
timestamp 1621261055
transform 1 0 32928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_339
timestamp 1621261055
transform 1 0 33696 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_347
timestamp 1621261055
transform 1 0 34464 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_355
timestamp 1621261055
transform 1 0 35232 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_363
timestamp 1621261055
transform 1 0 36000 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_380
timestamp 1621261055
transform 1 0 38112 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_371
timestamp 1621261055
transform 1 0 36768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_379
timestamp 1621261055
transform 1 0 37536 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_383
timestamp 1621261055
transform 1 0 37920 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_386
timestamp 1621261055
transform 1 0 38208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_394
timestamp 1621261055
transform 1 0 38976 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_402
timestamp 1621261055
transform 1 0 39744 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_410
timestamp 1621261055
transform 1 0 40512 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_418
timestamp 1621261055
transform 1 0 41280 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_426
timestamp 1621261055
transform 1 0 42048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_381
timestamp 1621261055
transform 1 0 43392 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_434
timestamp 1621261055
transform 1 0 42816 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_438
timestamp 1621261055
transform 1 0 43200 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_441
timestamp 1621261055
transform 1 0 43488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_449
timestamp 1621261055
transform 1 0 44256 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_457
timestamp 1621261055
transform 1 0 45024 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_382
timestamp 1621261055
transform 1 0 48672 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_465
timestamp 1621261055
transform 1 0 45792 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_473
timestamp 1621261055
transform 1 0 46560 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_481
timestamp 1621261055
transform 1 0 47328 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_489
timestamp 1621261055
transform 1 0 48096 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_493
timestamp 1621261055
transform 1 0 48480 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_496
timestamp 1621261055
transform 1 0 48768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_504
timestamp 1621261055
transform 1 0 49536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_512
timestamp 1621261055
transform 1 0 50304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_520
timestamp 1621261055
transform 1 0 51072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_528
timestamp 1621261055
transform 1 0 51840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_383
timestamp 1621261055
transform 1 0 53952 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_536
timestamp 1621261055
transform 1 0 52608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_544
timestamp 1621261055
transform 1 0 53376 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_548
timestamp 1621261055
transform 1 0 53760 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_551
timestamp 1621261055
transform 1 0 54048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_559
timestamp 1621261055
transform 1 0 54816 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_567
timestamp 1621261055
transform 1 0 55584 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_575
timestamp 1621261055
transform 1 0 56352 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_583
timestamp 1621261055
transform 1 0 57120 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_591
timestamp 1621261055
transform 1 0 57888 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_39
timestamp 1621261055
transform -1 0 58848 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_595
timestamp 1621261055
transform 1 0 58272 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_40
timestamp 1621261055
transform 1 0 1152 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_384
timestamp 1621261055
transform 1 0 3840 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_4
timestamp 1621261055
transform 1 0 1536 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_12
timestamp 1621261055
transform 1 0 2304 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_20
timestamp 1621261055
transform 1 0 3072 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_29
timestamp 1621261055
transform 1 0 3936 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_37
timestamp 1621261055
transform 1 0 4704 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_45
timestamp 1621261055
transform 1 0 5472 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_53
timestamp 1621261055
transform 1 0 6240 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_61
timestamp 1621261055
transform 1 0 7008 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_385
timestamp 1621261055
transform 1 0 9120 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_69
timestamp 1621261055
transform 1 0 7776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_77
timestamp 1621261055
transform 1 0 8544 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_81
timestamp 1621261055
transform 1 0 8928 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_84
timestamp 1621261055
transform 1 0 9216 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_92
timestamp 1621261055
transform 1 0 9984 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_100
timestamp 1621261055
transform 1 0 10752 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_108
timestamp 1621261055
transform 1 0 11520 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_116
timestamp 1621261055
transform 1 0 12288 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_124
timestamp 1621261055
transform 1 0 13056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_132
timestamp 1621261055
transform 1 0 13824 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_386
timestamp 1621261055
transform 1 0 14400 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_136
timestamp 1621261055
transform 1 0 14208 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_139
timestamp 1621261055
transform 1 0 14496 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_147
timestamp 1621261055
transform 1 0 15264 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_155
timestamp 1621261055
transform 1 0 16032 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_163
timestamp 1621261055
transform 1 0 16800 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_387
timestamp 1621261055
transform 1 0 19680 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_171
timestamp 1621261055
transform 1 0 17568 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_179
timestamp 1621261055
transform 1 0 18336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_187
timestamp 1621261055
transform 1 0 19104 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_191
timestamp 1621261055
transform 1 0 19488 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_194
timestamp 1621261055
transform 1 0 19776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_202
timestamp 1621261055
transform 1 0 20544 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_210
timestamp 1621261055
transform 1 0 21312 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_218
timestamp 1621261055
transform 1 0 22080 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_226
timestamp 1621261055
transform 1 0 22848 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_388
timestamp 1621261055
transform 1 0 24960 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_234
timestamp 1621261055
transform 1 0 23616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_242
timestamp 1621261055
transform 1 0 24384 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_246
timestamp 1621261055
transform 1 0 24768 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_249
timestamp 1621261055
transform 1 0 25056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_257
timestamp 1621261055
transform 1 0 25824 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_265
timestamp 1621261055
transform 1 0 26592 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_273
timestamp 1621261055
transform 1 0 27360 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_281
timestamp 1621261055
transform 1 0 28128 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_289
timestamp 1621261055
transform 1 0 28896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_297
timestamp 1621261055
transform 1 0 29664 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_389
timestamp 1621261055
transform 1 0 30240 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_301
timestamp 1621261055
transform 1 0 30048 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_304
timestamp 1621261055
transform 1 0 30336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_312
timestamp 1621261055
transform 1 0 31104 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_320
timestamp 1621261055
transform 1 0 31872 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_328
timestamp 1621261055
transform 1 0 32640 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_390
timestamp 1621261055
transform 1 0 35520 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_336
timestamp 1621261055
transform 1 0 33408 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_344
timestamp 1621261055
transform 1 0 34176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_352
timestamp 1621261055
transform 1 0 34944 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_356
timestamp 1621261055
transform 1 0 35328 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_359
timestamp 1621261055
transform 1 0 35616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_367
timestamp 1621261055
transform 1 0 36384 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_375
timestamp 1621261055
transform 1 0 37152 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_383
timestamp 1621261055
transform 1 0 37920 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_391
timestamp 1621261055
transform 1 0 38688 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_391
timestamp 1621261055
transform 1 0 40800 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_399
timestamp 1621261055
transform 1 0 39456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_407
timestamp 1621261055
transform 1 0 40224 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_411
timestamp 1621261055
transform 1 0 40608 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_414
timestamp 1621261055
transform 1 0 40896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_422
timestamp 1621261055
transform 1 0 41664 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_430
timestamp 1621261055
transform 1 0 42432 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_438
timestamp 1621261055
transform 1 0 43200 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_446
timestamp 1621261055
transform 1 0 43968 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_454
timestamp 1621261055
transform 1 0 44736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_462
timestamp 1621261055
transform 1 0 45504 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_392
timestamp 1621261055
transform 1 0 46080 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_466
timestamp 1621261055
transform 1 0 45888 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_469
timestamp 1621261055
transform 1 0 46176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_477
timestamp 1621261055
transform 1 0 46944 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_485
timestamp 1621261055
transform 1 0 47712 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_493
timestamp 1621261055
transform 1 0 48480 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_393
timestamp 1621261055
transform 1 0 51360 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_501
timestamp 1621261055
transform 1 0 49248 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_509
timestamp 1621261055
transform 1 0 50016 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_517
timestamp 1621261055
transform 1 0 50784 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_521
timestamp 1621261055
transform 1 0 51168 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_524
timestamp 1621261055
transform 1 0 51456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _023_
timestamp 1621261055
transform 1 0 53472 0 -1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_2
timestamp 1621261055
transform 1 0 53280 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_532
timestamp 1621261055
transform 1 0 52224 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_540
timestamp 1621261055
transform 1 0 52992 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_20_542
timestamp 1621261055
transform 1 0 53184 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_548
timestamp 1621261055
transform 1 0 53760 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_556
timestamp 1621261055
transform 1 0 54528 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_394
timestamp 1621261055
transform 1 0 56640 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_564
timestamp 1621261055
transform 1 0 55296 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_572
timestamp 1621261055
transform 1 0 56064 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_576
timestamp 1621261055
transform 1 0 56448 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_579
timestamp 1621261055
transform 1 0 56736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_587
timestamp 1621261055
transform 1 0 57504 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_41
timestamp 1621261055
transform -1 0 58848 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_595
timestamp 1621261055
transform 1 0 58272 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _049_
timestamp 1621261055
transform 1 0 2880 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_42
timestamp 1621261055
transform 1 0 1152 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_46
timestamp 1621261055
transform 1 0 2688 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_4
timestamp 1621261055
transform 1 0 1536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_12
timestamp 1621261055
transform 1 0 2304 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_21
timestamp 1621261055
transform 1 0 3168 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_29
timestamp 1621261055
transform 1 0 3936 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_395
timestamp 1621261055
transform 1 0 6432 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_37
timestamp 1621261055
transform 1 0 4704 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_45
timestamp 1621261055
transform 1 0 5472 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_53
timestamp 1621261055
transform 1 0 6240 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_56
timestamp 1621261055
transform 1 0 6528 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_64
timestamp 1621261055
transform 1 0 7296 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _074_
timestamp 1621261055
transform 1 0 10272 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_21_72
timestamp 1621261055
transform 1 0 8064 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_80
timestamp 1621261055
transform 1 0 8832 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_88
timestamp 1621261055
transform 1 0 9600 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_92
timestamp 1621261055
transform 1 0 9984 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_94
timestamp 1621261055
transform 1 0 10176 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_98
timestamp 1621261055
transform 1 0 10560 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_396
timestamp 1621261055
transform 1 0 11712 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_106
timestamp 1621261055
transform 1 0 11328 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_111
timestamp 1621261055
transform 1 0 11808 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_119
timestamp 1621261055
transform 1 0 12576 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_127
timestamp 1621261055
transform 1 0 13344 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_397
timestamp 1621261055
transform 1 0 16992 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_135
timestamp 1621261055
transform 1 0 14112 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_143
timestamp 1621261055
transform 1 0 14880 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_151
timestamp 1621261055
transform 1 0 15648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_159
timestamp 1621261055
transform 1 0 16416 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_163
timestamp 1621261055
transform 1 0 16800 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_166
timestamp 1621261055
transform 1 0 17088 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_174
timestamp 1621261055
transform 1 0 17856 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_182
timestamp 1621261055
transform 1 0 18624 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_190
timestamp 1621261055
transform 1 0 19392 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_198
timestamp 1621261055
transform 1 0 20160 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_398
timestamp 1621261055
transform 1 0 22272 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_206
timestamp 1621261055
transform 1 0 20928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_214
timestamp 1621261055
transform 1 0 21696 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_218
timestamp 1621261055
transform 1 0 22080 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_221
timestamp 1621261055
transform 1 0 22368 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_229
timestamp 1621261055
transform 1 0 23136 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_237
timestamp 1621261055
transform 1 0 23904 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_245
timestamp 1621261055
transform 1 0 24672 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_253
timestamp 1621261055
transform 1 0 25440 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_261
timestamp 1621261055
transform 1 0 26208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_399
timestamp 1621261055
transform 1 0 27552 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_269
timestamp 1621261055
transform 1 0 26976 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_273
timestamp 1621261055
transform 1 0 27360 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_276
timestamp 1621261055
transform 1 0 27648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_284
timestamp 1621261055
transform 1 0 28416 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_292
timestamp 1621261055
transform 1 0 29184 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_400
timestamp 1621261055
transform 1 0 32832 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_300
timestamp 1621261055
transform 1 0 29952 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_308
timestamp 1621261055
transform 1 0 30720 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_316
timestamp 1621261055
transform 1 0 31488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_324
timestamp 1621261055
transform 1 0 32256 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_328
timestamp 1621261055
transform 1 0 32640 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _067_
timestamp 1621261055
transform 1 0 35328 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_21_331
timestamp 1621261055
transform 1 0 32928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_339
timestamp 1621261055
transform 1 0 33696 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_347
timestamp 1621261055
transform 1 0 34464 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_21_355
timestamp 1621261055
transform 1 0 35232 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_359
timestamp 1621261055
transform 1 0 35616 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_401
timestamp 1621261055
transform 1 0 38112 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_367
timestamp 1621261055
transform 1 0 36384 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_375
timestamp 1621261055
transform 1 0 37152 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_383
timestamp 1621261055
transform 1 0 37920 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_386
timestamp 1621261055
transform 1 0 38208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_394
timestamp 1621261055
transform 1 0 38976 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_402
timestamp 1621261055
transform 1 0 39744 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_410
timestamp 1621261055
transform 1 0 40512 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_418
timestamp 1621261055
transform 1 0 41280 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_426
timestamp 1621261055
transform 1 0 42048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_402
timestamp 1621261055
transform 1 0 43392 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_434
timestamp 1621261055
transform 1 0 42816 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_438
timestamp 1621261055
transform 1 0 43200 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_441
timestamp 1621261055
transform 1 0 43488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_449
timestamp 1621261055
transform 1 0 44256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_457
timestamp 1621261055
transform 1 0 45024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _095_
timestamp 1621261055
transform 1 0 45888 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_403
timestamp 1621261055
transform 1 0 48672 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_21_465
timestamp 1621261055
transform 1 0 45792 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_469
timestamp 1621261055
transform 1 0 46176 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_477
timestamp 1621261055
transform 1 0 46944 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_485
timestamp 1621261055
transform 1 0 47712 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_493
timestamp 1621261055
transform 1 0 48480 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_496
timestamp 1621261055
transform 1 0 48768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_504
timestamp 1621261055
transform 1 0 49536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_512
timestamp 1621261055
transform 1 0 50304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_520
timestamp 1621261055
transform 1 0 51072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_528
timestamp 1621261055
transform 1 0 51840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _107_
timestamp 1621261055
transform 1 0 54432 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_404
timestamp 1621261055
transform 1 0 53952 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_536
timestamp 1621261055
transform 1 0 52608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_544
timestamp 1621261055
transform 1 0 53376 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_548
timestamp 1621261055
transform 1 0 53760 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_21_551
timestamp 1621261055
transform 1 0 54048 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_558
timestamp 1621261055
transform 1 0 54720 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_566
timestamp 1621261055
transform 1 0 55488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_574
timestamp 1621261055
transform 1 0 56256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_582
timestamp 1621261055
transform 1 0 57024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_590
timestamp 1621261055
transform 1 0 57792 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_594
timestamp 1621261055
transform 1 0 58176 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_43
timestamp 1621261055
transform -1 0 58848 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_21_596
timestamp 1621261055
transform 1 0 58368 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_44
timestamp 1621261055
transform 1 0 1152 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_405
timestamp 1621261055
transform 1 0 3840 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_4
timestamp 1621261055
transform 1 0 1536 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_12
timestamp 1621261055
transform 1 0 2304 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_20
timestamp 1621261055
transform 1 0 3072 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_29
timestamp 1621261055
transform 1 0 3936 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_37
timestamp 1621261055
transform 1 0 4704 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_45
timestamp 1621261055
transform 1 0 5472 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_53
timestamp 1621261055
transform 1 0 6240 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_61
timestamp 1621261055
transform 1 0 7008 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_406
timestamp 1621261055
transform 1 0 9120 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_69
timestamp 1621261055
transform 1 0 7776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_77
timestamp 1621261055
transform 1 0 8544 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_81
timestamp 1621261055
transform 1 0 8928 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_84
timestamp 1621261055
transform 1 0 9216 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_92
timestamp 1621261055
transform 1 0 9984 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_100
timestamp 1621261055
transform 1 0 10752 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_108
timestamp 1621261055
transform 1 0 11520 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_116
timestamp 1621261055
transform 1 0 12288 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_124
timestamp 1621261055
transform 1 0 13056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_132
timestamp 1621261055
transform 1 0 13824 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_407
timestamp 1621261055
transform 1 0 14400 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_136
timestamp 1621261055
transform 1 0 14208 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_139
timestamp 1621261055
transform 1 0 14496 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_147
timestamp 1621261055
transform 1 0 15264 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_155
timestamp 1621261055
transform 1 0 16032 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_163
timestamp 1621261055
transform 1 0 16800 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_408
timestamp 1621261055
transform 1 0 19680 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_171
timestamp 1621261055
transform 1 0 17568 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_179
timestamp 1621261055
transform 1 0 18336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_187
timestamp 1621261055
transform 1 0 19104 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_191
timestamp 1621261055
transform 1 0 19488 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_194
timestamp 1621261055
transform 1 0 19776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _191_
timestamp 1621261055
transform 1 0 22944 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_22_202
timestamp 1621261055
transform 1 0 20544 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_210
timestamp 1621261055
transform 1 0 21312 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_218
timestamp 1621261055
transform 1 0 22080 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_22_226
timestamp 1621261055
transform 1 0 22848 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_230
timestamp 1621261055
transform 1 0 23232 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_409
timestamp 1621261055
transform 1 0 24960 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_238
timestamp 1621261055
transform 1 0 24000 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_246
timestamp 1621261055
transform 1 0 24768 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_249
timestamp 1621261055
transform 1 0 25056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_257
timestamp 1621261055
transform 1 0 25824 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _020_
timestamp 1621261055
transform 1 0 27264 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_30
timestamp 1621261055
transform 1 0 27072 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_22_265
timestamp 1621261055
transform 1 0 26592 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_22_269
timestamp 1621261055
transform 1 0 26976 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_275
timestamp 1621261055
transform 1 0 27552 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_283
timestamp 1621261055
transform 1 0 28320 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_291
timestamp 1621261055
transform 1 0 29088 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_410
timestamp 1621261055
transform 1 0 30240 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_299
timestamp 1621261055
transform 1 0 29856 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_22_304
timestamp 1621261055
transform 1 0 30336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_312
timestamp 1621261055
transform 1 0 31104 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_320
timestamp 1621261055
transform 1 0 31872 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_328
timestamp 1621261055
transform 1 0 32640 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_411
timestamp 1621261055
transform 1 0 35520 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_336
timestamp 1621261055
transform 1 0 33408 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_344
timestamp 1621261055
transform 1 0 34176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_352
timestamp 1621261055
transform 1 0 34944 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_356
timestamp 1621261055
transform 1 0 35328 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_359
timestamp 1621261055
transform 1 0 35616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_367
timestamp 1621261055
transform 1 0 36384 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_375
timestamp 1621261055
transform 1 0 37152 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_383
timestamp 1621261055
transform 1 0 37920 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_391
timestamp 1621261055
transform 1 0 38688 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_412
timestamp 1621261055
transform 1 0 40800 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_399
timestamp 1621261055
transform 1 0 39456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_407
timestamp 1621261055
transform 1 0 40224 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_411
timestamp 1621261055
transform 1 0 40608 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_414
timestamp 1621261055
transform 1 0 40896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_422
timestamp 1621261055
transform 1 0 41664 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_430
timestamp 1621261055
transform 1 0 42432 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_438
timestamp 1621261055
transform 1 0 43200 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_446
timestamp 1621261055
transform 1 0 43968 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_454
timestamp 1621261055
transform 1 0 44736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_462
timestamp 1621261055
transform 1 0 45504 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _126_
timestamp 1621261055
transform 1 0 46560 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_413
timestamp 1621261055
transform 1 0 46080 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_466
timestamp 1621261055
transform 1 0 45888 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_22_469
timestamp 1621261055
transform 1 0 46176 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_22_476
timestamp 1621261055
transform 1 0 46848 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_484
timestamp 1621261055
transform 1 0 47616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_492
timestamp 1621261055
transform 1 0 48384 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_414
timestamp 1621261055
transform 1 0 51360 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_500
timestamp 1621261055
transform 1 0 49152 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_508
timestamp 1621261055
transform 1 0 49920 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_516
timestamp 1621261055
transform 1 0 50688 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_520
timestamp 1621261055
transform 1 0 51072 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_22_522
timestamp 1621261055
transform 1 0 51264 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_524
timestamp 1621261055
transform 1 0 51456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _082_
timestamp 1621261055
transform 1 0 53856 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_22_532
timestamp 1621261055
transform 1 0 52224 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_540
timestamp 1621261055
transform 1 0 52992 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_22_548
timestamp 1621261055
transform 1 0 53760 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_552
timestamp 1621261055
transform 1 0 54144 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_560
timestamp 1621261055
transform 1 0 54912 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_415
timestamp 1621261055
transform 1 0 56640 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_568
timestamp 1621261055
transform 1 0 55680 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_576
timestamp 1621261055
transform 1 0 56448 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_579
timestamp 1621261055
transform 1 0 56736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_587
timestamp 1621261055
transform 1 0 57504 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_45
timestamp 1621261055
transform -1 0 58848 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_595
timestamp 1621261055
transform 1 0 58272 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_4
timestamp 1621261055
transform 1 0 1536 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_4
timestamp 1621261055
transform 1 0 1536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_48
timestamp 1621261055
transform 1 0 1152 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_46
timestamp 1621261055
transform 1 0 1152 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_12
timestamp 1621261055
transform 1 0 2304 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_12
timestamp 1621261055
transform 1 0 2304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_20
timestamp 1621261055
transform 1 0 3072 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_20
timestamp 1621261055
transform 1 0 3072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_29
timestamp 1621261055
transform 1 0 3936 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_28
timestamp 1621261055
transform 1 0 3840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_426
timestamp 1621261055
transform 1 0 3840 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_24_43
timestamp 1621261055
transform 1 0 5280 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_41
timestamp 1621261055
transform 1 0 5088 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_37
timestamp 1621261055
transform 1 0 4704 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_44
timestamp 1621261055
transform 1 0 5376 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_36
timestamp 1621261055
transform 1 0 4608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_38
timestamp 1621261055
transform 1 0 5376 0 -1 19314
box -38 -49 230 715
use AOI22X1  AOI22X1
timestamp 1623610208
transform 1 0 5568 0 -1 19314
box 0 -48 1440 714
use sky130_fd_sc_ls__decap_8  FILLER_24_61
timestamp 1621261055
transform 1 0 7008 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_56
timestamp 1621261055
transform 1 0 6528 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_54
timestamp 1621261055
transform 1 0 6336 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_52
timestamp 1621261055
transform 1 0 6144 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_416
timestamp 1621261055
transform 1 0 6432 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_64
timestamp 1621261055
transform 1 0 7296 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_69
timestamp 1621261055
transform 1 0 7776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_72
timestamp 1621261055
transform 1 0 8064 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_81
timestamp 1621261055
transform 1 0 8928 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_77
timestamp 1621261055
transform 1 0 8544 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_80
timestamp 1621261055
transform 1 0 8832 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_427
timestamp 1621261055
transform 1 0 9120 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_92
timestamp 1621261055
transform 1 0 9984 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_84
timestamp 1621261055
transform 1 0 9216 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_88
timestamp 1621261055
transform 1 0 9600 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_96
timestamp 1621261055
transform 1 0 10368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_100
timestamp 1621261055
transform 1 0 10752 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_104
timestamp 1621261055
transform 1 0 11136 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_116
timestamp 1621261055
transform 1 0 12288 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_108
timestamp 1621261055
transform 1 0 11520 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_111
timestamp 1621261055
transform 1 0 11808 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_108
timestamp 1621261055
transform 1 0 11520 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_417
timestamp 1621261055
transform 1 0 11712 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_124
timestamp 1621261055
transform 1 0 13056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_119
timestamp 1621261055
transform 1 0 12576 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_132
timestamp 1621261055
transform 1 0 13824 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_127
timestamp 1621261055
transform 1 0 13344 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_139
timestamp 1621261055
transform 1 0 14496 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_136
timestamp 1621261055
transform 1 0 14208 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_135
timestamp 1621261055
transform 1 0 14112 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_428
timestamp 1621261055
transform 1 0 14400 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_147
timestamp 1621261055
transform 1 0 15264 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_143
timestamp 1621261055
transform 1 0 14880 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_155
timestamp 1621261055
transform 1 0 16032 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_151
timestamp 1621261055
transform 1 0 15648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_163
timestamp 1621261055
transform 1 0 16800 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_163
timestamp 1621261055
transform 1 0 16800 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_159
timestamp 1621261055
transform 1 0 16416 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_418
timestamp 1621261055
transform 1 0 16992 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_171
timestamp 1621261055
transform 1 0 17568 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_166
timestamp 1621261055
transform 1 0 17088 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_179
timestamp 1621261055
transform 1 0 18336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_182
timestamp 1621261055
transform 1 0 18624 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_174
timestamp 1621261055
transform 1 0 17856 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_191
timestamp 1621261055
transform 1 0 19488 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_187
timestamp 1621261055
transform 1 0 19104 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_190
timestamp 1621261055
transform 1 0 19392 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_194
timestamp 1621261055
transform 1 0 19776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_198
timestamp 1621261055
transform 1 0 20160 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_429
timestamp 1621261055
transform 1 0 19680 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_202
timestamp 1621261055
transform 1 0 20544 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_206
timestamp 1621261055
transform 1 0 20928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_210
timestamp 1621261055
transform 1 0 21312 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_214
timestamp 1621261055
transform 1 0 21696 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_218
timestamp 1621261055
transform 1 0 22080 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_221
timestamp 1621261055
transform 1 0 22368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_218
timestamp 1621261055
transform 1 0 22080 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_419
timestamp 1621261055
transform 1 0 22272 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_226
timestamp 1621261055
transform 1 0 22848 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_229
timestamp 1621261055
transform 1 0 23136 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_234
timestamp 1621261055
transform 1 0 23616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_237
timestamp 1621261055
transform 1 0 23904 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_246
timestamp 1621261055
transform 1 0 24768 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_242
timestamp 1621261055
transform 1 0 24384 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_245
timestamp 1621261055
transform 1 0 24672 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_430
timestamp 1621261055
transform 1 0 24960 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_257
timestamp 1621261055
transform 1 0 25824 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_249
timestamp 1621261055
transform 1 0 25056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_253
timestamp 1621261055
transform 1 0 25440 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_261
timestamp 1621261055
transform 1 0 26208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_265
timestamp 1621261055
transform 1 0 26592 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_269
timestamp 1621261055
transform 1 0 26976 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_281
timestamp 1621261055
transform 1 0 28128 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_273
timestamp 1621261055
transform 1 0 27360 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_276
timestamp 1621261055
transform 1 0 27648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_273
timestamp 1621261055
transform 1 0 27360 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_420
timestamp 1621261055
transform 1 0 27552 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_289
timestamp 1621261055
transform 1 0 28896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_284
timestamp 1621261055
transform 1 0 28416 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_297
timestamp 1621261055
transform 1 0 29664 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_292
timestamp 1621261055
transform 1 0 29184 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_304
timestamp 1621261055
transform 1 0 30336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_301
timestamp 1621261055
transform 1 0 30048 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_300
timestamp 1621261055
transform 1 0 29952 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_431
timestamp 1621261055
transform 1 0 30240 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_312
timestamp 1621261055
transform 1 0 31104 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_308
timestamp 1621261055
transform 1 0 30720 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_320
timestamp 1621261055
transform 1 0 31872 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_316
timestamp 1621261055
transform 1 0 31488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_328
timestamp 1621261055
transform 1 0 32640 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_328
timestamp 1621261055
transform 1 0 32640 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_324
timestamp 1621261055
transform 1 0 32256 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_421
timestamp 1621261055
transform 1 0 32832 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_336
timestamp 1621261055
transform 1 0 33408 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_331
timestamp 1621261055
transform 1 0 32928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_344
timestamp 1621261055
transform 1 0 34176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_343
timestamp 1621261055
transform 1 0 34080 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_339
timestamp 1621261055
transform 1 0 33696 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _205_
timestamp 1621261055
transform 1 0 33792 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_356
timestamp 1621261055
transform 1 0 35328 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_352
timestamp 1621261055
transform 1 0 34944 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_351
timestamp 1621261055
transform 1 0 34848 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_359
timestamp 1621261055
transform 1 0 35616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_359
timestamp 1621261055
transform 1 0 35616 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_432
timestamp 1621261055
transform 1 0 35520 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_367
timestamp 1621261055
transform 1 0 36384 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_367
timestamp 1621261055
transform 1 0 36384 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_375
timestamp 1621261055
transform 1 0 37152 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_375
timestamp 1621261055
transform 1 0 37152 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_383
timestamp 1621261055
transform 1 0 37920 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_386
timestamp 1621261055
transform 1 0 38208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_383
timestamp 1621261055
transform 1 0 37920 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_422
timestamp 1621261055
transform 1 0 38112 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_391
timestamp 1621261055
transform 1 0 38688 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_394
timestamp 1621261055
transform 1 0 38976 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_399
timestamp 1621261055
transform 1 0 39456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_402
timestamp 1621261055
transform 1 0 39744 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_411
timestamp 1621261055
transform 1 0 40608 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_407
timestamp 1621261055
transform 1 0 40224 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_410
timestamp 1621261055
transform 1 0 40512 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_433
timestamp 1621261055
transform 1 0 40800 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_422
timestamp 1621261055
transform 1 0 41664 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_414
timestamp 1621261055
transform 1 0 40896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_418
timestamp 1621261055
transform 1 0 41280 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_426
timestamp 1621261055
transform 1 0 42048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_430
timestamp 1621261055
transform 1 0 42432 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_434
timestamp 1621261055
transform 1 0 42816 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_446
timestamp 1621261055
transform 1 0 43968 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_438
timestamp 1621261055
transform 1 0 43200 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_441
timestamp 1621261055
transform 1 0 43488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_438
timestamp 1621261055
transform 1 0 43200 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_423
timestamp 1621261055
transform 1 0 43392 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_454
timestamp 1621261055
transform 1 0 44736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_449
timestamp 1621261055
transform 1 0 44256 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_462
timestamp 1621261055
transform 1 0 45504 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_457
timestamp 1621261055
transform 1 0 45024 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_469
timestamp 1621261055
transform 1 0 46176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_466
timestamp 1621261055
transform 1 0 45888 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_465
timestamp 1621261055
transform 1 0 45792 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_434
timestamp 1621261055
transform 1 0 46080 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_477
timestamp 1621261055
transform 1 0 46944 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_473
timestamp 1621261055
transform 1 0 46560 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_485
timestamp 1621261055
transform 1 0 47712 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_481
timestamp 1621261055
transform 1 0 47328 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_493
timestamp 1621261055
transform 1 0 48480 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_493
timestamp 1621261055
transform 1 0 48480 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_489
timestamp 1621261055
transform 1 0 48096 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_424
timestamp 1621261055
transform 1 0 48672 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_501
timestamp 1621261055
transform 1 0 49248 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_496
timestamp 1621261055
transform 1 0 48768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_509
timestamp 1621261055
transform 1 0 50016 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_512
timestamp 1621261055
transform 1 0 50304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_504
timestamp 1621261055
transform 1 0 49536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_521
timestamp 1621261055
transform 1 0 51168 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_517
timestamp 1621261055
transform 1 0 50784 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_520
timestamp 1621261055
transform 1 0 51072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_524
timestamp 1621261055
transform 1 0 51456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_528
timestamp 1621261055
transform 1 0 51840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_435
timestamp 1621261055
transform 1 0 51360 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_532
timestamp 1621261055
transform 1 0 52224 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_536
timestamp 1621261055
transform 1 0 52608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_540
timestamp 1621261055
transform 1 0 52992 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_544
timestamp 1621261055
transform 1 0 53376 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_548
timestamp 1621261055
transform 1 0 53760 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_551
timestamp 1621261055
transform 1 0 54048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_548
timestamp 1621261055
transform 1 0 53760 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_425
timestamp 1621261055
transform 1 0 53952 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_556
timestamp 1621261055
transform 1 0 54528 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_559
timestamp 1621261055
transform 1 0 54816 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_564
timestamp 1621261055
transform 1 0 55296 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_567
timestamp 1621261055
transform 1 0 55584 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_576
timestamp 1621261055
transform 1 0 56448 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_572
timestamp 1621261055
transform 1 0 56064 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_575
timestamp 1621261055
transform 1 0 56352 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_436
timestamp 1621261055
transform 1 0 56640 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_587
timestamp 1621261055
transform 1 0 57504 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_579
timestamp 1621261055
transform 1 0 56736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_583
timestamp 1621261055
transform 1 0 57120 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_591
timestamp 1621261055
transform 1 0 57888 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_47
timestamp 1621261055
transform -1 0 58848 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_49
timestamp 1621261055
transform -1 0 58848 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_595
timestamp 1621261055
transform 1 0 58272 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_595
timestamp 1621261055
transform 1 0 58272 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _078_
timestamp 1621261055
transform 1 0 1536 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_50
timestamp 1621261055
transform 1 0 1152 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_7
timestamp 1621261055
transform 1 0 1824 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_15
timestamp 1621261055
transform 1 0 2592 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_23
timestamp 1621261055
transform 1 0 3360 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_31
timestamp 1621261055
transform 1 0 4128 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_437
timestamp 1621261055
transform 1 0 6432 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_39
timestamp 1621261055
transform 1 0 4896 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_47
timestamp 1621261055
transform 1 0 5664 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_56
timestamp 1621261055
transform 1 0 6528 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_64
timestamp 1621261055
transform 1 0 7296 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _117_
timestamp 1621261055
transform 1 0 8256 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_72
timestamp 1621261055
transform 1 0 8064 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_77
timestamp 1621261055
transform 1 0 8544 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_85
timestamp 1621261055
transform 1 0 9312 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_93
timestamp 1621261055
transform 1 0 10080 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _140_
timestamp 1621261055
transform 1 0 13728 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_438
timestamp 1621261055
transform 1 0 11712 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_101
timestamp 1621261055
transform 1 0 10848 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_25_109
timestamp 1621261055
transform 1 0 11616 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_111
timestamp 1621261055
transform 1 0 11808 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_119
timestamp 1621261055
transform 1 0 12576 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_127
timestamp 1621261055
transform 1 0 13344 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_439
timestamp 1621261055
transform 1 0 16992 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_134
timestamp 1621261055
transform 1 0 14016 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_142
timestamp 1621261055
transform 1 0 14784 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_150
timestamp 1621261055
transform 1 0 15552 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_158
timestamp 1621261055
transform 1 0 16320 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_162
timestamp 1621261055
transform 1 0 16704 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_164
timestamp 1621261055
transform 1 0 16896 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_166
timestamp 1621261055
transform 1 0 17088 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_174
timestamp 1621261055
transform 1 0 17856 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_182
timestamp 1621261055
transform 1 0 18624 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_190
timestamp 1621261055
transform 1 0 19392 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_198
timestamp 1621261055
transform 1 0 20160 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_440
timestamp 1621261055
transform 1 0 22272 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_206
timestamp 1621261055
transform 1 0 20928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_214
timestamp 1621261055
transform 1 0 21696 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_218
timestamp 1621261055
transform 1 0 22080 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_221
timestamp 1621261055
transform 1 0 22368 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_229
timestamp 1621261055
transform 1 0 23136 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_237
timestamp 1621261055
transform 1 0 23904 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_245
timestamp 1621261055
transform 1 0 24672 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_253
timestamp 1621261055
transform 1 0 25440 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_261
timestamp 1621261055
transform 1 0 26208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _202_
timestamp 1621261055
transform 1 0 28032 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_441
timestamp 1621261055
transform 1 0 27552 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_269
timestamp 1621261055
transform 1 0 26976 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_273
timestamp 1621261055
transform 1 0 27360 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_25_276
timestamp 1621261055
transform 1 0 27648 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_283
timestamp 1621261055
transform 1 0 28320 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_291
timestamp 1621261055
transform 1 0 29088 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_442
timestamp 1621261055
transform 1 0 32832 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_299
timestamp 1621261055
transform 1 0 29856 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_307
timestamp 1621261055
transform 1 0 30624 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_315
timestamp 1621261055
transform 1 0 31392 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_323
timestamp 1621261055
transform 1 0 32160 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_327
timestamp 1621261055
transform 1 0 32544 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_329
timestamp 1621261055
transform 1 0 32736 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_331
timestamp 1621261055
transform 1 0 32928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_339
timestamp 1621261055
transform 1 0 33696 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_347
timestamp 1621261055
transform 1 0 34464 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_355
timestamp 1621261055
transform 1 0 35232 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_363
timestamp 1621261055
transform 1 0 36000 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _084_
timestamp 1621261055
transform 1 0 38688 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_443
timestamp 1621261055
transform 1 0 38112 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_371
timestamp 1621261055
transform 1 0 36768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_379
timestamp 1621261055
transform 1 0 37536 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_383
timestamp 1621261055
transform 1 0 37920 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_25_386
timestamp 1621261055
transform 1 0 38208 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_25_390
timestamp 1621261055
transform 1 0 38592 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_394
timestamp 1621261055
transform 1 0 38976 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_402
timestamp 1621261055
transform 1 0 39744 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_410
timestamp 1621261055
transform 1 0 40512 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_418
timestamp 1621261055
transform 1 0 41280 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_426
timestamp 1621261055
transform 1 0 42048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_444
timestamp 1621261055
transform 1 0 43392 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_434
timestamp 1621261055
transform 1 0 42816 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_438
timestamp 1621261055
transform 1 0 43200 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_441
timestamp 1621261055
transform 1 0 43488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_449
timestamp 1621261055
transform 1 0 44256 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_457
timestamp 1621261055
transform 1 0 45024 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_445
timestamp 1621261055
transform 1 0 48672 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_465
timestamp 1621261055
transform 1 0 45792 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_473
timestamp 1621261055
transform 1 0 46560 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_481
timestamp 1621261055
transform 1 0 47328 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_489
timestamp 1621261055
transform 1 0 48096 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_493
timestamp 1621261055
transform 1 0 48480 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_496
timestamp 1621261055
transform 1 0 48768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_504
timestamp 1621261055
transform 1 0 49536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_512
timestamp 1621261055
transform 1 0 50304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_520
timestamp 1621261055
transform 1 0 51072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_528
timestamp 1621261055
transform 1 0 51840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_446
timestamp 1621261055
transform 1 0 53952 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_536
timestamp 1621261055
transform 1 0 52608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_544
timestamp 1621261055
transform 1 0 53376 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_548
timestamp 1621261055
transform 1 0 53760 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_551
timestamp 1621261055
transform 1 0 54048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_559
timestamp 1621261055
transform 1 0 54816 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_567
timestamp 1621261055
transform 1 0 55584 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_575
timestamp 1621261055
transform 1 0 56352 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_583
timestamp 1621261055
transform 1 0 57120 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_591
timestamp 1621261055
transform 1 0 57888 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_51
timestamp 1621261055
transform -1 0 58848 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_595
timestamp 1621261055
transform 1 0 58272 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_52
timestamp 1621261055
transform 1 0 1152 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_447
timestamp 1621261055
transform 1 0 3840 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_4
timestamp 1621261055
transform 1 0 1536 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_12
timestamp 1621261055
transform 1 0 2304 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_20
timestamp 1621261055
transform 1 0 3072 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_29
timestamp 1621261055
transform 1 0 3936 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_37
timestamp 1621261055
transform 1 0 4704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_45
timestamp 1621261055
transform 1 0 5472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_53
timestamp 1621261055
transform 1 0 6240 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_61
timestamp 1621261055
transform 1 0 7008 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_448
timestamp 1621261055
transform 1 0 9120 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_69
timestamp 1621261055
transform 1 0 7776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_77
timestamp 1621261055
transform 1 0 8544 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_81
timestamp 1621261055
transform 1 0 8928 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_84
timestamp 1621261055
transform 1 0 9216 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_92
timestamp 1621261055
transform 1 0 9984 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_100
timestamp 1621261055
transform 1 0 10752 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_108
timestamp 1621261055
transform 1 0 11520 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_116
timestamp 1621261055
transform 1 0 12288 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_124
timestamp 1621261055
transform 1 0 13056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_132
timestamp 1621261055
transform 1 0 13824 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_449
timestamp 1621261055
transform 1 0 14400 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_136
timestamp 1621261055
transform 1 0 14208 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_139
timestamp 1621261055
transform 1 0 14496 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_147
timestamp 1621261055
transform 1 0 15264 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_155
timestamp 1621261055
transform 1 0 16032 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_163
timestamp 1621261055
transform 1 0 16800 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_450
timestamp 1621261055
transform 1 0 19680 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_171
timestamp 1621261055
transform 1 0 17568 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_179
timestamp 1621261055
transform 1 0 18336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_187
timestamp 1621261055
transform 1 0 19104 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_191
timestamp 1621261055
transform 1 0 19488 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_194
timestamp 1621261055
transform 1 0 19776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_202
timestamp 1621261055
transform 1 0 20544 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_210
timestamp 1621261055
transform 1 0 21312 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_218
timestamp 1621261055
transform 1 0 22080 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_226
timestamp 1621261055
transform 1 0 22848 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_451
timestamp 1621261055
transform 1 0 24960 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_234
timestamp 1621261055
transform 1 0 23616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_242
timestamp 1621261055
transform 1 0 24384 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_246
timestamp 1621261055
transform 1 0 24768 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_249
timestamp 1621261055
transform 1 0 25056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_257
timestamp 1621261055
transform 1 0 25824 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_265
timestamp 1621261055
transform 1 0 26592 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_273
timestamp 1621261055
transform 1 0 27360 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_281
timestamp 1621261055
transform 1 0 28128 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_289
timestamp 1621261055
transform 1 0 28896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_297
timestamp 1621261055
transform 1 0 29664 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_452
timestamp 1621261055
transform 1 0 30240 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_301
timestamp 1621261055
transform 1 0 30048 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_304
timestamp 1621261055
transform 1 0 30336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_312
timestamp 1621261055
transform 1 0 31104 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_320
timestamp 1621261055
transform 1 0 31872 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_328
timestamp 1621261055
transform 1 0 32640 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_453
timestamp 1621261055
transform 1 0 35520 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_336
timestamp 1621261055
transform 1 0 33408 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_344
timestamp 1621261055
transform 1 0 34176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_352
timestamp 1621261055
transform 1 0 34944 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_356
timestamp 1621261055
transform 1 0 35328 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_359
timestamp 1621261055
transform 1 0 35616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_367
timestamp 1621261055
transform 1 0 36384 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_375
timestamp 1621261055
transform 1 0 37152 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_383
timestamp 1621261055
transform 1 0 37920 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_391
timestamp 1621261055
transform 1 0 38688 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_454
timestamp 1621261055
transform 1 0 40800 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_399
timestamp 1621261055
transform 1 0 39456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_407
timestamp 1621261055
transform 1 0 40224 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_411
timestamp 1621261055
transform 1 0 40608 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_414
timestamp 1621261055
transform 1 0 40896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_422
timestamp 1621261055
transform 1 0 41664 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_430
timestamp 1621261055
transform 1 0 42432 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_438
timestamp 1621261055
transform 1 0 43200 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_446
timestamp 1621261055
transform 1 0 43968 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_454
timestamp 1621261055
transform 1 0 44736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_462
timestamp 1621261055
transform 1 0 45504 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_455
timestamp 1621261055
transform 1 0 46080 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_466
timestamp 1621261055
transform 1 0 45888 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_469
timestamp 1621261055
transform 1 0 46176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_477
timestamp 1621261055
transform 1 0 46944 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_485
timestamp 1621261055
transform 1 0 47712 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_493
timestamp 1621261055
transform 1 0 48480 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_456
timestamp 1621261055
transform 1 0 51360 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_501
timestamp 1621261055
transform 1 0 49248 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_509
timestamp 1621261055
transform 1 0 50016 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_517
timestamp 1621261055
transform 1 0 50784 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_521
timestamp 1621261055
transform 1 0 51168 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_524
timestamp 1621261055
transform 1 0 51456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_532
timestamp 1621261055
transform 1 0 52224 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_540
timestamp 1621261055
transform 1 0 52992 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_548
timestamp 1621261055
transform 1 0 53760 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_556
timestamp 1621261055
transform 1 0 54528 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_457
timestamp 1621261055
transform 1 0 56640 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_564
timestamp 1621261055
transform 1 0 55296 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_572
timestamp 1621261055
transform 1 0 56064 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_576
timestamp 1621261055
transform 1 0 56448 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_579
timestamp 1621261055
transform 1 0 56736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_587
timestamp 1621261055
transform 1 0 57504 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_53
timestamp 1621261055
transform -1 0 58848 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_595
timestamp 1621261055
transform 1 0 58272 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_54
timestamp 1621261055
transform 1 0 1152 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_4
timestamp 1621261055
transform 1 0 1536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_12
timestamp 1621261055
transform 1 0 2304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_20
timestamp 1621261055
transform 1 0 3072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_28
timestamp 1621261055
transform 1 0 3840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_458
timestamp 1621261055
transform 1 0 6432 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_36
timestamp 1621261055
transform 1 0 4608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_44
timestamp 1621261055
transform 1 0 5376 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_52
timestamp 1621261055
transform 1 0 6144 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_54
timestamp 1621261055
transform 1 0 6336 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_56
timestamp 1621261055
transform 1 0 6528 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_64
timestamp 1621261055
transform 1 0 7296 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_72
timestamp 1621261055
transform 1 0 8064 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_80
timestamp 1621261055
transform 1 0 8832 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_88
timestamp 1621261055
transform 1 0 9600 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_96
timestamp 1621261055
transform 1 0 10368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_459
timestamp 1621261055
transform 1 0 11712 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_104
timestamp 1621261055
transform 1 0 11136 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_108
timestamp 1621261055
transform 1 0 11520 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_111
timestamp 1621261055
transform 1 0 11808 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_119
timestamp 1621261055
transform 1 0 12576 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_127
timestamp 1621261055
transform 1 0 13344 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_460
timestamp 1621261055
transform 1 0 16992 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_135
timestamp 1621261055
transform 1 0 14112 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_143
timestamp 1621261055
transform 1 0 14880 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_151
timestamp 1621261055
transform 1 0 15648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_159
timestamp 1621261055
transform 1 0 16416 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_163
timestamp 1621261055
transform 1 0 16800 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_166
timestamp 1621261055
transform 1 0 17088 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_174
timestamp 1621261055
transform 1 0 17856 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_182
timestamp 1621261055
transform 1 0 18624 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_190
timestamp 1621261055
transform 1 0 19392 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_198
timestamp 1621261055
transform 1 0 20160 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_461
timestamp 1621261055
transform 1 0 22272 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_206
timestamp 1621261055
transform 1 0 20928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_214
timestamp 1621261055
transform 1 0 21696 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_218
timestamp 1621261055
transform 1 0 22080 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_221
timestamp 1621261055
transform 1 0 22368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_229
timestamp 1621261055
transform 1 0 23136 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_237
timestamp 1621261055
transform 1 0 23904 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_245
timestamp 1621261055
transform 1 0 24672 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_253
timestamp 1621261055
transform 1 0 25440 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_261
timestamp 1621261055
transform 1 0 26208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_462
timestamp 1621261055
transform 1 0 27552 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_269
timestamp 1621261055
transform 1 0 26976 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_273
timestamp 1621261055
transform 1 0 27360 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_276
timestamp 1621261055
transform 1 0 27648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_284
timestamp 1621261055
transform 1 0 28416 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_292
timestamp 1621261055
transform 1 0 29184 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_463
timestamp 1621261055
transform 1 0 32832 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_300
timestamp 1621261055
transform 1 0 29952 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_308
timestamp 1621261055
transform 1 0 30720 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_316
timestamp 1621261055
transform 1 0 31488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_324
timestamp 1621261055
transform 1 0 32256 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_328
timestamp 1621261055
transform 1 0 32640 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_331
timestamp 1621261055
transform 1 0 32928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_339
timestamp 1621261055
transform 1 0 33696 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_347
timestamp 1621261055
transform 1 0 34464 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_355
timestamp 1621261055
transform 1 0 35232 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_363
timestamp 1621261055
transform 1 0 36000 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _087_
timestamp 1621261055
transform 1 0 36864 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_464
timestamp 1621261055
transform 1 0 38112 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_27_371
timestamp 1621261055
transform 1 0 36768 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_375
timestamp 1621261055
transform 1 0 37152 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_383
timestamp 1621261055
transform 1 0 37920 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_386
timestamp 1621261055
transform 1 0 38208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_394
timestamp 1621261055
transform 1 0 38976 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_402
timestamp 1621261055
transform 1 0 39744 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_410
timestamp 1621261055
transform 1 0 40512 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_418
timestamp 1621261055
transform 1 0 41280 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_426
timestamp 1621261055
transform 1 0 42048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_465
timestamp 1621261055
transform 1 0 43392 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_434
timestamp 1621261055
transform 1 0 42816 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_438
timestamp 1621261055
transform 1 0 43200 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_441
timestamp 1621261055
transform 1 0 43488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_449
timestamp 1621261055
transform 1 0 44256 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_457
timestamp 1621261055
transform 1 0 45024 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _046_
timestamp 1621261055
transform -1 0 48000 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_466
timestamp 1621261055
transform 1 0 48672 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_40
timestamp 1621261055
transform -1 0 47712 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_465
timestamp 1621261055
transform 1 0 45792 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_473
timestamp 1621261055
transform 1 0 46560 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_481
timestamp 1621261055
transform 1 0 47328 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_27_488
timestamp 1621261055
transform 1 0 48000 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_492
timestamp 1621261055
transform 1 0 48384 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_494
timestamp 1621261055
transform 1 0 48576 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_496
timestamp 1621261055
transform 1 0 48768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_504
timestamp 1621261055
transform 1 0 49536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_512
timestamp 1621261055
transform 1 0 50304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_520
timestamp 1621261055
transform 1 0 51072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_528
timestamp 1621261055
transform 1 0 51840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_467
timestamp 1621261055
transform 1 0 53952 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_536
timestamp 1621261055
transform 1 0 52608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_544
timestamp 1621261055
transform 1 0 53376 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_548
timestamp 1621261055
transform 1 0 53760 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_551
timestamp 1621261055
transform 1 0 54048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_559
timestamp 1621261055
transform 1 0 54816 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_567
timestamp 1621261055
transform 1 0 55584 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_575
timestamp 1621261055
transform 1 0 56352 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_583
timestamp 1621261055
transform 1 0 57120 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_591
timestamp 1621261055
transform 1 0 57888 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_55
timestamp 1621261055
transform -1 0 58848 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_595
timestamp 1621261055
transform 1 0 58272 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_56
timestamp 1621261055
transform 1 0 1152 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_468
timestamp 1621261055
transform 1 0 3840 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_4
timestamp 1621261055
transform 1 0 1536 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_12
timestamp 1621261055
transform 1 0 2304 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_20
timestamp 1621261055
transform 1 0 3072 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_29
timestamp 1621261055
transform 1 0 3936 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _081_
timestamp 1621261055
transform 1 0 4896 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_37
timestamp 1621261055
transform 1 0 4704 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_42
timestamp 1621261055
transform 1 0 5184 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_50
timestamp 1621261055
transform 1 0 5952 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_58
timestamp 1621261055
transform 1 0 6720 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_66
timestamp 1621261055
transform 1 0 7488 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_469
timestamp 1621261055
transform 1 0 9120 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_74
timestamp 1621261055
transform 1 0 8256 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_28_82
timestamp 1621261055
transform 1 0 9024 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_84
timestamp 1621261055
transform 1 0 9216 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_92
timestamp 1621261055
transform 1 0 9984 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_100
timestamp 1621261055
transform 1 0 10752 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_108
timestamp 1621261055
transform 1 0 11520 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_116
timestamp 1621261055
transform 1 0 12288 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_124
timestamp 1621261055
transform 1 0 13056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_132
timestamp 1621261055
transform 1 0 13824 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _157_
timestamp 1621261055
transform 1 0 14880 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_470
timestamp 1621261055
transform 1 0 14400 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_136
timestamp 1621261055
transform 1 0 14208 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_28_139
timestamp 1621261055
transform 1 0 14496 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_28_146
timestamp 1621261055
transform 1 0 15168 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_154
timestamp 1621261055
transform 1 0 15936 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_162
timestamp 1621261055
transform 1 0 16704 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_471
timestamp 1621261055
transform 1 0 19680 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_170
timestamp 1621261055
transform 1 0 17472 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_178
timestamp 1621261055
transform 1 0 18240 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_186
timestamp 1621261055
transform 1 0 19008 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_190
timestamp 1621261055
transform 1 0 19392 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_28_192
timestamp 1621261055
transform 1 0 19584 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_194
timestamp 1621261055
transform 1 0 19776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_202
timestamp 1621261055
transform 1 0 20544 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_210
timestamp 1621261055
transform 1 0 21312 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_218
timestamp 1621261055
transform 1 0 22080 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_226
timestamp 1621261055
transform 1 0 22848 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_472
timestamp 1621261055
transform 1 0 24960 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_234
timestamp 1621261055
transform 1 0 23616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_242
timestamp 1621261055
transform 1 0 24384 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_246
timestamp 1621261055
transform 1 0 24768 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_249
timestamp 1621261055
transform 1 0 25056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_257
timestamp 1621261055
transform 1 0 25824 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_265
timestamp 1621261055
transform 1 0 26592 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_273
timestamp 1621261055
transform 1 0 27360 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_281
timestamp 1621261055
transform 1 0 28128 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_289
timestamp 1621261055
transform 1 0 28896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_297
timestamp 1621261055
transform 1 0 29664 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_473
timestamp 1621261055
transform 1 0 30240 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_301
timestamp 1621261055
transform 1 0 30048 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_304
timestamp 1621261055
transform 1 0 30336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_312
timestamp 1621261055
transform 1 0 31104 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_320
timestamp 1621261055
transform 1 0 31872 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_328
timestamp 1621261055
transform 1 0 32640 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_474
timestamp 1621261055
transform 1 0 35520 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_336
timestamp 1621261055
transform 1 0 33408 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_344
timestamp 1621261055
transform 1 0 34176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_352
timestamp 1621261055
transform 1 0 34944 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_356
timestamp 1621261055
transform 1 0 35328 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_359
timestamp 1621261055
transform 1 0 35616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_367
timestamp 1621261055
transform 1 0 36384 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_375
timestamp 1621261055
transform 1 0 37152 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_383
timestamp 1621261055
transform 1 0 37920 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_391
timestamp 1621261055
transform 1 0 38688 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_475
timestamp 1621261055
transform 1 0 40800 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_399
timestamp 1621261055
transform 1 0 39456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_407
timestamp 1621261055
transform 1 0 40224 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_411
timestamp 1621261055
transform 1 0 40608 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_414
timestamp 1621261055
transform 1 0 40896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_422
timestamp 1621261055
transform 1 0 41664 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_430
timestamp 1621261055
transform 1 0 42432 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_438
timestamp 1621261055
transform 1 0 43200 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_446
timestamp 1621261055
transform 1 0 43968 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_454
timestamp 1621261055
transform 1 0 44736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_462
timestamp 1621261055
transform 1 0 45504 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_476
timestamp 1621261055
transform 1 0 46080 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_466
timestamp 1621261055
transform 1 0 45888 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_469
timestamp 1621261055
transform 1 0 46176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_477
timestamp 1621261055
transform 1 0 46944 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_485
timestamp 1621261055
transform 1 0 47712 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_493
timestamp 1621261055
transform 1 0 48480 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_477
timestamp 1621261055
transform 1 0 51360 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_501
timestamp 1621261055
transform 1 0 49248 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_509
timestamp 1621261055
transform 1 0 50016 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_517
timestamp 1621261055
transform 1 0 50784 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_521
timestamp 1621261055
transform 1 0 51168 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_524
timestamp 1621261055
transform 1 0 51456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_532
timestamp 1621261055
transform 1 0 52224 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_540
timestamp 1621261055
transform 1 0 52992 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_548
timestamp 1621261055
transform 1 0 53760 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_556
timestamp 1621261055
transform 1 0 54528 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_478
timestamp 1621261055
transform 1 0 56640 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_564
timestamp 1621261055
transform 1 0 55296 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_572
timestamp 1621261055
transform 1 0 56064 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_576
timestamp 1621261055
transform 1 0 56448 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_579
timestamp 1621261055
transform 1 0 56736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_587
timestamp 1621261055
transform 1 0 57504 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_57
timestamp 1621261055
transform -1 0 58848 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_595
timestamp 1621261055
transform 1 0 58272 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_58
timestamp 1621261055
transform 1 0 1152 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_4
timestamp 1621261055
transform 1 0 1536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_12
timestamp 1621261055
transform 1 0 2304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_20
timestamp 1621261055
transform 1 0 3072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_28
timestamp 1621261055
transform 1 0 3840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_479
timestamp 1621261055
transform 1 0 6432 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_36
timestamp 1621261055
transform 1 0 4608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_44
timestamp 1621261055
transform 1 0 5376 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_52
timestamp 1621261055
transform 1 0 6144 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_54
timestamp 1621261055
transform 1 0 6336 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_56
timestamp 1621261055
transform 1 0 6528 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_64
timestamp 1621261055
transform 1 0 7296 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_72
timestamp 1621261055
transform 1 0 8064 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_80
timestamp 1621261055
transform 1 0 8832 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_88
timestamp 1621261055
transform 1 0 9600 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_96
timestamp 1621261055
transform 1 0 10368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_480
timestamp 1621261055
transform 1 0 11712 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_104
timestamp 1621261055
transform 1 0 11136 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_108
timestamp 1621261055
transform 1 0 11520 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_111
timestamp 1621261055
transform 1 0 11808 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_119
timestamp 1621261055
transform 1 0 12576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_127
timestamp 1621261055
transform 1 0 13344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _086_
timestamp 1621261055
transform 1 0 14880 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_481
timestamp 1621261055
transform 1 0 16992 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_135
timestamp 1621261055
transform 1 0 14112 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_146
timestamp 1621261055
transform 1 0 15168 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_154
timestamp 1621261055
transform 1 0 15936 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_162
timestamp 1621261055
transform 1 0 16704 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_164
timestamp 1621261055
transform 1 0 16896 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_166
timestamp 1621261055
transform 1 0 17088 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_174
timestamp 1621261055
transform 1 0 17856 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_182
timestamp 1621261055
transform 1 0 18624 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_190
timestamp 1621261055
transform 1 0 19392 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_198
timestamp 1621261055
transform 1 0 20160 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _146_
timestamp 1621261055
transform 1 0 20352 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_482
timestamp 1621261055
transform 1 0 22272 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_203
timestamp 1621261055
transform 1 0 20640 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_211
timestamp 1621261055
transform 1 0 21408 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_29_219
timestamp 1621261055
transform 1 0 22176 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_221
timestamp 1621261055
transform 1 0 22368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_229
timestamp 1621261055
transform 1 0 23136 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_237
timestamp 1621261055
transform 1 0 23904 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_245
timestamp 1621261055
transform 1 0 24672 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_253
timestamp 1621261055
transform 1 0 25440 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_261
timestamp 1621261055
transform 1 0 26208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_483
timestamp 1621261055
transform 1 0 27552 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_269
timestamp 1621261055
transform 1 0 26976 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_273
timestamp 1621261055
transform 1 0 27360 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_276
timestamp 1621261055
transform 1 0 27648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_284
timestamp 1621261055
transform 1 0 28416 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_292
timestamp 1621261055
transform 1 0 29184 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_484
timestamp 1621261055
transform 1 0 32832 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_300
timestamp 1621261055
transform 1 0 29952 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_308
timestamp 1621261055
transform 1 0 30720 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_316
timestamp 1621261055
transform 1 0 31488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_324
timestamp 1621261055
transform 1 0 32256 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_328
timestamp 1621261055
transform 1 0 32640 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _079_
timestamp 1621261055
transform 1 0 34752 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_29_331
timestamp 1621261055
transform 1 0 32928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_339
timestamp 1621261055
transform 1 0 33696 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_347
timestamp 1621261055
transform 1 0 34464 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_349
timestamp 1621261055
transform 1 0 34656 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_353
timestamp 1621261055
transform 1 0 35040 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_361
timestamp 1621261055
transform 1 0 35808 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_485
timestamp 1621261055
transform 1 0 38112 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_369
timestamp 1621261055
transform 1 0 36576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_377
timestamp 1621261055
transform 1 0 37344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_386
timestamp 1621261055
transform 1 0 38208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_394
timestamp 1621261055
transform 1 0 38976 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_402
timestamp 1621261055
transform 1 0 39744 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_410
timestamp 1621261055
transform 1 0 40512 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_418
timestamp 1621261055
transform 1 0 41280 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_426
timestamp 1621261055
transform 1 0 42048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_486
timestamp 1621261055
transform 1 0 43392 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_434
timestamp 1621261055
transform 1 0 42816 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_438
timestamp 1621261055
transform 1 0 43200 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_441
timestamp 1621261055
transform 1 0 43488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_449
timestamp 1621261055
transform 1 0 44256 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_457
timestamp 1621261055
transform 1 0 45024 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_487
timestamp 1621261055
transform 1 0 48672 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_465
timestamp 1621261055
transform 1 0 45792 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_473
timestamp 1621261055
transform 1 0 46560 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_481
timestamp 1621261055
transform 1 0 47328 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_489
timestamp 1621261055
transform 1 0 48096 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_493
timestamp 1621261055
transform 1 0 48480 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_496
timestamp 1621261055
transform 1 0 48768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_504
timestamp 1621261055
transform 1 0 49536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_512
timestamp 1621261055
transform 1 0 50304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_520
timestamp 1621261055
transform 1 0 51072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_528
timestamp 1621261055
transform 1 0 51840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_488
timestamp 1621261055
transform 1 0 53952 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_536
timestamp 1621261055
transform 1 0 52608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_544
timestamp 1621261055
transform 1 0 53376 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_548
timestamp 1621261055
transform 1 0 53760 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_551
timestamp 1621261055
transform 1 0 54048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_559
timestamp 1621261055
transform 1 0 54816 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_567
timestamp 1621261055
transform 1 0 55584 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_575
timestamp 1621261055
transform 1 0 56352 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_583
timestamp 1621261055
transform 1 0 57120 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_591
timestamp 1621261055
transform 1 0 57888 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_59
timestamp 1621261055
transform -1 0 58848 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_595
timestamp 1621261055
transform 1 0 58272 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_4
timestamp 1621261055
transform 1 0 1536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_4
timestamp 1621261055
transform 1 0 1536 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_62
timestamp 1621261055
transform 1 0 1152 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_60
timestamp 1621261055
transform 1 0 1152 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_12
timestamp 1621261055
transform 1 0 2304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_12
timestamp 1621261055
transform 1 0 2304 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_20
timestamp 1621261055
transform 1 0 3072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_20
timestamp 1621261055
transform 1 0 3072 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_28
timestamp 1621261055
transform 1 0 3840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_29
timestamp 1621261055
transform 1 0 3936 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_489
timestamp 1621261055
transform 1 0 3840 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_36
timestamp 1621261055
transform 1 0 4608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_37
timestamp 1621261055
transform 1 0 4704 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_44
timestamp 1621261055
transform 1 0 5376 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_45
timestamp 1621261055
transform 1 0 5472 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_56
timestamp 1621261055
transform 1 0 6528 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_54
timestamp 1621261055
transform 1 0 6336 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_52
timestamp 1621261055
transform 1 0 6144 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_53
timestamp 1621261055
transform 1 0 6240 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_500
timestamp 1621261055
transform 1 0 6432 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_64
timestamp 1621261055
transform 1 0 7296 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_61
timestamp 1621261055
transform 1 0 7008 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_74
timestamp 1621261055
transform 1 0 8256 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_72
timestamp 1621261055
transform 1 0 8064 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_73
timestamp 1621261055
transform 1 0 8160 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_69
timestamp 1621261055
transform 1 0 7776 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_78
timestamp 1621261055
transform 1 0 8640 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_79
timestamp 1621261055
transform 1 0 8736 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_30_75
timestamp 1621261055
transform 1 0 8352 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_490
timestamp 1621261055
transform 1 0 9120 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _193_
timestamp 1621261055
transform 1 0 8448 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _105_
timestamp 1621261055
transform 1 0 8352 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_86
timestamp 1621261055
transform 1 0 9408 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_92
timestamp 1621261055
transform 1 0 9984 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_84
timestamp 1621261055
transform 1 0 9216 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_94
timestamp 1621261055
transform 1 0 10176 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_102
timestamp 1621261055
transform 1 0 10944 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_100
timestamp 1621261055
transform 1 0 10752 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_111
timestamp 1621261055
transform 1 0 11808 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_116
timestamp 1621261055
transform 1 0 12288 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_108
timestamp 1621261055
transform 1 0 11520 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_501
timestamp 1621261055
transform 1 0 11712 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_119
timestamp 1621261055
transform 1 0 12576 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_124
timestamp 1621261055
transform 1 0 13056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_131
timestamp 1621261055
transform 1 0 13728 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_127
timestamp 1621261055
transform 1 0 13344 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_132
timestamp 1621261055
transform 1 0 13824 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _122_
timestamp 1621261055
transform 1 0 13440 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_139
timestamp 1621261055
transform 1 0 14496 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_139
timestamp 1621261055
transform 1 0 14496 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_136
timestamp 1621261055
transform 1 0 14208 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_491
timestamp 1621261055
transform 1 0 14400 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_147
timestamp 1621261055
transform 1 0 15264 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_147
timestamp 1621261055
transform 1 0 15264 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_155
timestamp 1621261055
transform 1 0 16032 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_155
timestamp 1621261055
transform 1 0 16032 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_163
timestamp 1621261055
transform 1 0 16800 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_163
timestamp 1621261055
transform 1 0 16800 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_502
timestamp 1621261055
transform 1 0 16992 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_166
timestamp 1621261055
transform 1 0 17088 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_171
timestamp 1621261055
transform 1 0 17568 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_182
timestamp 1621261055
transform 1 0 18624 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_174
timestamp 1621261055
transform 1 0 17856 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_179
timestamp 1621261055
transform 1 0 18336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_190
timestamp 1621261055
transform 1 0 19392 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_191
timestamp 1621261055
transform 1 0 19488 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_187
timestamp 1621261055
transform 1 0 19104 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_198
timestamp 1621261055
transform 1 0 20160 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_198
timestamp 1621261055
transform 1 0 20160 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_194
timestamp 1621261055
transform 1 0 19776 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_492
timestamp 1621261055
transform 1 0 19680 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_206
timestamp 1621261055
transform 1 0 20928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_205
timestamp 1621261055
transform 1 0 20832 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_25
timestamp 1621261055
transform -1 0 20544 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _014_
timestamp 1621261055
transform -1 0 20832 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_31_214
timestamp 1621261055
transform 1 0 21696 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_213
timestamp 1621261055
transform 1 0 21600 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_221
timestamp 1621261055
transform 1 0 22368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_218
timestamp 1621261055
transform 1 0 22080 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_221
timestamp 1621261055
transform 1 0 22368 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_503
timestamp 1621261055
transform 1 0 22272 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_229
timestamp 1621261055
transform 1 0 23136 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_229
timestamp 1621261055
transform 1 0 23136 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_237
timestamp 1621261055
transform 1 0 23904 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_239
timestamp 1621261055
transform 1 0 24096 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_235
timestamp 1621261055
transform 1 0 23712 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_233
timestamp 1621261055
transform 1 0 23520 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _068_
timestamp 1621261055
transform 1 0 23808 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_245
timestamp 1621261055
transform 1 0 24672 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_247
timestamp 1621261055
transform 1 0 24864 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_493
timestamp 1621261055
transform 1 0 24960 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_253
timestamp 1621261055
transform 1 0 25440 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_257
timestamp 1621261055
transform 1 0 25824 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_249
timestamp 1621261055
transform 1 0 25056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_261
timestamp 1621261055
transform 1 0 26208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_269
timestamp 1621261055
transform 1 0 26976 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_265
timestamp 1621261055
transform 1 0 26592 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_276
timestamp 1621261055
transform 1 0 27648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_273
timestamp 1621261055
transform 1 0 27360 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_281
timestamp 1621261055
transform 1 0 28128 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_273
timestamp 1621261055
transform 1 0 27360 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_504
timestamp 1621261055
transform 1 0 27552 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_284
timestamp 1621261055
transform 1 0 28416 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_289
timestamp 1621261055
transform 1 0 28896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_292
timestamp 1621261055
transform 1 0 29184 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_297
timestamp 1621261055
transform 1 0 29664 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_300
timestamp 1621261055
transform 1 0 29952 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_304
timestamp 1621261055
transform 1 0 30336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_301
timestamp 1621261055
transform 1 0 30048 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_494
timestamp 1621261055
transform 1 0 30240 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_308
timestamp 1621261055
transform 1 0 30720 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_312
timestamp 1621261055
transform 1 0 31104 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_316
timestamp 1621261055
transform 1 0 31488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_320
timestamp 1621261055
transform 1 0 31872 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_328
timestamp 1621261055
transform 1 0 32640 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_324
timestamp 1621261055
transform 1 0 32256 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_328
timestamp 1621261055
transform 1 0 32640 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_505
timestamp 1621261055
transform 1 0 32832 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_331
timestamp 1621261055
transform 1 0 32928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_336
timestamp 1621261055
transform 1 0 33408 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_347
timestamp 1621261055
transform 1 0 34464 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_339
timestamp 1621261055
transform 1 0 33696 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_344
timestamp 1621261055
transform 1 0 34176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_355
timestamp 1621261055
transform 1 0 35232 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_356
timestamp 1621261055
transform 1 0 35328 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_352
timestamp 1621261055
transform 1 0 34944 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_363
timestamp 1621261055
transform 1 0 36000 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_363
timestamp 1621261055
transform 1 0 36000 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_359
timestamp 1621261055
transform 1 0 35616 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_495
timestamp 1621261055
transform 1 0 35520 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_371
timestamp 1621261055
transform 1 0 36768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_367
timestamp 1621261055
transform 1 0 36384 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _188_
timestamp 1621261055
transform 1 0 36096 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_31_379
timestamp 1621261055
transform 1 0 37536 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_375
timestamp 1621261055
transform 1 0 37152 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_386
timestamp 1621261055
transform 1 0 38208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_383
timestamp 1621261055
transform 1 0 37920 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_383
timestamp 1621261055
transform 1 0 37920 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_506
timestamp 1621261055
transform 1 0 38112 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_394
timestamp 1621261055
transform 1 0 38976 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_391
timestamp 1621261055
transform 1 0 38688 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_402
timestamp 1621261055
transform 1 0 39744 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_399
timestamp 1621261055
transform 1 0 39456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_410
timestamp 1621261055
transform 1 0 40512 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_411
timestamp 1621261055
transform 1 0 40608 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_407
timestamp 1621261055
transform 1 0 40224 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_496
timestamp 1621261055
transform 1 0 40800 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_31_418
timestamp 1621261055
transform 1 0 41280 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_422
timestamp 1621261055
transform 1 0 41664 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_414
timestamp 1621261055
transform 1 0 40896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _090_
timestamp 1621261055
transform 1 0 41664 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_425
timestamp 1621261055
transform 1 0 41952 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_437
timestamp 1621261055
transform 1 0 43104 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_433
timestamp 1621261055
transform 1 0 42720 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_430
timestamp 1621261055
transform 1 0 42432 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_441
timestamp 1621261055
transform 1 0 43488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_439
timestamp 1621261055
transform 1 0 43296 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_446
timestamp 1621261055
transform 1 0 43968 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_438
timestamp 1621261055
transform 1 0 43200 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_507
timestamp 1621261055
transform 1 0 43392 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_449
timestamp 1621261055
transform 1 0 44256 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_454
timestamp 1621261055
transform 1 0 44736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_459
timestamp 1621261055
transform 1 0 45216 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_457
timestamp 1621261055
transform 1 0 45024 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_462
timestamp 1621261055
transform 1 0 45504 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _195_
timestamp 1621261055
transform 1 0 45312 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_463
timestamp 1621261055
transform 1 0 45600 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_469
timestamp 1621261055
transform 1 0 46176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_466
timestamp 1621261055
transform 1 0 45888 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_497
timestamp 1621261055
transform 1 0 46080 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_479
timestamp 1621261055
transform 1 0 47136 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_471
timestamp 1621261055
transform 1 0 46368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_477
timestamp 1621261055
transform 1 0 46944 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_487
timestamp 1621261055
transform 1 0 47904 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_485
timestamp 1621261055
transform 1 0 47712 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_493
timestamp 1621261055
transform 1 0 48480 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_508
timestamp 1621261055
transform 1 0 48672 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_496
timestamp 1621261055
transform 1 0 48768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_501
timestamp 1621261055
transform 1 0 49248 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_512
timestamp 1621261055
transform 1 0 50304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_504
timestamp 1621261055
transform 1 0 49536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_509
timestamp 1621261055
transform 1 0 50016 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_520
timestamp 1621261055
transform 1 0 51072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_521
timestamp 1621261055
transform 1 0 51168 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_517
timestamp 1621261055
transform 1 0 50784 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_528
timestamp 1621261055
transform 1 0 51840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_524
timestamp 1621261055
transform 1 0 51456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_498
timestamp 1621261055
transform 1 0 51360 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_536
timestamp 1621261055
transform 1 0 52608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_532
timestamp 1621261055
transform 1 0 52224 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_544
timestamp 1621261055
transform 1 0 53376 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_540
timestamp 1621261055
transform 1 0 52992 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_551
timestamp 1621261055
transform 1 0 54048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_548
timestamp 1621261055
transform 1 0 53760 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_548
timestamp 1621261055
transform 1 0 53760 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_509
timestamp 1621261055
transform 1 0 53952 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_559
timestamp 1621261055
transform 1 0 54816 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_556
timestamp 1621261055
transform 1 0 54528 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_567
timestamp 1621261055
transform 1 0 55584 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_564
timestamp 1621261055
transform 1 0 55296 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_575
timestamp 1621261055
transform 1 0 56352 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_576
timestamp 1621261055
transform 1 0 56448 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_572
timestamp 1621261055
transform 1 0 56064 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_499
timestamp 1621261055
transform 1 0 56640 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_583
timestamp 1621261055
transform 1 0 57120 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_586
timestamp 1621261055
transform 1 0 57408 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_579
timestamp 1621261055
transform 1 0 56736 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _150_
timestamp 1621261055
transform 1 0 57120 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_31_591
timestamp 1621261055
transform 1 0 57888 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_594
timestamp 1621261055
transform 1 0 58176 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_61
timestamp 1621261055
transform -1 0 58848 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_63
timestamp 1621261055
transform -1 0 58848 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_30_596
timestamp 1621261055
transform 1 0 58368 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_595
timestamp 1621261055
transform 1 0 58272 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_64
timestamp 1621261055
transform 1 0 1152 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_510
timestamp 1621261055
transform 1 0 3840 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_4
timestamp 1621261055
transform 1 0 1536 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_12
timestamp 1621261055
transform 1 0 2304 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_20
timestamp 1621261055
transform 1 0 3072 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_29
timestamp 1621261055
transform 1 0 3936 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_37
timestamp 1621261055
transform 1 0 4704 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_45
timestamp 1621261055
transform 1 0 5472 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_53
timestamp 1621261055
transform 1 0 6240 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_61
timestamp 1621261055
transform 1 0 7008 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_511
timestamp 1621261055
transform 1 0 9120 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_69
timestamp 1621261055
transform 1 0 7776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_77
timestamp 1621261055
transform 1 0 8544 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_81
timestamp 1621261055
transform 1 0 8928 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_84
timestamp 1621261055
transform 1 0 9216 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_92
timestamp 1621261055
transform 1 0 9984 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_100
timestamp 1621261055
transform 1 0 10752 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_108
timestamp 1621261055
transform 1 0 11520 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_116
timestamp 1621261055
transform 1 0 12288 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_124
timestamp 1621261055
transform 1 0 13056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_132
timestamp 1621261055
transform 1 0 13824 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_512
timestamp 1621261055
transform 1 0 14400 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_136
timestamp 1621261055
transform 1 0 14208 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_139
timestamp 1621261055
transform 1 0 14496 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_147
timestamp 1621261055
transform 1 0 15264 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_155
timestamp 1621261055
transform 1 0 16032 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_163
timestamp 1621261055
transform 1 0 16800 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_513
timestamp 1621261055
transform 1 0 19680 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_171
timestamp 1621261055
transform 1 0 17568 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_179
timestamp 1621261055
transform 1 0 18336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_187
timestamp 1621261055
transform 1 0 19104 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_191
timestamp 1621261055
transform 1 0 19488 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_194
timestamp 1621261055
transform 1 0 19776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_202
timestamp 1621261055
transform 1 0 20544 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_210
timestamp 1621261055
transform 1 0 21312 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_218
timestamp 1621261055
transform 1 0 22080 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_226
timestamp 1621261055
transform 1 0 22848 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_514
timestamp 1621261055
transform 1 0 24960 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_234
timestamp 1621261055
transform 1 0 23616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_242
timestamp 1621261055
transform 1 0 24384 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_246
timestamp 1621261055
transform 1 0 24768 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_249
timestamp 1621261055
transform 1 0 25056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_257
timestamp 1621261055
transform 1 0 25824 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_265
timestamp 1621261055
transform 1 0 26592 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_273
timestamp 1621261055
transform 1 0 27360 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_281
timestamp 1621261055
transform 1 0 28128 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_289
timestamp 1621261055
transform 1 0 28896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_297
timestamp 1621261055
transform 1 0 29664 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_515
timestamp 1621261055
transform 1 0 30240 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_301
timestamp 1621261055
transform 1 0 30048 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_304
timestamp 1621261055
transform 1 0 30336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_312
timestamp 1621261055
transform 1 0 31104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_320
timestamp 1621261055
transform 1 0 31872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_328
timestamp 1621261055
transform 1 0 32640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_516
timestamp 1621261055
transform 1 0 35520 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_336
timestamp 1621261055
transform 1 0 33408 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_344
timestamp 1621261055
transform 1 0 34176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_352
timestamp 1621261055
transform 1 0 34944 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_356
timestamp 1621261055
transform 1 0 35328 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_359
timestamp 1621261055
transform 1 0 35616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_367
timestamp 1621261055
transform 1 0 36384 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_375
timestamp 1621261055
transform 1 0 37152 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_383
timestamp 1621261055
transform 1 0 37920 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_391
timestamp 1621261055
transform 1 0 38688 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_517
timestamp 1621261055
transform 1 0 40800 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_399
timestamp 1621261055
transform 1 0 39456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_407
timestamp 1621261055
transform 1 0 40224 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_411
timestamp 1621261055
transform 1 0 40608 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_414
timestamp 1621261055
transform 1 0 40896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_422
timestamp 1621261055
transform 1 0 41664 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_430
timestamp 1621261055
transform 1 0 42432 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_438
timestamp 1621261055
transform 1 0 43200 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_446
timestamp 1621261055
transform 1 0 43968 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_454
timestamp 1621261055
transform 1 0 44736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_462
timestamp 1621261055
transform 1 0 45504 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_518
timestamp 1621261055
transform 1 0 46080 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_466
timestamp 1621261055
transform 1 0 45888 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_469
timestamp 1621261055
transform 1 0 46176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_477
timestamp 1621261055
transform 1 0 46944 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_485
timestamp 1621261055
transform 1 0 47712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_493
timestamp 1621261055
transform 1 0 48480 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_519
timestamp 1621261055
transform 1 0 51360 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_501
timestamp 1621261055
transform 1 0 49248 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_509
timestamp 1621261055
transform 1 0 50016 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_517
timestamp 1621261055
transform 1 0 50784 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_521
timestamp 1621261055
transform 1 0 51168 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_524
timestamp 1621261055
transform 1 0 51456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_532
timestamp 1621261055
transform 1 0 52224 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_540
timestamp 1621261055
transform 1 0 52992 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_548
timestamp 1621261055
transform 1 0 53760 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_556
timestamp 1621261055
transform 1 0 54528 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_520
timestamp 1621261055
transform 1 0 56640 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_564
timestamp 1621261055
transform 1 0 55296 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_572
timestamp 1621261055
transform 1 0 56064 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_576
timestamp 1621261055
transform 1 0 56448 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_579
timestamp 1621261055
transform 1 0 56736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_587
timestamp 1621261055
transform 1 0 57504 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_65
timestamp 1621261055
transform -1 0 58848 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_595
timestamp 1621261055
transform 1 0 58272 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_66
timestamp 1621261055
transform 1 0 1152 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_4
timestamp 1621261055
transform 1 0 1536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_12
timestamp 1621261055
transform 1 0 2304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_20
timestamp 1621261055
transform 1 0 3072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_28
timestamp 1621261055
transform 1 0 3840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_521
timestamp 1621261055
transform 1 0 6432 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_36
timestamp 1621261055
transform 1 0 4608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_44
timestamp 1621261055
transform 1 0 5376 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_52
timestamp 1621261055
transform 1 0 6144 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_54
timestamp 1621261055
transform 1 0 6336 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_56
timestamp 1621261055
transform 1 0 6528 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_64
timestamp 1621261055
transform 1 0 7296 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_72
timestamp 1621261055
transform 1 0 8064 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_80
timestamp 1621261055
transform 1 0 8832 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_88
timestamp 1621261055
transform 1 0 9600 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_96
timestamp 1621261055
transform 1 0 10368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_522
timestamp 1621261055
transform 1 0 11712 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_104
timestamp 1621261055
transform 1 0 11136 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_108
timestamp 1621261055
transform 1 0 11520 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_111
timestamp 1621261055
transform 1 0 11808 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_119
timestamp 1621261055
transform 1 0 12576 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_127
timestamp 1621261055
transform 1 0 13344 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _096_
timestamp 1621261055
transform 1 0 15456 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_523
timestamp 1621261055
transform 1 0 16992 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_135
timestamp 1621261055
transform 1 0 14112 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_143
timestamp 1621261055
transform 1 0 14880 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_147
timestamp 1621261055
transform 1 0 15264 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_152
timestamp 1621261055
transform 1 0 15744 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_160
timestamp 1621261055
transform 1 0 16512 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_33_164
timestamp 1621261055
transform 1 0 16896 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_166
timestamp 1621261055
transform 1 0 17088 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_174
timestamp 1621261055
transform 1 0 17856 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_182
timestamp 1621261055
transform 1 0 18624 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_190
timestamp 1621261055
transform 1 0 19392 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_198
timestamp 1621261055
transform 1 0 20160 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_524
timestamp 1621261055
transform 1 0 22272 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_206
timestamp 1621261055
transform 1 0 20928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_214
timestamp 1621261055
transform 1 0 21696 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_218
timestamp 1621261055
transform 1 0 22080 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_221
timestamp 1621261055
transform 1 0 22368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_229
timestamp 1621261055
transform 1 0 23136 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_8
timestamp 1621261055
transform 1 0 26496 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_237
timestamp 1621261055
transform 1 0 23904 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_245
timestamp 1621261055
transform 1 0 24672 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_253
timestamp 1621261055
transform 1 0 25440 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_261
timestamp 1621261055
transform 1 0 26208 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_263
timestamp 1621261055
transform 1 0 26400 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _029_
timestamp 1621261055
transform 1 0 26688 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_525
timestamp 1621261055
transform 1 0 27552 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_269
timestamp 1621261055
transform 1 0 26976 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_273
timestamp 1621261055
transform 1 0 27360 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_276
timestamp 1621261055
transform 1 0 27648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_284
timestamp 1621261055
transform 1 0 28416 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_292
timestamp 1621261055
transform 1 0 29184 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_526
timestamp 1621261055
transform 1 0 32832 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_300
timestamp 1621261055
transform 1 0 29952 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_308
timestamp 1621261055
transform 1 0 30720 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_316
timestamp 1621261055
transform 1 0 31488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_324
timestamp 1621261055
transform 1 0 32256 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_328
timestamp 1621261055
transform 1 0 32640 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_331
timestamp 1621261055
transform 1 0 32928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_339
timestamp 1621261055
transform 1 0 33696 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_347
timestamp 1621261055
transform 1 0 34464 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_355
timestamp 1621261055
transform 1 0 35232 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_363
timestamp 1621261055
transform 1 0 36000 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _101_
timestamp 1621261055
transform 1 0 36480 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_527
timestamp 1621261055
transform 1 0 38112 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_33_367
timestamp 1621261055
transform 1 0 36384 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_371
timestamp 1621261055
transform 1 0 36768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_379
timestamp 1621261055
transform 1 0 37536 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_383
timestamp 1621261055
transform 1 0 37920 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_386
timestamp 1621261055
transform 1 0 38208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_394
timestamp 1621261055
transform 1 0 38976 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_402
timestamp 1621261055
transform 1 0 39744 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_410
timestamp 1621261055
transform 1 0 40512 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_418
timestamp 1621261055
transform 1 0 41280 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_426
timestamp 1621261055
transform 1 0 42048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_528
timestamp 1621261055
transform 1 0 43392 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_434
timestamp 1621261055
transform 1 0 42816 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_438
timestamp 1621261055
transform 1 0 43200 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_441
timestamp 1621261055
transform 1 0 43488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_449
timestamp 1621261055
transform 1 0 44256 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_457
timestamp 1621261055
transform 1 0 45024 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_529
timestamp 1621261055
transform 1 0 48672 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_465
timestamp 1621261055
transform 1 0 45792 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_473
timestamp 1621261055
transform 1 0 46560 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_481
timestamp 1621261055
transform 1 0 47328 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_489
timestamp 1621261055
transform 1 0 48096 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_493
timestamp 1621261055
transform 1 0 48480 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_496
timestamp 1621261055
transform 1 0 48768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_504
timestamp 1621261055
transform 1 0 49536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_512
timestamp 1621261055
transform 1 0 50304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_520
timestamp 1621261055
transform 1 0 51072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_528
timestamp 1621261055
transform 1 0 51840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_530
timestamp 1621261055
transform 1 0 53952 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_536
timestamp 1621261055
transform 1 0 52608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_544
timestamp 1621261055
transform 1 0 53376 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_548
timestamp 1621261055
transform 1 0 53760 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_551
timestamp 1621261055
transform 1 0 54048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_559
timestamp 1621261055
transform 1 0 54816 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_567
timestamp 1621261055
transform 1 0 55584 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_575
timestamp 1621261055
transform 1 0 56352 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_583
timestamp 1621261055
transform 1 0 57120 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_591
timestamp 1621261055
transform 1 0 57888 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_67
timestamp 1621261055
transform -1 0 58848 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_595
timestamp 1621261055
transform 1 0 58272 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_68
timestamp 1621261055
transform 1 0 1152 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_531
timestamp 1621261055
transform 1 0 3840 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_36
timestamp 1621261055
transform 1 0 4320 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_4
timestamp 1621261055
transform 1 0 1536 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_12
timestamp 1621261055
transform 1 0 2304 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_20
timestamp 1621261055
transform 1 0 3072 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_29
timestamp 1621261055
transform 1 0 3936 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _045_
timestamp 1621261055
transform 1 0 4512 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _139_
timestamp 1621261055
transform 1 0 5184 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_34_38
timestamp 1621261055
transform 1 0 4800 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_45
timestamp 1621261055
transform 1 0 5472 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_53
timestamp 1621261055
transform 1 0 6240 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_61
timestamp 1621261055
transform 1 0 7008 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_532
timestamp 1621261055
transform 1 0 9120 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_69
timestamp 1621261055
transform 1 0 7776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_77
timestamp 1621261055
transform 1 0 8544 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_81
timestamp 1621261055
transform 1 0 8928 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_84
timestamp 1621261055
transform 1 0 9216 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_92
timestamp 1621261055
transform 1 0 9984 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _041_
timestamp 1621261055
transform 1 0 13632 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_71
timestamp 1621261055
transform 1 0 13440 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_100
timestamp 1621261055
transform 1 0 10752 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_108
timestamp 1621261055
transform 1 0 11520 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_116
timestamp 1621261055
transform 1 0 12288 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_124
timestamp 1621261055
transform 1 0 13056 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_533
timestamp 1621261055
transform 1 0 14400 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_133
timestamp 1621261055
transform 1 0 13920 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_34_137
timestamp 1621261055
transform 1 0 14304 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_139
timestamp 1621261055
transform 1 0 14496 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_147
timestamp 1621261055
transform 1 0 15264 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_155
timestamp 1621261055
transform 1 0 16032 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_163
timestamp 1621261055
transform 1 0 16800 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_534
timestamp 1621261055
transform 1 0 19680 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_171
timestamp 1621261055
transform 1 0 17568 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_179
timestamp 1621261055
transform 1 0 18336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_187
timestamp 1621261055
transform 1 0 19104 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_191
timestamp 1621261055
transform 1 0 19488 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_194
timestamp 1621261055
transform 1 0 19776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_202
timestamp 1621261055
transform 1 0 20544 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_210
timestamp 1621261055
transform 1 0 21312 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_218
timestamp 1621261055
transform 1 0 22080 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_226
timestamp 1621261055
transform 1 0 22848 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_535
timestamp 1621261055
transform 1 0 24960 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_234
timestamp 1621261055
transform 1 0 23616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_242
timestamp 1621261055
transform 1 0 24384 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_246
timestamp 1621261055
transform 1 0 24768 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_249
timestamp 1621261055
transform 1 0 25056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_257
timestamp 1621261055
transform 1 0 25824 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_265
timestamp 1621261055
transform 1 0 26592 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_273
timestamp 1621261055
transform 1 0 27360 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_281
timestamp 1621261055
transform 1 0 28128 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_289
timestamp 1621261055
transform 1 0 28896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_297
timestamp 1621261055
transform 1 0 29664 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_536
timestamp 1621261055
transform 1 0 30240 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_301
timestamp 1621261055
transform 1 0 30048 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_304
timestamp 1621261055
transform 1 0 30336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_312
timestamp 1621261055
transform 1 0 31104 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_320
timestamp 1621261055
transform 1 0 31872 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_328
timestamp 1621261055
transform 1 0 32640 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_537
timestamp 1621261055
transform 1 0 35520 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_336
timestamp 1621261055
transform 1 0 33408 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_344
timestamp 1621261055
transform 1 0 34176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_352
timestamp 1621261055
transform 1 0 34944 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_356
timestamp 1621261055
transform 1 0 35328 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_359
timestamp 1621261055
transform 1 0 35616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_367
timestamp 1621261055
transform 1 0 36384 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_375
timestamp 1621261055
transform 1 0 37152 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_383
timestamp 1621261055
transform 1 0 37920 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_391
timestamp 1621261055
transform 1 0 38688 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _112_
timestamp 1621261055
transform 1 0 39552 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_538
timestamp 1621261055
transform 1 0 40800 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_34_399
timestamp 1621261055
transform 1 0 39456 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_403
timestamp 1621261055
transform 1 0 39840 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_411
timestamp 1621261055
transform 1 0 40608 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_414
timestamp 1621261055
transform 1 0 40896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_422
timestamp 1621261055
transform 1 0 41664 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_430
timestamp 1621261055
transform 1 0 42432 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_438
timestamp 1621261055
transform 1 0 43200 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_446
timestamp 1621261055
transform 1 0 43968 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_454
timestamp 1621261055
transform 1 0 44736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_462
timestamp 1621261055
transform 1 0 45504 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_539
timestamp 1621261055
transform 1 0 46080 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_466
timestamp 1621261055
transform 1 0 45888 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_469
timestamp 1621261055
transform 1 0 46176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_477
timestamp 1621261055
transform 1 0 46944 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_485
timestamp 1621261055
transform 1 0 47712 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_493
timestamp 1621261055
transform 1 0 48480 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_540
timestamp 1621261055
transform 1 0 51360 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_501
timestamp 1621261055
transform 1 0 49248 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_509
timestamp 1621261055
transform 1 0 50016 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_517
timestamp 1621261055
transform 1 0 50784 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_521
timestamp 1621261055
transform 1 0 51168 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_524
timestamp 1621261055
transform 1 0 51456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_532
timestamp 1621261055
transform 1 0 52224 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_540
timestamp 1621261055
transform 1 0 52992 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_548
timestamp 1621261055
transform 1 0 53760 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_556
timestamp 1621261055
transform 1 0 54528 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_541
timestamp 1621261055
transform 1 0 56640 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_564
timestamp 1621261055
transform 1 0 55296 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_572
timestamp 1621261055
transform 1 0 56064 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_576
timestamp 1621261055
transform 1 0 56448 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_579
timestamp 1621261055
transform 1 0 56736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_587
timestamp 1621261055
transform 1 0 57504 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_69
timestamp 1621261055
transform -1 0 58848 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_595
timestamp 1621261055
transform 1 0 58272 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_70
timestamp 1621261055
transform 1 0 1152 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_4
timestamp 1621261055
transform 1 0 1536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_12
timestamp 1621261055
transform 1 0 2304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_20
timestamp 1621261055
transform 1 0 3072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_28
timestamp 1621261055
transform 1 0 3840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_542
timestamp 1621261055
transform 1 0 6432 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_36
timestamp 1621261055
transform 1 0 4608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_44
timestamp 1621261055
transform 1 0 5376 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_52
timestamp 1621261055
transform 1 0 6144 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_54
timestamp 1621261055
transform 1 0 6336 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_56
timestamp 1621261055
transform 1 0 6528 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_64
timestamp 1621261055
transform 1 0 7296 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_72
timestamp 1621261055
transform 1 0 8064 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_80
timestamp 1621261055
transform 1 0 8832 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_88
timestamp 1621261055
transform 1 0 9600 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_96
timestamp 1621261055
transform 1 0 10368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_543
timestamp 1621261055
transform 1 0 11712 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_104
timestamp 1621261055
transform 1 0 11136 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_108
timestamp 1621261055
transform 1 0 11520 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_111
timestamp 1621261055
transform 1 0 11808 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_119
timestamp 1621261055
transform 1 0 12576 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_127
timestamp 1621261055
transform 1 0 13344 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_544
timestamp 1621261055
transform 1 0 16992 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_135
timestamp 1621261055
transform 1 0 14112 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_143
timestamp 1621261055
transform 1 0 14880 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_151
timestamp 1621261055
transform 1 0 15648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_159
timestamp 1621261055
transform 1 0 16416 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_163
timestamp 1621261055
transform 1 0 16800 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_166
timestamp 1621261055
transform 1 0 17088 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_174
timestamp 1621261055
transform 1 0 17856 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_182
timestamp 1621261055
transform 1 0 18624 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_190
timestamp 1621261055
transform 1 0 19392 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_198
timestamp 1621261055
transform 1 0 20160 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_545
timestamp 1621261055
transform 1 0 22272 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_206
timestamp 1621261055
transform 1 0 20928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_214
timestamp 1621261055
transform 1 0 21696 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_218
timestamp 1621261055
transform 1 0 22080 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_221
timestamp 1621261055
transform 1 0 22368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_229
timestamp 1621261055
transform 1 0 23136 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_237
timestamp 1621261055
transform 1 0 23904 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_245
timestamp 1621261055
transform 1 0 24672 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_253
timestamp 1621261055
transform 1 0 25440 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_261
timestamp 1621261055
transform 1 0 26208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_546
timestamp 1621261055
transform 1 0 27552 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_269
timestamp 1621261055
transform 1 0 26976 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_273
timestamp 1621261055
transform 1 0 27360 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_276
timestamp 1621261055
transform 1 0 27648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_284
timestamp 1621261055
transform 1 0 28416 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_292
timestamp 1621261055
transform 1 0 29184 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_547
timestamp 1621261055
transform 1 0 32832 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_300
timestamp 1621261055
transform 1 0 29952 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_308
timestamp 1621261055
transform 1 0 30720 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_316
timestamp 1621261055
transform 1 0 31488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_324
timestamp 1621261055
transform 1 0 32256 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_328
timestamp 1621261055
transform 1 0 32640 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_331
timestamp 1621261055
transform 1 0 32928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_339
timestamp 1621261055
transform 1 0 33696 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_347
timestamp 1621261055
transform 1 0 34464 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_355
timestamp 1621261055
transform 1 0 35232 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_363
timestamp 1621261055
transform 1 0 36000 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_548
timestamp 1621261055
transform 1 0 38112 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_371
timestamp 1621261055
transform 1 0 36768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_379
timestamp 1621261055
transform 1 0 37536 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_383
timestamp 1621261055
transform 1 0 37920 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_386
timestamp 1621261055
transform 1 0 38208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_394
timestamp 1621261055
transform 1 0 38976 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _155_
timestamp 1621261055
transform 1 0 39936 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_402
timestamp 1621261055
transform 1 0 39744 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_407
timestamp 1621261055
transform 1 0 40224 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_415
timestamp 1621261055
transform 1 0 40992 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_423
timestamp 1621261055
transform 1 0 41760 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_549
timestamp 1621261055
transform 1 0 43392 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_431
timestamp 1621261055
transform 1 0 42528 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_35_439
timestamp 1621261055
transform 1 0 43296 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_441
timestamp 1621261055
transform 1 0 43488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_449
timestamp 1621261055
transform 1 0 44256 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_457
timestamp 1621261055
transform 1 0 45024 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _154_
timestamp 1621261055
transform 1 0 47520 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_550
timestamp 1621261055
transform 1 0 48672 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_465
timestamp 1621261055
transform 1 0 45792 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_473
timestamp 1621261055
transform 1 0 46560 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_481
timestamp 1621261055
transform 1 0 47328 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_486
timestamp 1621261055
transform 1 0 47808 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_35_494
timestamp 1621261055
transform 1 0 48576 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_496
timestamp 1621261055
transform 1 0 48768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_504
timestamp 1621261055
transform 1 0 49536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_512
timestamp 1621261055
transform 1 0 50304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_520
timestamp 1621261055
transform 1 0 51072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_528
timestamp 1621261055
transform 1 0 51840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _128_
timestamp 1621261055
transform 1 0 54432 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_551
timestamp 1621261055
transform 1 0 53952 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_536
timestamp 1621261055
transform 1 0 52608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_544
timestamp 1621261055
transform 1 0 53376 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_548
timestamp 1621261055
transform 1 0 53760 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_35_551
timestamp 1621261055
transform 1 0 54048 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_558
timestamp 1621261055
transform 1 0 54720 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_566
timestamp 1621261055
transform 1 0 55488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_574
timestamp 1621261055
transform 1 0 56256 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_582
timestamp 1621261055
transform 1 0 57024 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_590
timestamp 1621261055
transform 1 0 57792 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_594
timestamp 1621261055
transform 1 0 58176 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_71
timestamp 1621261055
transform -1 0 58848 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_35_596
timestamp 1621261055
transform 1 0 58368 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_72
timestamp 1621261055
transform 1 0 1152 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_552
timestamp 1621261055
transform 1 0 3840 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_4
timestamp 1621261055
transform 1 0 1536 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_12
timestamp 1621261055
transform 1 0 2304 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_20
timestamp 1621261055
transform 1 0 3072 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_29
timestamp 1621261055
transform 1 0 3936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_37
timestamp 1621261055
transform 1 0 4704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_45
timestamp 1621261055
transform 1 0 5472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_53
timestamp 1621261055
transform 1 0 6240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_61
timestamp 1621261055
transform 1 0 7008 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_553
timestamp 1621261055
transform 1 0 9120 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_69
timestamp 1621261055
transform 1 0 7776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_77
timestamp 1621261055
transform 1 0 8544 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_81
timestamp 1621261055
transform 1 0 8928 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_84
timestamp 1621261055
transform 1 0 9216 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_92
timestamp 1621261055
transform 1 0 9984 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _148_
timestamp 1621261055
transform 1 0 12288 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_36_100
timestamp 1621261055
transform 1 0 10752 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_108
timestamp 1621261055
transform 1 0 11520 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_119
timestamp 1621261055
transform 1 0 12576 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_127
timestamp 1621261055
transform 1 0 13344 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_554
timestamp 1621261055
transform 1 0 14400 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_135
timestamp 1621261055
transform 1 0 14112 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_36_137
timestamp 1621261055
transform 1 0 14304 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_139
timestamp 1621261055
transform 1 0 14496 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_147
timestamp 1621261055
transform 1 0 15264 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_155
timestamp 1621261055
transform 1 0 16032 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_163
timestamp 1621261055
transform 1 0 16800 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_555
timestamp 1621261055
transform 1 0 19680 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_171
timestamp 1621261055
transform 1 0 17568 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_179
timestamp 1621261055
transform 1 0 18336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_187
timestamp 1621261055
transform 1 0 19104 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_191
timestamp 1621261055
transform 1 0 19488 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_194
timestamp 1621261055
transform 1 0 19776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_202
timestamp 1621261055
transform 1 0 20544 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_210
timestamp 1621261055
transform 1 0 21312 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_218
timestamp 1621261055
transform 1 0 22080 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_226
timestamp 1621261055
transform 1 0 22848 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_556
timestamp 1621261055
transform 1 0 24960 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_234
timestamp 1621261055
transform 1 0 23616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_242
timestamp 1621261055
transform 1 0 24384 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_246
timestamp 1621261055
transform 1 0 24768 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_249
timestamp 1621261055
transform 1 0 25056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_257
timestamp 1621261055
transform 1 0 25824 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_265
timestamp 1621261055
transform 1 0 26592 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_273
timestamp 1621261055
transform 1 0 27360 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_281
timestamp 1621261055
transform 1 0 28128 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_289
timestamp 1621261055
transform 1 0 28896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_297
timestamp 1621261055
transform 1 0 29664 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_557
timestamp 1621261055
transform 1 0 30240 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_301
timestamp 1621261055
transform 1 0 30048 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_304
timestamp 1621261055
transform 1 0 30336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_312
timestamp 1621261055
transform 1 0 31104 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_320
timestamp 1621261055
transform 1 0 31872 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_328
timestamp 1621261055
transform 1 0 32640 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_558
timestamp 1621261055
transform 1 0 35520 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_336
timestamp 1621261055
transform 1 0 33408 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_344
timestamp 1621261055
transform 1 0 34176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_352
timestamp 1621261055
transform 1 0 34944 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_356
timestamp 1621261055
transform 1 0 35328 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_359
timestamp 1621261055
transform 1 0 35616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _052_
timestamp 1621261055
transform 1 0 37824 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_53
timestamp 1621261055
transform 1 0 37632 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_367
timestamp 1621261055
transform 1 0 36384 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_375
timestamp 1621261055
transform 1 0 37152 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_36_379
timestamp 1621261055
transform 1 0 37536 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_385
timestamp 1621261055
transform 1 0 38112 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_393
timestamp 1621261055
transform 1 0 38880 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_559
timestamp 1621261055
transform 1 0 40800 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_401
timestamp 1621261055
transform 1 0 39648 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_409
timestamp 1621261055
transform 1 0 40416 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_414
timestamp 1621261055
transform 1 0 40896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_422
timestamp 1621261055
transform 1 0 41664 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_430
timestamp 1621261055
transform 1 0 42432 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_438
timestamp 1621261055
transform 1 0 43200 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_446
timestamp 1621261055
transform 1 0 43968 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_454
timestamp 1621261055
transform 1 0 44736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_462
timestamp 1621261055
transform 1 0 45504 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_560
timestamp 1621261055
transform 1 0 46080 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_466
timestamp 1621261055
transform 1 0 45888 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_469
timestamp 1621261055
transform 1 0 46176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_477
timestamp 1621261055
transform 1 0 46944 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_485
timestamp 1621261055
transform 1 0 47712 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_493
timestamp 1621261055
transform 1 0 48480 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_561
timestamp 1621261055
transform 1 0 51360 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_501
timestamp 1621261055
transform 1 0 49248 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_509
timestamp 1621261055
transform 1 0 50016 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_517
timestamp 1621261055
transform 1 0 50784 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_521
timestamp 1621261055
transform 1 0 51168 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_524
timestamp 1621261055
transform 1 0 51456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_532
timestamp 1621261055
transform 1 0 52224 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_540
timestamp 1621261055
transform 1 0 52992 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_548
timestamp 1621261055
transform 1 0 53760 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_556
timestamp 1621261055
transform 1 0 54528 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_562
timestamp 1621261055
transform 1 0 56640 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_564
timestamp 1621261055
transform 1 0 55296 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_572
timestamp 1621261055
transform 1 0 56064 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_576
timestamp 1621261055
transform 1 0 56448 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_579
timestamp 1621261055
transform 1 0 56736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_587
timestamp 1621261055
transform 1 0 57504 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_73
timestamp 1621261055
transform -1 0 58848 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_595
timestamp 1621261055
transform 1 0 58272 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_74
timestamp 1621261055
transform 1 0 1152 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_4
timestamp 1621261055
transform 1 0 1536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_12
timestamp 1621261055
transform 1 0 2304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_20
timestamp 1621261055
transform 1 0 3072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_28
timestamp 1621261055
transform 1 0 3840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_563
timestamp 1621261055
transform 1 0 6432 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_36
timestamp 1621261055
transform 1 0 4608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_44
timestamp 1621261055
transform 1 0 5376 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_52
timestamp 1621261055
transform 1 0 6144 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_54
timestamp 1621261055
transform 1 0 6336 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_56
timestamp 1621261055
transform 1 0 6528 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_64
timestamp 1621261055
transform 1 0 7296 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_72
timestamp 1621261055
transform 1 0 8064 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_80
timestamp 1621261055
transform 1 0 8832 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_88
timestamp 1621261055
transform 1 0 9600 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_96
timestamp 1621261055
transform 1 0 10368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_564
timestamp 1621261055
transform 1 0 11712 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_104
timestamp 1621261055
transform 1 0 11136 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_108
timestamp 1621261055
transform 1 0 11520 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_111
timestamp 1621261055
transform 1 0 11808 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_119
timestamp 1621261055
transform 1 0 12576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_127
timestamp 1621261055
transform 1 0 13344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_565
timestamp 1621261055
transform 1 0 16992 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_135
timestamp 1621261055
transform 1 0 14112 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_143
timestamp 1621261055
transform 1 0 14880 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_151
timestamp 1621261055
transform 1 0 15648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_159
timestamp 1621261055
transform 1 0 16416 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_163
timestamp 1621261055
transform 1 0 16800 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_166
timestamp 1621261055
transform 1 0 17088 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_174
timestamp 1621261055
transform 1 0 17856 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_182
timestamp 1621261055
transform 1 0 18624 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_190
timestamp 1621261055
transform 1 0 19392 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_198
timestamp 1621261055
transform 1 0 20160 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_566
timestamp 1621261055
transform 1 0 22272 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_206
timestamp 1621261055
transform 1 0 20928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_214
timestamp 1621261055
transform 1 0 21696 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_218
timestamp 1621261055
transform 1 0 22080 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_221
timestamp 1621261055
transform 1 0 22368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_229
timestamp 1621261055
transform 1 0 23136 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_237
timestamp 1621261055
transform 1 0 23904 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_245
timestamp 1621261055
transform 1 0 24672 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_253
timestamp 1621261055
transform 1 0 25440 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_261
timestamp 1621261055
transform 1 0 26208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_567
timestamp 1621261055
transform 1 0 27552 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_269
timestamp 1621261055
transform 1 0 26976 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_273
timestamp 1621261055
transform 1 0 27360 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_276
timestamp 1621261055
transform 1 0 27648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_284
timestamp 1621261055
transform 1 0 28416 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_292
timestamp 1621261055
transform 1 0 29184 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_568
timestamp 1621261055
transform 1 0 32832 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_300
timestamp 1621261055
transform 1 0 29952 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_308
timestamp 1621261055
transform 1 0 30720 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_316
timestamp 1621261055
transform 1 0 31488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_324
timestamp 1621261055
transform 1 0 32256 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_328
timestamp 1621261055
transform 1 0 32640 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_331
timestamp 1621261055
transform 1 0 32928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_339
timestamp 1621261055
transform 1 0 33696 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_347
timestamp 1621261055
transform 1 0 34464 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_355
timestamp 1621261055
transform 1 0 35232 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_363
timestamp 1621261055
transform 1 0 36000 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_569
timestamp 1621261055
transform 1 0 38112 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_371
timestamp 1621261055
transform 1 0 36768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_379
timestamp 1621261055
transform 1 0 37536 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_383
timestamp 1621261055
transform 1 0 37920 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_386
timestamp 1621261055
transform 1 0 38208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_394
timestamp 1621261055
transform 1 0 38976 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_402
timestamp 1621261055
transform 1 0 39744 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_410
timestamp 1621261055
transform 1 0 40512 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_418
timestamp 1621261055
transform 1 0 41280 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_426
timestamp 1621261055
transform 1 0 42048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_570
timestamp 1621261055
transform 1 0 43392 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_434
timestamp 1621261055
transform 1 0 42816 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_438
timestamp 1621261055
transform 1 0 43200 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_441
timestamp 1621261055
transform 1 0 43488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_449
timestamp 1621261055
transform 1 0 44256 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_457
timestamp 1621261055
transform 1 0 45024 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_571
timestamp 1621261055
transform 1 0 48672 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_465
timestamp 1621261055
transform 1 0 45792 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_473
timestamp 1621261055
transform 1 0 46560 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_481
timestamp 1621261055
transform 1 0 47328 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_489
timestamp 1621261055
transform 1 0 48096 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_493
timestamp 1621261055
transform 1 0 48480 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_496
timestamp 1621261055
transform 1 0 48768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_504
timestamp 1621261055
transform 1 0 49536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_512
timestamp 1621261055
transform 1 0 50304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_520
timestamp 1621261055
transform 1 0 51072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_528
timestamp 1621261055
transform 1 0 51840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_572
timestamp 1621261055
transform 1 0 53952 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_536
timestamp 1621261055
transform 1 0 52608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_544
timestamp 1621261055
transform 1 0 53376 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_548
timestamp 1621261055
transform 1 0 53760 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_551
timestamp 1621261055
transform 1 0 54048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_559
timestamp 1621261055
transform 1 0 54816 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_567
timestamp 1621261055
transform 1 0 55584 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_575
timestamp 1621261055
transform 1 0 56352 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_583
timestamp 1621261055
transform 1 0 57120 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_591
timestamp 1621261055
transform 1 0 57888 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_75
timestamp 1621261055
transform -1 0 58848 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_595
timestamp 1621261055
transform 1 0 58272 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_4
timestamp 1621261055
transform 1 0 1536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_4
timestamp 1621261055
transform 1 0 1536 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_78
timestamp 1621261055
transform 1 0 1152 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_76
timestamp 1621261055
transform 1 0 1152 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_12
timestamp 1621261055
transform 1 0 2304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_12
timestamp 1621261055
transform 1 0 2304 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_20
timestamp 1621261055
transform 1 0 3072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_20
timestamp 1621261055
transform 1 0 3072 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_28
timestamp 1621261055
transform 1 0 3840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_29
timestamp 1621261055
transform 1 0 3936 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_573
timestamp 1621261055
transform 1 0 3840 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_36
timestamp 1621261055
transform 1 0 4608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_37
timestamp 1621261055
transform 1 0 4704 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_44
timestamp 1621261055
transform 1 0 5376 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_49
timestamp 1621261055
transform 1 0 5856 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_45
timestamp 1621261055
transform 1 0 5472 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_56
timestamp 1621261055
transform 1 0 6528 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_54
timestamp 1621261055
transform 1 0 6336 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_52
timestamp 1621261055
transform 1 0 6144 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_54
timestamp 1621261055
transform 1 0 6336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_584
timestamp 1621261055
transform 1 0 6432 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _180_
timestamp 1621261055
transform 1 0 6048 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_64
timestamp 1621261055
transform 1 0 7296 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_62
timestamp 1621261055
transform 1 0 7104 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_72
timestamp 1621261055
transform 1 0 8064 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_70
timestamp 1621261055
transform 1 0 7872 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_80
timestamp 1621261055
transform 1 0 8832 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_38_82
timestamp 1621261055
transform 1 0 9024 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_78
timestamp 1621261055
transform 1 0 8640 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_98
timestamp 1621261055
transform 1 0 8928 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_574
timestamp 1621261055
transform 1 0 9120 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _178_
timestamp 1621261055
transform 1 0 9120 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_86
timestamp 1621261055
transform 1 0 9408 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_92
timestamp 1621261055
transform 1 0 9984 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_84
timestamp 1621261055
transform 1 0 9216 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_94
timestamp 1621261055
transform 1 0 10176 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_102
timestamp 1621261055
transform 1 0 10944 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_100
timestamp 1621261055
transform 1 0 10752 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_111
timestamp 1621261055
transform 1 0 11808 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_116
timestamp 1621261055
transform 1 0 12288 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_108
timestamp 1621261055
transform 1 0 11520 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_585
timestamp 1621261055
transform 1 0 11712 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_119
timestamp 1621261055
transform 1 0 12576 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_124
timestamp 1621261055
transform 1 0 13056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_127
timestamp 1621261055
transform 1 0 13344 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_132
timestamp 1621261055
transform 1 0 13824 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_135
timestamp 1621261055
transform 1 0 14112 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_139
timestamp 1621261055
transform 1 0 14496 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_136
timestamp 1621261055
transform 1 0 14208 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_575
timestamp 1621261055
transform 1 0 14400 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_143
timestamp 1621261055
transform 1 0 14880 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_147
timestamp 1621261055
transform 1 0 15264 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_151
timestamp 1621261055
transform 1 0 15648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_155
timestamp 1621261055
transform 1 0 16032 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_163
timestamp 1621261055
transform 1 0 16800 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_159
timestamp 1621261055
transform 1 0 16416 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_163
timestamp 1621261055
transform 1 0 16800 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_586
timestamp 1621261055
transform 1 0 16992 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_166
timestamp 1621261055
transform 1 0 17088 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_171
timestamp 1621261055
transform 1 0 17568 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_182
timestamp 1621261055
transform 1 0 18624 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_174
timestamp 1621261055
transform 1 0 17856 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_179
timestamp 1621261055
transform 1 0 18336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_190
timestamp 1621261055
transform 1 0 19392 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_191
timestamp 1621261055
transform 1 0 19488 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_187
timestamp 1621261055
transform 1 0 19104 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_198
timestamp 1621261055
transform 1 0 20160 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_194
timestamp 1621261055
transform 1 0 19776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_576
timestamp 1621261055
transform 1 0 19680 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_206
timestamp 1621261055
transform 1 0 20928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_202
timestamp 1621261055
transform 1 0 20544 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_214
timestamp 1621261055
transform 1 0 21696 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_210
timestamp 1621261055
transform 1 0 21312 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_221
timestamp 1621261055
transform 1 0 22368 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_218
timestamp 1621261055
transform 1 0 22080 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_218
timestamp 1621261055
transform 1 0 22080 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_587
timestamp 1621261055
transform 1 0 22272 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_229
timestamp 1621261055
transform 1 0 23136 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_226
timestamp 1621261055
transform 1 0 22848 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_237
timestamp 1621261055
transform 1 0 23904 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_234
timestamp 1621261055
transform 1 0 23616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_245
timestamp 1621261055
transform 1 0 24672 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_246
timestamp 1621261055
transform 1 0 24768 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_242
timestamp 1621261055
transform 1 0 24384 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_577
timestamp 1621261055
transform 1 0 24960 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_253
timestamp 1621261055
transform 1 0 25440 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_257
timestamp 1621261055
transform 1 0 25824 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_249
timestamp 1621261055
transform 1 0 25056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_261
timestamp 1621261055
transform 1 0 26208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_269
timestamp 1621261055
transform 1 0 26976 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_265
timestamp 1621261055
transform 1 0 26592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_276
timestamp 1621261055
transform 1 0 27648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_273
timestamp 1621261055
transform 1 0 27360 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_281
timestamp 1621261055
transform 1 0 28128 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_273
timestamp 1621261055
transform 1 0 27360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_588
timestamp 1621261055
transform 1 0 27552 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_290
timestamp 1621261055
transform 1 0 28992 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_286
timestamp 1621261055
transform 1 0 28608 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_284
timestamp 1621261055
transform 1 0 28416 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_289
timestamp 1621261055
transform 1 0 28896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _075_
timestamp 1621261055
transform 1 0 28704 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_38_297
timestamp 1621261055
transform 1 0 29664 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_298
timestamp 1621261055
transform 1 0 29760 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_304
timestamp 1621261055
transform 1 0 30336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_301
timestamp 1621261055
transform 1 0 30048 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_578
timestamp 1621261055
transform 1 0 30240 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_314
timestamp 1621261055
transform 1 0 31296 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_306
timestamp 1621261055
transform 1 0 30528 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_312
timestamp 1621261055
transform 1 0 31104 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_322
timestamp 1621261055
transform 1 0 32064 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_320
timestamp 1621261055
transform 1 0 31872 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_328
timestamp 1621261055
transform 1 0 32640 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_589
timestamp 1621261055
transform 1 0 32832 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_331
timestamp 1621261055
transform 1 0 32928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_336
timestamp 1621261055
transform 1 0 33408 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_347
timestamp 1621261055
transform 1 0 34464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_339
timestamp 1621261055
transform 1 0 33696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_344
timestamp 1621261055
transform 1 0 34176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_355
timestamp 1621261055
transform 1 0 35232 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_356
timestamp 1621261055
transform 1 0 35328 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_352
timestamp 1621261055
transform 1 0 34944 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_363
timestamp 1621261055
transform 1 0 36000 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_359
timestamp 1621261055
transform 1 0 35616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_579
timestamp 1621261055
transform 1 0 35520 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_371
timestamp 1621261055
transform 1 0 36768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_367
timestamp 1621261055
transform 1 0 36384 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_379
timestamp 1621261055
transform 1 0 37536 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_375
timestamp 1621261055
transform 1 0 37152 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_386
timestamp 1621261055
transform 1 0 38208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_383
timestamp 1621261055
transform 1 0 37920 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_388
timestamp 1621261055
transform 1 0 38400 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_0
timestamp 1621261055
transform 1 0 37920 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_590
timestamp 1621261055
transform 1 0 38112 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _022_
timestamp 1621261055
transform 1 0 38112 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_394
timestamp 1621261055
transform 1 0 38976 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_396
timestamp 1621261055
transform 1 0 39168 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_580
timestamp 1621261055
transform 1 0 40800 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_404
timestamp 1621261055
transform 1 0 39936 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_38_412
timestamp 1621261055
transform 1 0 40704 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_414
timestamp 1621261055
transform 1 0 40896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_422
timestamp 1621261055
transform 1 0 41664 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_402
timestamp 1621261055
transform 1 0 39744 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_410
timestamp 1621261055
transform 1 0 40512 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_418
timestamp 1621261055
transform 1 0 41280 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_426
timestamp 1621261055
transform 1 0 42048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_434
timestamp 1621261055
transform 1 0 42816 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_430
timestamp 1621261055
transform 1 0 42432 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_441
timestamp 1621261055
transform 1 0 43488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_438
timestamp 1621261055
transform 1 0 43200 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_446
timestamp 1621261055
transform 1 0 43968 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_438
timestamp 1621261055
transform 1 0 43200 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_591
timestamp 1621261055
transform 1 0 43392 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_449
timestamp 1621261055
transform 1 0 44256 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_454
timestamp 1621261055
transform 1 0 44736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_457
timestamp 1621261055
transform 1 0 45024 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_462
timestamp 1621261055
transform 1 0 45504 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_465
timestamp 1621261055
transform 1 0 45792 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_469
timestamp 1621261055
transform 1 0 46176 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_466
timestamp 1621261055
transform 1 0 45888 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_581
timestamp 1621261055
transform 1 0 46080 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_473
timestamp 1621261055
transform 1 0 46560 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_476
timestamp 1621261055
transform 1 0 46848 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_51
timestamp 1621261055
transform -1 0 46560 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _050_
timestamp 1621261055
transform -1 0 46848 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_481
timestamp 1621261055
transform 1 0 47328 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_484
timestamp 1621261055
transform 1 0 47616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_493
timestamp 1621261055
transform 1 0 48480 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_489
timestamp 1621261055
transform 1 0 48096 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_492
timestamp 1621261055
transform 1 0 48384 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_592
timestamp 1621261055
transform 1 0 48672 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_496
timestamp 1621261055
transform 1 0 48768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_500
timestamp 1621261055
transform 1 0 49152 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_512
timestamp 1621261055
transform 1 0 50304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_504
timestamp 1621261055
transform 1 0 49536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_508
timestamp 1621261055
transform 1 0 49920 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_520
timestamp 1621261055
transform 1 0 51072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_520
timestamp 1621261055
transform 1 0 51072 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_516
timestamp 1621261055
transform 1 0 50688 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_528
timestamp 1621261055
transform 1 0 51840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_524
timestamp 1621261055
transform 1 0 51456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_38_522
timestamp 1621261055
transform 1 0 51264 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_582
timestamp 1621261055
transform 1 0 51360 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_536
timestamp 1621261055
transform 1 0 52608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_532
timestamp 1621261055
transform 1 0 52224 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_544
timestamp 1621261055
transform 1 0 53376 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_540
timestamp 1621261055
transform 1 0 52992 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_551
timestamp 1621261055
transform 1 0 54048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_548
timestamp 1621261055
transform 1 0 53760 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_548
timestamp 1621261055
transform 1 0 53760 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_593
timestamp 1621261055
transform 1 0 53952 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_559
timestamp 1621261055
transform 1 0 54816 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_556
timestamp 1621261055
transform 1 0 54528 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_567
timestamp 1621261055
transform 1 0 55584 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_564
timestamp 1621261055
transform 1 0 55296 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_575
timestamp 1621261055
transform 1 0 56352 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_576
timestamp 1621261055
transform 1 0 56448 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_572
timestamp 1621261055
transform 1 0 56064 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_583
timestamp 1621261055
transform 1 0 56640 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_583
timestamp 1621261055
transform 1 0 57120 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_586
timestamp 1621261055
transform 1 0 57408 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_38_579
timestamp 1621261055
transform 1 0 56736 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _169_
timestamp 1621261055
transform 1 0 57120 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_39_591
timestamp 1621261055
transform 1 0 57888 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_38_593
timestamp 1621261055
transform 1 0 58080 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _088_
timestamp 1621261055
transform 1 0 57792 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_77
timestamp 1621261055
transform -1 0 58848 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_79
timestamp 1621261055
transform -1 0 58848 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_595
timestamp 1621261055
transform 1 0 58272 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_80
timestamp 1621261055
transform 1 0 1152 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_594
timestamp 1621261055
transform 1 0 3840 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_4
timestamp 1621261055
transform 1 0 1536 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_12
timestamp 1621261055
transform 1 0 2304 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_20
timestamp 1621261055
transform 1 0 3072 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_29
timestamp 1621261055
transform 1 0 3936 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_37
timestamp 1621261055
transform 1 0 4704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_45
timestamp 1621261055
transform 1 0 5472 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_53
timestamp 1621261055
transform 1 0 6240 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_61
timestamp 1621261055
transform 1 0 7008 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_595
timestamp 1621261055
transform 1 0 9120 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_69
timestamp 1621261055
transform 1 0 7776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_77
timestamp 1621261055
transform 1 0 8544 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_81
timestamp 1621261055
transform 1 0 8928 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_84
timestamp 1621261055
transform 1 0 9216 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_92
timestamp 1621261055
transform 1 0 9984 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_100
timestamp 1621261055
transform 1 0 10752 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_108
timestamp 1621261055
transform 1 0 11520 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_116
timestamp 1621261055
transform 1 0 12288 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_124
timestamp 1621261055
transform 1 0 13056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_132
timestamp 1621261055
transform 1 0 13824 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_596
timestamp 1621261055
transform 1 0 14400 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_136
timestamp 1621261055
transform 1 0 14208 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_139
timestamp 1621261055
transform 1 0 14496 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_147
timestamp 1621261055
transform 1 0 15264 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_155
timestamp 1621261055
transform 1 0 16032 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_163
timestamp 1621261055
transform 1 0 16800 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_597
timestamp 1621261055
transform 1 0 19680 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_171
timestamp 1621261055
transform 1 0 17568 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_179
timestamp 1621261055
transform 1 0 18336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_187
timestamp 1621261055
transform 1 0 19104 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_191
timestamp 1621261055
transform 1 0 19488 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_194
timestamp 1621261055
transform 1 0 19776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_202
timestamp 1621261055
transform 1 0 20544 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_210
timestamp 1621261055
transform 1 0 21312 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_218
timestamp 1621261055
transform 1 0 22080 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_226
timestamp 1621261055
transform 1 0 22848 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_598
timestamp 1621261055
transform 1 0 24960 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_234
timestamp 1621261055
transform 1 0 23616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_242
timestamp 1621261055
transform 1 0 24384 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_246
timestamp 1621261055
transform 1 0 24768 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_249
timestamp 1621261055
transform 1 0 25056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_257
timestamp 1621261055
transform 1 0 25824 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _030_
timestamp 1621261055
transform 1 0 28032 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_10
timestamp 1621261055
transform 1 0 27840 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_265
timestamp 1621261055
transform 1 0 26592 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_273
timestamp 1621261055
transform 1 0 27360 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_40_277
timestamp 1621261055
transform 1 0 27744 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_283
timestamp 1621261055
transform 1 0 28320 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_291
timestamp 1621261055
transform 1 0 29088 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_599
timestamp 1621261055
transform 1 0 30240 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_299
timestamp 1621261055
transform 1 0 29856 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_40_304
timestamp 1621261055
transform 1 0 30336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_312
timestamp 1621261055
transform 1 0 31104 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_320
timestamp 1621261055
transform 1 0 31872 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_328
timestamp 1621261055
transform 1 0 32640 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_600
timestamp 1621261055
transform 1 0 35520 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_336
timestamp 1621261055
transform 1 0 33408 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_344
timestamp 1621261055
transform 1 0 34176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_352
timestamp 1621261055
transform 1 0 34944 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_356
timestamp 1621261055
transform 1 0 35328 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_359
timestamp 1621261055
transform 1 0 35616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_367
timestamp 1621261055
transform 1 0 36384 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_375
timestamp 1621261055
transform 1 0 37152 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_383
timestamp 1621261055
transform 1 0 37920 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_391
timestamp 1621261055
transform 1 0 38688 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_601
timestamp 1621261055
transform 1 0 40800 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_399
timestamp 1621261055
transform 1 0 39456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_407
timestamp 1621261055
transform 1 0 40224 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_411
timestamp 1621261055
transform 1 0 40608 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_414
timestamp 1621261055
transform 1 0 40896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_422
timestamp 1621261055
transform 1 0 41664 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_430
timestamp 1621261055
transform 1 0 42432 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_438
timestamp 1621261055
transform 1 0 43200 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_446
timestamp 1621261055
transform 1 0 43968 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_454
timestamp 1621261055
transform 1 0 44736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_462
timestamp 1621261055
transform 1 0 45504 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_602
timestamp 1621261055
transform 1 0 46080 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_466
timestamp 1621261055
transform 1 0 45888 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_469
timestamp 1621261055
transform 1 0 46176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_477
timestamp 1621261055
transform 1 0 46944 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_485
timestamp 1621261055
transform 1 0 47712 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_493
timestamp 1621261055
transform 1 0 48480 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_603
timestamp 1621261055
transform 1 0 51360 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_501
timestamp 1621261055
transform 1 0 49248 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_509
timestamp 1621261055
transform 1 0 50016 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_517
timestamp 1621261055
transform 1 0 50784 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_521
timestamp 1621261055
transform 1 0 51168 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_524
timestamp 1621261055
transform 1 0 51456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_532
timestamp 1621261055
transform 1 0 52224 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_540
timestamp 1621261055
transform 1 0 52992 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_548
timestamp 1621261055
transform 1 0 53760 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_556
timestamp 1621261055
transform 1 0 54528 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_604
timestamp 1621261055
transform 1 0 56640 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_564
timestamp 1621261055
transform 1 0 55296 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_572
timestamp 1621261055
transform 1 0 56064 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_576
timestamp 1621261055
transform 1 0 56448 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_579
timestamp 1621261055
transform 1 0 56736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_587
timestamp 1621261055
transform 1 0 57504 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_81
timestamp 1621261055
transform -1 0 58848 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_595
timestamp 1621261055
transform 1 0 58272 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_82
timestamp 1621261055
transform 1 0 1152 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_4
timestamp 1621261055
transform 1 0 1536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_12
timestamp 1621261055
transform 1 0 2304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_20
timestamp 1621261055
transform 1 0 3072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_28
timestamp 1621261055
transform 1 0 3840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_605
timestamp 1621261055
transform 1 0 6432 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_36
timestamp 1621261055
transform 1 0 4608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_44
timestamp 1621261055
transform 1 0 5376 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_52
timestamp 1621261055
transform 1 0 6144 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_41_54
timestamp 1621261055
transform 1 0 6336 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_56
timestamp 1621261055
transform 1 0 6528 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_64
timestamp 1621261055
transform 1 0 7296 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_72
timestamp 1621261055
transform 1 0 8064 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_80
timestamp 1621261055
transform 1 0 8832 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_88
timestamp 1621261055
transform 1 0 9600 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_96
timestamp 1621261055
transform 1 0 10368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_606
timestamp 1621261055
transform 1 0 11712 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_104
timestamp 1621261055
transform 1 0 11136 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_108
timestamp 1621261055
transform 1 0 11520 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_111
timestamp 1621261055
transform 1 0 11808 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_119
timestamp 1621261055
transform 1 0 12576 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_127
timestamp 1621261055
transform 1 0 13344 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_607
timestamp 1621261055
transform 1 0 16992 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_135
timestamp 1621261055
transform 1 0 14112 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_143
timestamp 1621261055
transform 1 0 14880 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_151
timestamp 1621261055
transform 1 0 15648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_159
timestamp 1621261055
transform 1 0 16416 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_163
timestamp 1621261055
transform 1 0 16800 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_166
timestamp 1621261055
transform 1 0 17088 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_174
timestamp 1621261055
transform 1 0 17856 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_182
timestamp 1621261055
transform 1 0 18624 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_190
timestamp 1621261055
transform 1 0 19392 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_198
timestamp 1621261055
transform 1 0 20160 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _036_
timestamp 1621261055
transform 1 0 20640 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_608
timestamp 1621261055
transform 1 0 22272 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_41_202
timestamp 1621261055
transform 1 0 20544 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_206
timestamp 1621261055
transform 1 0 20928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_214
timestamp 1621261055
transform 1 0 21696 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_218
timestamp 1621261055
transform 1 0 22080 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_221
timestamp 1621261055
transform 1 0 22368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_229
timestamp 1621261055
transform 1 0 23136 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_237
timestamp 1621261055
transform 1 0 23904 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_245
timestamp 1621261055
transform 1 0 24672 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_253
timestamp 1621261055
transform 1 0 25440 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_261
timestamp 1621261055
transform 1 0 26208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_609
timestamp 1621261055
transform 1 0 27552 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_269
timestamp 1621261055
transform 1 0 26976 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_273
timestamp 1621261055
transform 1 0 27360 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_276
timestamp 1621261055
transform 1 0 27648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_284
timestamp 1621261055
transform 1 0 28416 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_292
timestamp 1621261055
transform 1 0 29184 0 1 29970
box -38 -49 806 715
use INVX1  INVX1
timestamp 1623610208
transform 1 0 29952 0 1 29970
box 0 -48 576 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_610
timestamp 1621261055
transform 1 0 32832 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_306
timestamp 1621261055
transform 1 0 30528 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_314
timestamp 1621261055
transform 1 0 31296 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_322
timestamp 1621261055
transform 1 0 32064 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_331
timestamp 1621261055
transform 1 0 32928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_339
timestamp 1621261055
transform 1 0 33696 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_347
timestamp 1621261055
transform 1 0 34464 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_355
timestamp 1621261055
transform 1 0 35232 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_363
timestamp 1621261055
transform 1 0 36000 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_611
timestamp 1621261055
transform 1 0 38112 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_371
timestamp 1621261055
transform 1 0 36768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_379
timestamp 1621261055
transform 1 0 37536 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_383
timestamp 1621261055
transform 1 0 37920 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_386
timestamp 1621261055
transform 1 0 38208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_394
timestamp 1621261055
transform 1 0 38976 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_402
timestamp 1621261055
transform 1 0 39744 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_410
timestamp 1621261055
transform 1 0 40512 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_418
timestamp 1621261055
transform 1 0 41280 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_426
timestamp 1621261055
transform 1 0 42048 0 1 29970
box -38 -49 806 715
use OAI22X1  OAI22X1
timestamp 1623610208
transform 1 0 44352 0 1 29970
box 0 -48 1440 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_612
timestamp 1621261055
transform 1 0 43392 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_434
timestamp 1621261055
transform 1 0 42816 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_438
timestamp 1621261055
transform 1 0 43200 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_441
timestamp 1621261055
transform 1 0 43488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_41_449
timestamp 1621261055
transform 1 0 44256 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _156_
timestamp 1621261055
transform 1 0 46560 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_613
timestamp 1621261055
transform 1 0 48672 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_465
timestamp 1621261055
transform 1 0 45792 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_476
timestamp 1621261055
transform 1 0 46848 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_484
timestamp 1621261055
transform 1 0 47616 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_492
timestamp 1621261055
transform 1 0 48384 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_41_494
timestamp 1621261055
transform 1 0 48576 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_496
timestamp 1621261055
transform 1 0 48768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_504
timestamp 1621261055
transform 1 0 49536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_512
timestamp 1621261055
transform 1 0 50304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_520
timestamp 1621261055
transform 1 0 51072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_528
timestamp 1621261055
transform 1 0 51840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_614
timestamp 1621261055
transform 1 0 53952 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_536
timestamp 1621261055
transform 1 0 52608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_544
timestamp 1621261055
transform 1 0 53376 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_548
timestamp 1621261055
transform 1 0 53760 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_551
timestamp 1621261055
transform 1 0 54048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_559
timestamp 1621261055
transform 1 0 54816 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_567
timestamp 1621261055
transform 1 0 55584 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_575
timestamp 1621261055
transform 1 0 56352 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_583
timestamp 1621261055
transform 1 0 57120 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_591
timestamp 1621261055
transform 1 0 57888 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_83
timestamp 1621261055
transform -1 0 58848 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_595
timestamp 1621261055
transform 1 0 58272 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_84
timestamp 1621261055
transform 1 0 1152 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_615
timestamp 1621261055
transform 1 0 3840 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_4
timestamp 1621261055
transform 1 0 1536 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_12
timestamp 1621261055
transform 1 0 2304 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_20
timestamp 1621261055
transform 1 0 3072 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_29
timestamp 1621261055
transform 1 0 3936 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_37
timestamp 1621261055
transform 1 0 4704 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_45
timestamp 1621261055
transform 1 0 5472 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_53
timestamp 1621261055
transform 1 0 6240 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_61
timestamp 1621261055
transform 1 0 7008 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_616
timestamp 1621261055
transform 1 0 9120 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_69
timestamp 1621261055
transform 1 0 7776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_77
timestamp 1621261055
transform 1 0 8544 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_81
timestamp 1621261055
transform 1 0 8928 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_84
timestamp 1621261055
transform 1 0 9216 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_92
timestamp 1621261055
transform 1 0 9984 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_100
timestamp 1621261055
transform 1 0 10752 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_108
timestamp 1621261055
transform 1 0 11520 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_116
timestamp 1621261055
transform 1 0 12288 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_124
timestamp 1621261055
transform 1 0 13056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_132
timestamp 1621261055
transform 1 0 13824 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_617
timestamp 1621261055
transform 1 0 14400 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_136
timestamp 1621261055
transform 1 0 14208 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_139
timestamp 1621261055
transform 1 0 14496 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_147
timestamp 1621261055
transform 1 0 15264 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_155
timestamp 1621261055
transform 1 0 16032 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_163
timestamp 1621261055
transform 1 0 16800 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_618
timestamp 1621261055
transform 1 0 19680 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_171
timestamp 1621261055
transform 1 0 17568 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_179
timestamp 1621261055
transform 1 0 18336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_187
timestamp 1621261055
transform 1 0 19104 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_191
timestamp 1621261055
transform 1 0 19488 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_194
timestamp 1621261055
transform 1 0 19776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _015_
timestamp 1621261055
transform 1 0 23040 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_202
timestamp 1621261055
transform 1 0 20544 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_210
timestamp 1621261055
transform 1 0 21312 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_218
timestamp 1621261055
transform 1 0 22080 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_226
timestamp 1621261055
transform 1 0 22848 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_231
timestamp 1621261055
transform 1 0 23328 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_619
timestamp 1621261055
transform 1 0 24960 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_239
timestamp 1621261055
transform 1 0 24096 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_42_247
timestamp 1621261055
transform 1 0 24864 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_249
timestamp 1621261055
transform 1 0 25056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_257
timestamp 1621261055
transform 1 0 25824 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_265
timestamp 1621261055
transform 1 0 26592 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_273
timestamp 1621261055
transform 1 0 27360 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_281
timestamp 1621261055
transform 1 0 28128 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_289
timestamp 1621261055
transform 1 0 28896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_297
timestamp 1621261055
transform 1 0 29664 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_620
timestamp 1621261055
transform 1 0 30240 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_301
timestamp 1621261055
transform 1 0 30048 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_304
timestamp 1621261055
transform 1 0 30336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_312
timestamp 1621261055
transform 1 0 31104 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_320
timestamp 1621261055
transform 1 0 31872 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_328
timestamp 1621261055
transform 1 0 32640 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_621
timestamp 1621261055
transform 1 0 35520 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_336
timestamp 1621261055
transform 1 0 33408 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_344
timestamp 1621261055
transform 1 0 34176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_352
timestamp 1621261055
transform 1 0 34944 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_356
timestamp 1621261055
transform 1 0 35328 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_359
timestamp 1621261055
transform 1 0 35616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_367
timestamp 1621261055
transform 1 0 36384 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_375
timestamp 1621261055
transform 1 0 37152 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_383
timestamp 1621261055
transform 1 0 37920 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_391
timestamp 1621261055
transform 1 0 38688 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_622
timestamp 1621261055
transform 1 0 40800 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_399
timestamp 1621261055
transform 1 0 39456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_407
timestamp 1621261055
transform 1 0 40224 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_411
timestamp 1621261055
transform 1 0 40608 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_414
timestamp 1621261055
transform 1 0 40896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_422
timestamp 1621261055
transform 1 0 41664 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_430
timestamp 1621261055
transform 1 0 42432 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_438
timestamp 1621261055
transform 1 0 43200 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_446
timestamp 1621261055
transform 1 0 43968 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_454
timestamp 1621261055
transform 1 0 44736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_462
timestamp 1621261055
transform 1 0 45504 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_623
timestamp 1621261055
transform 1 0 46080 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_466
timestamp 1621261055
transform 1 0 45888 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_469
timestamp 1621261055
transform 1 0 46176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_477
timestamp 1621261055
transform 1 0 46944 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_485
timestamp 1621261055
transform 1 0 47712 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_493
timestamp 1621261055
transform 1 0 48480 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_624
timestamp 1621261055
transform 1 0 51360 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_501
timestamp 1621261055
transform 1 0 49248 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_509
timestamp 1621261055
transform 1 0 50016 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_517
timestamp 1621261055
transform 1 0 50784 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_521
timestamp 1621261055
transform 1 0 51168 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_524
timestamp 1621261055
transform 1 0 51456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_532
timestamp 1621261055
transform 1 0 52224 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_540
timestamp 1621261055
transform 1 0 52992 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_548
timestamp 1621261055
transform 1 0 53760 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_556
timestamp 1621261055
transform 1 0 54528 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_625
timestamp 1621261055
transform 1 0 56640 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_564
timestamp 1621261055
transform 1 0 55296 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_572
timestamp 1621261055
transform 1 0 56064 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_576
timestamp 1621261055
transform 1 0 56448 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_579
timestamp 1621261055
transform 1 0 56736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_587
timestamp 1621261055
transform 1 0 57504 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_85
timestamp 1621261055
transform -1 0 58848 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_595
timestamp 1621261055
transform 1 0 58272 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_86
timestamp 1621261055
transform 1 0 1152 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_43_4
timestamp 1621261055
transform 1 0 1536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_12
timestamp 1621261055
transform 1 0 2304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_20
timestamp 1621261055
transform 1 0 3072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_28
timestamp 1621261055
transform 1 0 3840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_626
timestamp 1621261055
transform 1 0 6432 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_36
timestamp 1621261055
transform 1 0 4608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_44
timestamp 1621261055
transform 1 0 5376 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_52
timestamp 1621261055
transform 1 0 6144 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_54
timestamp 1621261055
transform 1 0 6336 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_56
timestamp 1621261055
transform 1 0 6528 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_64
timestamp 1621261055
transform 1 0 7296 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_72
timestamp 1621261055
transform 1 0 8064 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_80
timestamp 1621261055
transform 1 0 8832 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_88
timestamp 1621261055
transform 1 0 9600 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_96
timestamp 1621261055
transform 1 0 10368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_627
timestamp 1621261055
transform 1 0 11712 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_104
timestamp 1621261055
transform 1 0 11136 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_108
timestamp 1621261055
transform 1 0 11520 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_111
timestamp 1621261055
transform 1 0 11808 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_119
timestamp 1621261055
transform 1 0 12576 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_127
timestamp 1621261055
transform 1 0 13344 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_628
timestamp 1621261055
transform 1 0 16992 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_135
timestamp 1621261055
transform 1 0 14112 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_143
timestamp 1621261055
transform 1 0 14880 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_151
timestamp 1621261055
transform 1 0 15648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_159
timestamp 1621261055
transform 1 0 16416 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_163
timestamp 1621261055
transform 1 0 16800 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_166
timestamp 1621261055
transform 1 0 17088 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_174
timestamp 1621261055
transform 1 0 17856 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_182
timestamp 1621261055
transform 1 0 18624 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_190
timestamp 1621261055
transform 1 0 19392 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_198
timestamp 1621261055
transform 1 0 20160 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_629
timestamp 1621261055
transform 1 0 22272 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_206
timestamp 1621261055
transform 1 0 20928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_214
timestamp 1621261055
transform 1 0 21696 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_218
timestamp 1621261055
transform 1 0 22080 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_221
timestamp 1621261055
transform 1 0 22368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_229
timestamp 1621261055
transform 1 0 23136 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _141_
timestamp 1621261055
transform 1 0 26304 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_43_237
timestamp 1621261055
transform 1 0 23904 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_245
timestamp 1621261055
transform 1 0 24672 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_253
timestamp 1621261055
transform 1 0 25440 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_43_261
timestamp 1621261055
transform 1 0 26208 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_630
timestamp 1621261055
transform 1 0 27552 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_265
timestamp 1621261055
transform 1 0 26592 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_273
timestamp 1621261055
transform 1 0 27360 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_276
timestamp 1621261055
transform 1 0 27648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_284
timestamp 1621261055
transform 1 0 28416 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_292
timestamp 1621261055
transform 1 0 29184 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_631
timestamp 1621261055
transform 1 0 32832 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_300
timestamp 1621261055
transform 1 0 29952 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_308
timestamp 1621261055
transform 1 0 30720 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_316
timestamp 1621261055
transform 1 0 31488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_324
timestamp 1621261055
transform 1 0 32256 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_328
timestamp 1621261055
transform 1 0 32640 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_331
timestamp 1621261055
transform 1 0 32928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_339
timestamp 1621261055
transform 1 0 33696 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_347
timestamp 1621261055
transform 1 0 34464 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_355
timestamp 1621261055
transform 1 0 35232 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_363
timestamp 1621261055
transform 1 0 36000 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_632
timestamp 1621261055
transform 1 0 38112 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_371
timestamp 1621261055
transform 1 0 36768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_379
timestamp 1621261055
transform 1 0 37536 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_383
timestamp 1621261055
transform 1 0 37920 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_386
timestamp 1621261055
transform 1 0 38208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_394
timestamp 1621261055
transform 1 0 38976 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_402
timestamp 1621261055
transform 1 0 39744 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_410
timestamp 1621261055
transform 1 0 40512 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_418
timestamp 1621261055
transform 1 0 41280 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_426
timestamp 1621261055
transform 1 0 42048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_633
timestamp 1621261055
transform 1 0 43392 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_434
timestamp 1621261055
transform 1 0 42816 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_438
timestamp 1621261055
transform 1 0 43200 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_441
timestamp 1621261055
transform 1 0 43488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_449
timestamp 1621261055
transform 1 0 44256 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_457
timestamp 1621261055
transform 1 0 45024 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_634
timestamp 1621261055
transform 1 0 48672 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_465
timestamp 1621261055
transform 1 0 45792 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_473
timestamp 1621261055
transform 1 0 46560 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_481
timestamp 1621261055
transform 1 0 47328 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_489
timestamp 1621261055
transform 1 0 48096 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_493
timestamp 1621261055
transform 1 0 48480 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_496
timestamp 1621261055
transform 1 0 48768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_504
timestamp 1621261055
transform 1 0 49536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_512
timestamp 1621261055
transform 1 0 50304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_520
timestamp 1621261055
transform 1 0 51072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_528
timestamp 1621261055
transform 1 0 51840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_635
timestamp 1621261055
transform 1 0 53952 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_536
timestamp 1621261055
transform 1 0 52608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_544
timestamp 1621261055
transform 1 0 53376 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_548
timestamp 1621261055
transform 1 0 53760 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_551
timestamp 1621261055
transform 1 0 54048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_559
timestamp 1621261055
transform 1 0 54816 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _171_
timestamp 1621261055
transform 1 0 57120 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_43_567
timestamp 1621261055
transform 1 0 55584 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_575
timestamp 1621261055
transform 1 0 56352 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_586
timestamp 1621261055
transform 1 0 57408 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_594
timestamp 1621261055
transform 1 0 58176 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_87
timestamp 1621261055
transform -1 0 58848 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_43_596
timestamp 1621261055
transform 1 0 58368 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_88
timestamp 1621261055
transform 1 0 1152 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_636
timestamp 1621261055
transform 1 0 3840 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_4
timestamp 1621261055
transform 1 0 1536 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_12
timestamp 1621261055
transform 1 0 2304 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_20
timestamp 1621261055
transform 1 0 3072 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_29
timestamp 1621261055
transform 1 0 3936 0 -1 32634
box -38 -49 806 715
use MUX2X1  MUX2X1
timestamp 1623610208
transform 1 0 5856 0 -1 32634
box 0 -48 1728 714
use sky130_fd_sc_ls__decap_8  FILLER_44_37
timestamp 1621261055
transform 1 0 4704 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_45
timestamp 1621261055
transform 1 0 5472 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_637
timestamp 1621261055
transform 1 0 9120 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_67
timestamp 1621261055
transform 1 0 7584 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_75
timestamp 1621261055
transform 1 0 8352 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_84
timestamp 1621261055
transform 1 0 9216 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_92
timestamp 1621261055
transform 1 0 9984 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _143_
timestamp 1621261055
transform 1 0 12864 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_44_100
timestamp 1621261055
transform 1 0 10752 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_108
timestamp 1621261055
transform 1 0 11520 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_116
timestamp 1621261055
transform 1 0 12288 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_120
timestamp 1621261055
transform 1 0 12672 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_125
timestamp 1621261055
transform 1 0 13152 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_638
timestamp 1621261055
transform 1 0 14400 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_133
timestamp 1621261055
transform 1 0 13920 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_44_137
timestamp 1621261055
transform 1 0 14304 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_139
timestamp 1621261055
transform 1 0 14496 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_147
timestamp 1621261055
transform 1 0 15264 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_155
timestamp 1621261055
transform 1 0 16032 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_163
timestamp 1621261055
transform 1 0 16800 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_639
timestamp 1621261055
transform 1 0 19680 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_171
timestamp 1621261055
transform 1 0 17568 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_179
timestamp 1621261055
transform 1 0 18336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_187
timestamp 1621261055
transform 1 0 19104 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_191
timestamp 1621261055
transform 1 0 19488 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_194
timestamp 1621261055
transform 1 0 19776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_202
timestamp 1621261055
transform 1 0 20544 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_210
timestamp 1621261055
transform 1 0 21312 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_218
timestamp 1621261055
transform 1 0 22080 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_226
timestamp 1621261055
transform 1 0 22848 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_640
timestamp 1621261055
transform 1 0 24960 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_234
timestamp 1621261055
transform 1 0 23616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_242
timestamp 1621261055
transform 1 0 24384 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_246
timestamp 1621261055
transform 1 0 24768 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_249
timestamp 1621261055
transform 1 0 25056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_257
timestamp 1621261055
transform 1 0 25824 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_265
timestamp 1621261055
transform 1 0 26592 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_273
timestamp 1621261055
transform 1 0 27360 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_281
timestamp 1621261055
transform 1 0 28128 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_289
timestamp 1621261055
transform 1 0 28896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_297
timestamp 1621261055
transform 1 0 29664 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_641
timestamp 1621261055
transform 1 0 30240 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_301
timestamp 1621261055
transform 1 0 30048 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_304
timestamp 1621261055
transform 1 0 30336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_312
timestamp 1621261055
transform 1 0 31104 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_320
timestamp 1621261055
transform 1 0 31872 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_328
timestamp 1621261055
transform 1 0 32640 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_642
timestamp 1621261055
transform 1 0 35520 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_336
timestamp 1621261055
transform 1 0 33408 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_344
timestamp 1621261055
transform 1 0 34176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_352
timestamp 1621261055
transform 1 0 34944 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_356
timestamp 1621261055
transform 1 0 35328 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_359
timestamp 1621261055
transform 1 0 35616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_367
timestamp 1621261055
transform 1 0 36384 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_375
timestamp 1621261055
transform 1 0 37152 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_383
timestamp 1621261055
transform 1 0 37920 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_391
timestamp 1621261055
transform 1 0 38688 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_643
timestamp 1621261055
transform 1 0 40800 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_399
timestamp 1621261055
transform 1 0 39456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_407
timestamp 1621261055
transform 1 0 40224 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_411
timestamp 1621261055
transform 1 0 40608 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_414
timestamp 1621261055
transform 1 0 40896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_422
timestamp 1621261055
transform 1 0 41664 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_430
timestamp 1621261055
transform 1 0 42432 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_438
timestamp 1621261055
transform 1 0 43200 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_446
timestamp 1621261055
transform 1 0 43968 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_454
timestamp 1621261055
transform 1 0 44736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_462
timestamp 1621261055
transform 1 0 45504 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_644
timestamp 1621261055
transform 1 0 46080 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_466
timestamp 1621261055
transform 1 0 45888 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_469
timestamp 1621261055
transform 1 0 46176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_477
timestamp 1621261055
transform 1 0 46944 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_485
timestamp 1621261055
transform 1 0 47712 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_493
timestamp 1621261055
transform 1 0 48480 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_645
timestamp 1621261055
transform 1 0 51360 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_501
timestamp 1621261055
transform 1 0 49248 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_509
timestamp 1621261055
transform 1 0 50016 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_517
timestamp 1621261055
transform 1 0 50784 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_521
timestamp 1621261055
transform 1 0 51168 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_524
timestamp 1621261055
transform 1 0 51456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_532
timestamp 1621261055
transform 1 0 52224 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_540
timestamp 1621261055
transform 1 0 52992 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_548
timestamp 1621261055
transform 1 0 53760 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_556
timestamp 1621261055
transform 1 0 54528 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_646
timestamp 1621261055
transform 1 0 56640 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_564
timestamp 1621261055
transform 1 0 55296 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_572
timestamp 1621261055
transform 1 0 56064 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_576
timestamp 1621261055
transform 1 0 56448 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_579
timestamp 1621261055
transform 1 0 56736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_587
timestamp 1621261055
transform 1 0 57504 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_89
timestamp 1621261055
transform -1 0 58848 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_595
timestamp 1621261055
transform 1 0 58272 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_90
timestamp 1621261055
transform 1 0 1152 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_4
timestamp 1621261055
transform 1 0 1536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_12
timestamp 1621261055
transform 1 0 2304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_20
timestamp 1621261055
transform 1 0 3072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_28
timestamp 1621261055
transform 1 0 3840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_647
timestamp 1621261055
transform 1 0 6432 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_36
timestamp 1621261055
transform 1 0 4608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_44
timestamp 1621261055
transform 1 0 5376 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_52
timestamp 1621261055
transform 1 0 6144 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_54
timestamp 1621261055
transform 1 0 6336 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_56
timestamp 1621261055
transform 1 0 6528 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_64
timestamp 1621261055
transform 1 0 7296 0 1 32634
box -38 -49 806 715
use AOI21X1  AOI21X1
timestamp 1623610208
transform 1 0 8160 0 1 32634
box 0 -48 1152 714
use sky130_fd_sc_ls__fill_1  FILLER_45_72
timestamp 1621261055
transform 1 0 8064 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_85
timestamp 1621261055
transform 1 0 9312 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_93
timestamp 1621261055
transform 1 0 10080 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_648
timestamp 1621261055
transform 1 0 11712 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_101
timestamp 1621261055
transform 1 0 10848 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_45_109
timestamp 1621261055
transform 1 0 11616 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_111
timestamp 1621261055
transform 1 0 11808 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_119
timestamp 1621261055
transform 1 0 12576 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_127
timestamp 1621261055
transform 1 0 13344 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_649
timestamp 1621261055
transform 1 0 16992 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_135
timestamp 1621261055
transform 1 0 14112 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_143
timestamp 1621261055
transform 1 0 14880 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_151
timestamp 1621261055
transform 1 0 15648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_159
timestamp 1621261055
transform 1 0 16416 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_163
timestamp 1621261055
transform 1 0 16800 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_166
timestamp 1621261055
transform 1 0 17088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_174
timestamp 1621261055
transform 1 0 17856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_182
timestamp 1621261055
transform 1 0 18624 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_190
timestamp 1621261055
transform 1 0 19392 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_198
timestamp 1621261055
transform 1 0 20160 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_650
timestamp 1621261055
transform 1 0 22272 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_206
timestamp 1621261055
transform 1 0 20928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_214
timestamp 1621261055
transform 1 0 21696 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_218
timestamp 1621261055
transform 1 0 22080 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_221
timestamp 1621261055
transform 1 0 22368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_229
timestamp 1621261055
transform 1 0 23136 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_237
timestamp 1621261055
transform 1 0 23904 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_245
timestamp 1621261055
transform 1 0 24672 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_253
timestamp 1621261055
transform 1 0 25440 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_261
timestamp 1621261055
transform 1 0 26208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_651
timestamp 1621261055
transform 1 0 27552 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_269
timestamp 1621261055
transform 1 0 26976 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_273
timestamp 1621261055
transform 1 0 27360 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_276
timestamp 1621261055
transform 1 0 27648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_284
timestamp 1621261055
transform 1 0 28416 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_292
timestamp 1621261055
transform 1 0 29184 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_652
timestamp 1621261055
transform 1 0 32832 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_300
timestamp 1621261055
transform 1 0 29952 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_308
timestamp 1621261055
transform 1 0 30720 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_316
timestamp 1621261055
transform 1 0 31488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_324
timestamp 1621261055
transform 1 0 32256 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_328
timestamp 1621261055
transform 1 0 32640 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_331
timestamp 1621261055
transform 1 0 32928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_339
timestamp 1621261055
transform 1 0 33696 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_347
timestamp 1621261055
transform 1 0 34464 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_355
timestamp 1621261055
transform 1 0 35232 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_363
timestamp 1621261055
transform 1 0 36000 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_653
timestamp 1621261055
transform 1 0 38112 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_371
timestamp 1621261055
transform 1 0 36768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_379
timestamp 1621261055
transform 1 0 37536 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_383
timestamp 1621261055
transform 1 0 37920 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_386
timestamp 1621261055
transform 1 0 38208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_394
timestamp 1621261055
transform 1 0 38976 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_402
timestamp 1621261055
transform 1 0 39744 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_410
timestamp 1621261055
transform 1 0 40512 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_418
timestamp 1621261055
transform 1 0 41280 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_426
timestamp 1621261055
transform 1 0 42048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_654
timestamp 1621261055
transform 1 0 43392 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_434
timestamp 1621261055
transform 1 0 42816 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_438
timestamp 1621261055
transform 1 0 43200 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_441
timestamp 1621261055
transform 1 0 43488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_449
timestamp 1621261055
transform 1 0 44256 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_457
timestamp 1621261055
transform 1 0 45024 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_655
timestamp 1621261055
transform 1 0 48672 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_465
timestamp 1621261055
transform 1 0 45792 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_473
timestamp 1621261055
transform 1 0 46560 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_481
timestamp 1621261055
transform 1 0 47328 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_489
timestamp 1621261055
transform 1 0 48096 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_493
timestamp 1621261055
transform 1 0 48480 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_496
timestamp 1621261055
transform 1 0 48768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_504
timestamp 1621261055
transform 1 0 49536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_512
timestamp 1621261055
transform 1 0 50304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_520
timestamp 1621261055
transform 1 0 51072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_528
timestamp 1621261055
transform 1 0 51840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_656
timestamp 1621261055
transform 1 0 53952 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_536
timestamp 1621261055
transform 1 0 52608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_544
timestamp 1621261055
transform 1 0 53376 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_548
timestamp 1621261055
transform 1 0 53760 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_551
timestamp 1621261055
transform 1 0 54048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_559
timestamp 1621261055
transform 1 0 54816 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _034_
timestamp 1621261055
transform 1 0 57120 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_45_567
timestamp 1621261055
transform 1 0 55584 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_575
timestamp 1621261055
transform 1 0 56352 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_586
timestamp 1621261055
transform 1 0 57408 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_594
timestamp 1621261055
transform 1 0 58176 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_91
timestamp 1621261055
transform -1 0 58848 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_45_596
timestamp 1621261055
transform 1 0 58368 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_4
timestamp 1621261055
transform 1 0 1536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_4
timestamp 1621261055
transform 1 0 1536 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_94
timestamp 1621261055
transform 1 0 1152 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_92
timestamp 1621261055
transform 1 0 1152 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_12
timestamp 1621261055
transform 1 0 2304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_12
timestamp 1621261055
transform 1 0 2304 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_20
timestamp 1621261055
transform 1 0 3072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_20
timestamp 1621261055
transform 1 0 3072 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_28
timestamp 1621261055
transform 1 0 3840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_29
timestamp 1621261055
transform 1 0 3936 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_657
timestamp 1621261055
transform 1 0 3840 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_36
timestamp 1621261055
transform 1 0 4608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_37
timestamp 1621261055
transform 1 0 4704 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_44
timestamp 1621261055
transform 1 0 5376 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_45
timestamp 1621261055
transform 1 0 5472 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_56
timestamp 1621261055
transform 1 0 6528 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_54
timestamp 1621261055
transform 1 0 6336 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_52
timestamp 1621261055
transform 1 0 6144 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_53
timestamp 1621261055
transform 1 0 6240 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_668
timestamp 1621261055
transform 1 0 6432 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_64
timestamp 1621261055
transform 1 0 7296 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_61
timestamp 1621261055
transform 1 0 7008 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_72
timestamp 1621261055
transform 1 0 8064 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_69
timestamp 1621261055
transform 1 0 7776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_80
timestamp 1621261055
transform 1 0 8832 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_81
timestamp 1621261055
transform 1 0 8928 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_77
timestamp 1621261055
transform 1 0 8544 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_658
timestamp 1621261055
transform 1 0 9120 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_88
timestamp 1621261055
transform 1 0 9600 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_92
timestamp 1621261055
transform 1 0 9984 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_84
timestamp 1621261055
transform 1 0 9216 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_96
timestamp 1621261055
transform 1 0 10368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_104
timestamp 1621261055
transform 1 0 11136 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_100
timestamp 1621261055
transform 1 0 10752 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_111
timestamp 1621261055
transform 1 0 11808 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_108
timestamp 1621261055
transform 1 0 11520 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_116
timestamp 1621261055
transform 1 0 12288 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_108
timestamp 1621261055
transform 1 0 11520 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_669
timestamp 1621261055
transform 1 0 11712 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_119
timestamp 1621261055
transform 1 0 12576 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_124
timestamp 1621261055
transform 1 0 13056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_127
timestamp 1621261055
transform 1 0 13344 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_132
timestamp 1621261055
transform 1 0 13824 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_135
timestamp 1621261055
transform 1 0 14112 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_139
timestamp 1621261055
transform 1 0 14496 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_136
timestamp 1621261055
transform 1 0 14208 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_659
timestamp 1621261055
transform 1 0 14400 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_143
timestamp 1621261055
transform 1 0 14880 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_147
timestamp 1621261055
transform 1 0 15264 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_151
timestamp 1621261055
transform 1 0 15648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_155
timestamp 1621261055
transform 1 0 16032 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_163
timestamp 1621261055
transform 1 0 16800 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_159
timestamp 1621261055
transform 1 0 16416 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_163
timestamp 1621261055
transform 1 0 16800 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_670
timestamp 1621261055
transform 1 0 16992 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_166
timestamp 1621261055
transform 1 0 17088 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_171
timestamp 1621261055
transform 1 0 17568 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_182
timestamp 1621261055
transform 1 0 18624 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_174
timestamp 1621261055
transform 1 0 17856 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_179
timestamp 1621261055
transform 1 0 18336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_190
timestamp 1621261055
transform 1 0 19392 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_191
timestamp 1621261055
transform 1 0 19488 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_187
timestamp 1621261055
transform 1 0 19104 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_198
timestamp 1621261055
transform 1 0 20160 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_194
timestamp 1621261055
transform 1 0 19776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_660
timestamp 1621261055
transform 1 0 19680 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_206
timestamp 1621261055
transform 1 0 20928 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_202
timestamp 1621261055
transform 1 0 20544 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_211
timestamp 1621261055
transform 1 0 21408 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_210
timestamp 1621261055
transform 1 0 21312 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _121_
timestamp 1621261055
transform 1 0 21120 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_221
timestamp 1621261055
transform 1 0 22368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_219
timestamp 1621261055
transform 1 0 22176 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_218
timestamp 1621261055
transform 1 0 22080 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_671
timestamp 1621261055
transform 1 0 22272 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_229
timestamp 1621261055
transform 1 0 23136 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_226
timestamp 1621261055
transform 1 0 22848 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_237
timestamp 1621261055
transform 1 0 23904 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_234
timestamp 1621261055
transform 1 0 23616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_245
timestamp 1621261055
transform 1 0 24672 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_246
timestamp 1621261055
transform 1 0 24768 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_242
timestamp 1621261055
transform 1 0 24384 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_661
timestamp 1621261055
transform 1 0 24960 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_253
timestamp 1621261055
transform 1 0 25440 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_257
timestamp 1621261055
transform 1 0 25824 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_249
timestamp 1621261055
transform 1 0 25056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_261
timestamp 1621261055
transform 1 0 26208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_269
timestamp 1621261055
transform 1 0 26976 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_265
timestamp 1621261055
transform 1 0 26592 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_276
timestamp 1621261055
transform 1 0 27648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_273
timestamp 1621261055
transform 1 0 27360 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_281
timestamp 1621261055
transform 1 0 28128 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_273
timestamp 1621261055
transform 1 0 27360 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_672
timestamp 1621261055
transform 1 0 27552 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_284
timestamp 1621261055
transform 1 0 28416 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_289
timestamp 1621261055
transform 1 0 28896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_292
timestamp 1621261055
transform 1 0 29184 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_297
timestamp 1621261055
transform 1 0 29664 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_300
timestamp 1621261055
transform 1 0 29952 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_304
timestamp 1621261055
transform 1 0 30336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_301
timestamp 1621261055
transform 1 0 30048 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_662
timestamp 1621261055
transform 1 0 30240 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_308
timestamp 1621261055
transform 1 0 30720 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_312
timestamp 1621261055
transform 1 0 31104 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_316
timestamp 1621261055
transform 1 0 31488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_320
timestamp 1621261055
transform 1 0 31872 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_328
timestamp 1621261055
transform 1 0 32640 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_324
timestamp 1621261055
transform 1 0 32256 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_328
timestamp 1621261055
transform 1 0 32640 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_673
timestamp 1621261055
transform 1 0 32832 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_331
timestamp 1621261055
transform 1 0 32928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_336
timestamp 1621261055
transform 1 0 33408 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_347
timestamp 1621261055
transform 1 0 34464 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_339
timestamp 1621261055
transform 1 0 33696 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_344
timestamp 1621261055
transform 1 0 34176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_355
timestamp 1621261055
transform 1 0 35232 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_356
timestamp 1621261055
transform 1 0 35328 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_352
timestamp 1621261055
transform 1 0 34944 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_47_363
timestamp 1621261055
transform 1 0 36000 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_359
timestamp 1621261055
transform 1 0 35616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_663
timestamp 1621261055
transform 1 0 35520 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_371
timestamp 1621261055
transform 1 0 36768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_367
timestamp 1621261055
transform 1 0 36384 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_367
timestamp 1621261055
transform 1 0 36384 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _176_
timestamp 1621261055
transform 1 0 36480 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_47_379
timestamp 1621261055
transform 1 0 37536 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_375
timestamp 1621261055
transform 1 0 37152 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_386
timestamp 1621261055
transform 1 0 38208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_383
timestamp 1621261055
transform 1 0 37920 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_383
timestamp 1621261055
transform 1 0 37920 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_674
timestamp 1621261055
transform 1 0 38112 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_394
timestamp 1621261055
transform 1 0 38976 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_391
timestamp 1621261055
transform 1 0 38688 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_402
timestamp 1621261055
transform 1 0 39744 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_399
timestamp 1621261055
transform 1 0 39456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_410
timestamp 1621261055
transform 1 0 40512 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_411
timestamp 1621261055
transform 1 0 40608 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_407
timestamp 1621261055
transform 1 0 40224 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_664
timestamp 1621261055
transform 1 0 40800 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_418
timestamp 1621261055
transform 1 0 41280 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_422
timestamp 1621261055
transform 1 0 41664 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_414
timestamp 1621261055
transform 1 0 40896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_426
timestamp 1621261055
transform 1 0 42048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_434
timestamp 1621261055
transform 1 0 42816 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_430
timestamp 1621261055
transform 1 0 42432 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_441
timestamp 1621261055
transform 1 0 43488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_438
timestamp 1621261055
transform 1 0 43200 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_446
timestamp 1621261055
transform 1 0 43968 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_438
timestamp 1621261055
transform 1 0 43200 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_675
timestamp 1621261055
transform 1 0 43392 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_449
timestamp 1621261055
transform 1 0 44256 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_454
timestamp 1621261055
transform 1 0 44736 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_457
timestamp 1621261055
transform 1 0 45024 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_460
timestamp 1621261055
transform 1 0 45312 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_458
timestamp 1621261055
transform 1 0 45120 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _129_
timestamp 1621261055
transform 1 0 45408 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_465
timestamp 1621261055
transform 1 0 45792 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_469
timestamp 1621261055
transform 1 0 46176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_464
timestamp 1621261055
transform 1 0 45696 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_665
timestamp 1621261055
transform 1 0 46080 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_473
timestamp 1621261055
transform 1 0 46560 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_477
timestamp 1621261055
transform 1 0 46944 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_481
timestamp 1621261055
transform 1 0 47328 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_485
timestamp 1621261055
transform 1 0 47712 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_493
timestamp 1621261055
transform 1 0 48480 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_489
timestamp 1621261055
transform 1 0 48096 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_493
timestamp 1621261055
transform 1 0 48480 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_676
timestamp 1621261055
transform 1 0 48672 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_496
timestamp 1621261055
transform 1 0 48768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_501
timestamp 1621261055
transform 1 0 49248 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_512
timestamp 1621261055
transform 1 0 50304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_504
timestamp 1621261055
transform 1 0 49536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_509
timestamp 1621261055
transform 1 0 50016 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_520
timestamp 1621261055
transform 1 0 51072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_521
timestamp 1621261055
transform 1 0 51168 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_517
timestamp 1621261055
transform 1 0 50784 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_528
timestamp 1621261055
transform 1 0 51840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_524
timestamp 1621261055
transform 1 0 51456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_666
timestamp 1621261055
transform 1 0 51360 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_536
timestamp 1621261055
transform 1 0 52608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_534
timestamp 1621261055
transform 1 0 52416 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_532
timestamp 1621261055
transform 1 0 52224 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_139
timestamp 1621261055
transform -1 0 52704 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_544
timestamp 1621261055
transform 1 0 53376 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_540
timestamp 1621261055
transform 1 0 52992 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _104_
timestamp 1621261055
transform -1 0 52992 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_551
timestamp 1621261055
transform 1 0 54048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_548
timestamp 1621261055
transform 1 0 53760 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_548
timestamp 1621261055
transform 1 0 53760 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_677
timestamp 1621261055
transform 1 0 53952 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_559
timestamp 1621261055
transform 1 0 54816 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_556
timestamp 1621261055
transform 1 0 54528 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_567
timestamp 1621261055
transform 1 0 55584 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_564
timestamp 1621261055
transform 1 0 55296 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_575
timestamp 1621261055
transform 1 0 56352 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_576
timestamp 1621261055
transform 1 0 56448 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_572
timestamp 1621261055
transform 1 0 56064 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_667
timestamp 1621261055
transform 1 0 56640 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_583
timestamp 1621261055
transform 1 0 57120 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_587
timestamp 1621261055
transform 1 0 57504 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_579
timestamp 1621261055
transform 1 0 56736 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_591
timestamp 1621261055
transform 1 0 57888 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_93
timestamp 1621261055
transform -1 0 58848 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_95
timestamp 1621261055
transform -1 0 58848 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_595
timestamp 1621261055
transform 1 0 58272 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_595
timestamp 1621261055
transform 1 0 58272 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _024_
timestamp 1621261055
transform 1 0 4320 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_96
timestamp 1621261055
transform 1 0 1152 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_678
timestamp 1621261055
transform 1 0 3840 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_4
timestamp 1621261055
transform 1 0 1536 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_12
timestamp 1621261055
transform 1 0 2304 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_20
timestamp 1621261055
transform 1 0 3072 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_29
timestamp 1621261055
transform 1 0 3936 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_36
timestamp 1621261055
transform 1 0 4608 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_44
timestamp 1621261055
transform 1 0 5376 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_52
timestamp 1621261055
transform 1 0 6144 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_60
timestamp 1621261055
transform 1 0 6912 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_679
timestamp 1621261055
transform 1 0 9120 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_68
timestamp 1621261055
transform 1 0 7680 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_76
timestamp 1621261055
transform 1 0 8448 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_80
timestamp 1621261055
transform 1 0 8832 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_82
timestamp 1621261055
transform 1 0 9024 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_84
timestamp 1621261055
transform 1 0 9216 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_92
timestamp 1621261055
transform 1 0 9984 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_100
timestamp 1621261055
transform 1 0 10752 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_108
timestamp 1621261055
transform 1 0 11520 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_116
timestamp 1621261055
transform 1 0 12288 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_124
timestamp 1621261055
transform 1 0 13056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_132
timestamp 1621261055
transform 1 0 13824 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_680
timestamp 1621261055
transform 1 0 14400 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_136
timestamp 1621261055
transform 1 0 14208 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_139
timestamp 1621261055
transform 1 0 14496 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_147
timestamp 1621261055
transform 1 0 15264 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_155
timestamp 1621261055
transform 1 0 16032 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_163
timestamp 1621261055
transform 1 0 16800 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _103_
timestamp 1621261055
transform 1 0 17568 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_681
timestamp 1621261055
transform 1 0 19680 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_174
timestamp 1621261055
transform 1 0 17856 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_182
timestamp 1621261055
transform 1 0 18624 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_190
timestamp 1621261055
transform 1 0 19392 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_192
timestamp 1621261055
transform 1 0 19584 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_194
timestamp 1621261055
transform 1 0 19776 0 -1 35298
box -38 -49 806 715
use OR2X1  OR2X1
timestamp 1623610208
transform -1 0 22176 0 -1 35298
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_109
timestamp 1621261055
transform -1 0 21024 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_202
timestamp 1621261055
transform 1 0 20544 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_204
timestamp 1621261055
transform 1 0 20736 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_219
timestamp 1621261055
transform 1 0 22176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_227
timestamp 1621261055
transform 1 0 22944 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_682
timestamp 1621261055
transform 1 0 24960 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_235
timestamp 1621261055
transform 1 0 23712 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_243
timestamp 1621261055
transform 1 0 24480 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_48_247
timestamp 1621261055
transform 1 0 24864 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_249
timestamp 1621261055
transform 1 0 25056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_257
timestamp 1621261055
transform 1 0 25824 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_265
timestamp 1621261055
transform 1 0 26592 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_273
timestamp 1621261055
transform 1 0 27360 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_281
timestamp 1621261055
transform 1 0 28128 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_289
timestamp 1621261055
transform 1 0 28896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_297
timestamp 1621261055
transform 1 0 29664 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_683
timestamp 1621261055
transform 1 0 30240 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_301
timestamp 1621261055
transform 1 0 30048 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_304
timestamp 1621261055
transform 1 0 30336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_312
timestamp 1621261055
transform 1 0 31104 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_320
timestamp 1621261055
transform 1 0 31872 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_328
timestamp 1621261055
transform 1 0 32640 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_684
timestamp 1621261055
transform 1 0 35520 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_336
timestamp 1621261055
transform 1 0 33408 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_344
timestamp 1621261055
transform 1 0 34176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_352
timestamp 1621261055
transform 1 0 34944 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_356
timestamp 1621261055
transform 1 0 35328 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_359
timestamp 1621261055
transform 1 0 35616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_367
timestamp 1621261055
transform 1 0 36384 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_375
timestamp 1621261055
transform 1 0 37152 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_383
timestamp 1621261055
transform 1 0 37920 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_391
timestamp 1621261055
transform 1 0 38688 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_685
timestamp 1621261055
transform 1 0 40800 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_399
timestamp 1621261055
transform 1 0 39456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_407
timestamp 1621261055
transform 1 0 40224 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_411
timestamp 1621261055
transform 1 0 40608 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_414
timestamp 1621261055
transform 1 0 40896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_422
timestamp 1621261055
transform 1 0 41664 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_430
timestamp 1621261055
transform 1 0 42432 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_438
timestamp 1621261055
transform 1 0 43200 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_446
timestamp 1621261055
transform 1 0 43968 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_454
timestamp 1621261055
transform 1 0 44736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_462
timestamp 1621261055
transform 1 0 45504 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_686
timestamp 1621261055
transform 1 0 46080 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_466
timestamp 1621261055
transform 1 0 45888 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_469
timestamp 1621261055
transform 1 0 46176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_477
timestamp 1621261055
transform 1 0 46944 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_485
timestamp 1621261055
transform 1 0 47712 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_493
timestamp 1621261055
transform 1 0 48480 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _071_
timestamp 1621261055
transform -1 0 50496 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_687
timestamp 1621261055
transform 1 0 51360 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_105
timestamp 1621261055
transform -1 0 50208 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_501
timestamp 1621261055
transform 1 0 49248 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_514
timestamp 1621261055
transform 1 0 50496 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_48_522
timestamp 1621261055
transform 1 0 51264 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_524
timestamp 1621261055
transform 1 0 51456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_532
timestamp 1621261055
transform 1 0 52224 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_540
timestamp 1621261055
transform 1 0 52992 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_548
timestamp 1621261055
transform 1 0 53760 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_556
timestamp 1621261055
transform 1 0 54528 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_688
timestamp 1621261055
transform 1 0 56640 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_564
timestamp 1621261055
transform 1 0 55296 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_572
timestamp 1621261055
transform 1 0 56064 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_576
timestamp 1621261055
transform 1 0 56448 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_579
timestamp 1621261055
transform 1 0 56736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_587
timestamp 1621261055
transform 1 0 57504 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_97
timestamp 1621261055
transform -1 0 58848 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_595
timestamp 1621261055
transform 1 0 58272 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _125_
timestamp 1621261055
transform 1 0 2400 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_98
timestamp 1621261055
transform 1 0 1152 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_160
timestamp 1621261055
transform 1 0 2208 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_49_4
timestamp 1621261055
transform 1 0 1536 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_8
timestamp 1621261055
transform 1 0 1920 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_10
timestamp 1621261055
transform 1 0 2112 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_16
timestamp 1621261055
transform 1 0 2688 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_24
timestamp 1621261055
transform 1 0 3456 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_32
timestamp 1621261055
transform 1 0 4224 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_689
timestamp 1621261055
transform 1 0 6432 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_40
timestamp 1621261055
transform 1 0 4992 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_48
timestamp 1621261055
transform 1 0 5760 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_52
timestamp 1621261055
transform 1 0 6144 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_54
timestamp 1621261055
transform 1 0 6336 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_56
timestamp 1621261055
transform 1 0 6528 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_64
timestamp 1621261055
transform 1 0 7296 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _004_
timestamp 1621261055
transform 1 0 9408 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_49_72
timestamp 1621261055
transform 1 0 8064 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_80
timestamp 1621261055
transform 1 0 8832 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_84
timestamp 1621261055
transform 1 0 9216 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_89
timestamp 1621261055
transform 1 0 9696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_97
timestamp 1621261055
transform 1 0 10464 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_690
timestamp 1621261055
transform 1 0 11712 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_105
timestamp 1621261055
transform 1 0 11232 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_49_109
timestamp 1621261055
transform 1 0 11616 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_111
timestamp 1621261055
transform 1 0 11808 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_119
timestamp 1621261055
transform 1 0 12576 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_127
timestamp 1621261055
transform 1 0 13344 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_691
timestamp 1621261055
transform 1 0 16992 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_135
timestamp 1621261055
transform 1 0 14112 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_143
timestamp 1621261055
transform 1 0 14880 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_151
timestamp 1621261055
transform 1 0 15648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_159
timestamp 1621261055
transform 1 0 16416 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_163
timestamp 1621261055
transform 1 0 16800 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_166
timestamp 1621261055
transform 1 0 17088 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_174
timestamp 1621261055
transform 1 0 17856 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_182
timestamp 1621261055
transform 1 0 18624 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_190
timestamp 1621261055
transform 1 0 19392 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_49_198
timestamp 1621261055
transform 1 0 20160 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_206
timestamp 1621261055
transform 1 0 20928 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_49_202
timestamp 1621261055
transform 1 0 20544 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _166_
timestamp 1621261055
transform 1 0 20256 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_49_214
timestamp 1621261055
transform 1 0 21696 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_49_208
timestamp 1621261055
transform 1 0 21120 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_144
timestamp 1621261055
transform 1 0 21216 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _115_
timestamp 1621261055
transform 1 0 21408 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_49_221
timestamp 1621261055
transform 1 0 22368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_218
timestamp 1621261055
transform 1 0 22080 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_692
timestamp 1621261055
transform 1 0 22272 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_229
timestamp 1621261055
transform 1 0 23136 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_237
timestamp 1621261055
transform 1 0 23904 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_245
timestamp 1621261055
transform 1 0 24672 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_253
timestamp 1621261055
transform 1 0 25440 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_261
timestamp 1621261055
transform 1 0 26208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_693
timestamp 1621261055
transform 1 0 27552 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_269
timestamp 1621261055
transform 1 0 26976 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_273
timestamp 1621261055
transform 1 0 27360 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_276
timestamp 1621261055
transform 1 0 27648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_284
timestamp 1621261055
transform 1 0 28416 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_292
timestamp 1621261055
transform 1 0 29184 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_694
timestamp 1621261055
transform 1 0 32832 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_300
timestamp 1621261055
transform 1 0 29952 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_308
timestamp 1621261055
transform 1 0 30720 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_316
timestamp 1621261055
transform 1 0 31488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_324
timestamp 1621261055
transform 1 0 32256 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_328
timestamp 1621261055
transform 1 0 32640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_331
timestamp 1621261055
transform 1 0 32928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_339
timestamp 1621261055
transform 1 0 33696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_347
timestamp 1621261055
transform 1 0 34464 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_355
timestamp 1621261055
transform 1 0 35232 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_363
timestamp 1621261055
transform 1 0 36000 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_695
timestamp 1621261055
transform 1 0 38112 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_371
timestamp 1621261055
transform 1 0 36768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_379
timestamp 1621261055
transform 1 0 37536 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_383
timestamp 1621261055
transform 1 0 37920 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_386
timestamp 1621261055
transform 1 0 38208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_394
timestamp 1621261055
transform 1 0 38976 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_402
timestamp 1621261055
transform 1 0 39744 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_410
timestamp 1621261055
transform 1 0 40512 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_418
timestamp 1621261055
transform 1 0 41280 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_426
timestamp 1621261055
transform 1 0 42048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _134_
timestamp 1621261055
transform -1 0 45312 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_696
timestamp 1621261055
transform 1 0 43392 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_170
timestamp 1621261055
transform -1 0 45024 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_49_434
timestamp 1621261055
transform 1 0 42816 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_438
timestamp 1621261055
transform 1 0 43200 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_441
timestamp 1621261055
transform 1 0 43488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_449
timestamp 1621261055
transform 1 0 44256 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_453
timestamp 1621261055
transform 1 0 44640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_460
timestamp 1621261055
transform 1 0 45312 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_697
timestamp 1621261055
transform 1 0 48672 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_468
timestamp 1621261055
transform 1 0 46080 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_476
timestamp 1621261055
transform 1 0 46848 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_484
timestamp 1621261055
transform 1 0 47616 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_492
timestamp 1621261055
transform 1 0 48384 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_494
timestamp 1621261055
transform 1 0 48576 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _097_
timestamp 1621261055
transform -1 0 51648 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _147_
timestamp 1621261055
transform -1 0 49440 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_133
timestamp 1621261055
transform -1 0 51360 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_181
timestamp 1621261055
transform -1 0 49152 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_496
timestamp 1621261055
transform 1 0 48768 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_503
timestamp 1621261055
transform 1 0 49440 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_511
timestamp 1621261055
transform 1 0 50208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_519
timestamp 1621261055
transform 1 0 50976 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_526
timestamp 1621261055
transform 1 0 51648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_698
timestamp 1621261055
transform 1 0 53952 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_534
timestamp 1621261055
transform 1 0 52416 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_542
timestamp 1621261055
transform 1 0 53184 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_551
timestamp 1621261055
transform 1 0 54048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_559
timestamp 1621261055
transform 1 0 54816 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_567
timestamp 1621261055
transform 1 0 55584 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_575
timestamp 1621261055
transform 1 0 56352 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_583
timestamp 1621261055
transform 1 0 57120 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_591
timestamp 1621261055
transform 1 0 57888 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_99
timestamp 1621261055
transform -1 0 58848 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_595
timestamp 1621261055
transform 1 0 58272 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_146
timestamp 1621261055
transform 1 0 1536 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_100
timestamp 1621261055
transform 1 0 1152 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _116_
timestamp 1621261055
transform 1 0 1728 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_50_15
timestamp 1621261055
transform 1 0 2592 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_13
timestamp 1621261055
transform 1 0 2400 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_9
timestamp 1621261055
transform 1 0 2016 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _000_
timestamp 1621261055
transform 1 0 2688 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_50_19
timestamp 1621261055
transform 1 0 2976 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_29
timestamp 1621261055
transform 1 0 3936 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_50_27
timestamp 1621261055
transform 1 0 3744 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_699
timestamp 1621261055
transform 1 0 3840 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_37
timestamp 1621261055
transform 1 0 4704 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_45
timestamp 1621261055
transform 1 0 5472 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_53
timestamp 1621261055
transform 1 0 6240 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_61
timestamp 1621261055
transform 1 0 7008 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_700
timestamp 1621261055
transform 1 0 9120 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_69
timestamp 1621261055
transform 1 0 7776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_77
timestamp 1621261055
transform 1 0 8544 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_81
timestamp 1621261055
transform 1 0 8928 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_84
timestamp 1621261055
transform 1 0 9216 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_92
timestamp 1621261055
transform 1 0 9984 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_100
timestamp 1621261055
transform 1 0 10752 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_108
timestamp 1621261055
transform 1 0 11520 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_116
timestamp 1621261055
transform 1 0 12288 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_124
timestamp 1621261055
transform 1 0 13056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_132
timestamp 1621261055
transform 1 0 13824 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_701
timestamp 1621261055
transform 1 0 14400 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_136
timestamp 1621261055
transform 1 0 14208 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_139
timestamp 1621261055
transform 1 0 14496 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_147
timestamp 1621261055
transform 1 0 15264 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_155
timestamp 1621261055
transform 1 0 16032 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_163
timestamp 1621261055
transform 1 0 16800 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_702
timestamp 1621261055
transform 1 0 19680 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_171
timestamp 1621261055
transform 1 0 17568 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_179
timestamp 1621261055
transform 1 0 18336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_187
timestamp 1621261055
transform 1 0 19104 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_191
timestamp 1621261055
transform 1 0 19488 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_194
timestamp 1621261055
transform 1 0 19776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _200_
timestamp 1621261055
transform -1 0 22848 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_202
timestamp 1621261055
transform -1 0 22560 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_202
timestamp 1621261055
transform 1 0 20544 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_210
timestamp 1621261055
transform 1 0 21312 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_218
timestamp 1621261055
transform 1 0 22080 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_220
timestamp 1621261055
transform 1 0 22272 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_226
timestamp 1621261055
transform 1 0 22848 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_703
timestamp 1621261055
transform 1 0 24960 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_234
timestamp 1621261055
transform 1 0 23616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_242
timestamp 1621261055
transform 1 0 24384 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_246
timestamp 1621261055
transform 1 0 24768 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_249
timestamp 1621261055
transform 1 0 25056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_257
timestamp 1621261055
transform 1 0 25824 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_265
timestamp 1621261055
transform 1 0 26592 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_273
timestamp 1621261055
transform 1 0 27360 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_281
timestamp 1621261055
transform 1 0 28128 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_289
timestamp 1621261055
transform 1 0 28896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_297
timestamp 1621261055
transform 1 0 29664 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_704
timestamp 1621261055
transform 1 0 30240 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_301
timestamp 1621261055
transform 1 0 30048 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_304
timestamp 1621261055
transform 1 0 30336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_312
timestamp 1621261055
transform 1 0 31104 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_320
timestamp 1621261055
transform 1 0 31872 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_328
timestamp 1621261055
transform 1 0 32640 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_705
timestamp 1621261055
transform 1 0 35520 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_336
timestamp 1621261055
transform 1 0 33408 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_344
timestamp 1621261055
transform 1 0 34176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_352
timestamp 1621261055
transform 1 0 34944 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_356
timestamp 1621261055
transform 1 0 35328 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_359
timestamp 1621261055
transform 1 0 35616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _172_
timestamp 1621261055
transform 1 0 38304 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_50_367
timestamp 1621261055
transform 1 0 36384 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_375
timestamp 1621261055
transform 1 0 37152 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_383
timestamp 1621261055
transform 1 0 37920 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_390
timestamp 1621261055
transform 1 0 38592 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_706
timestamp 1621261055
transform 1 0 40800 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_398
timestamp 1621261055
transform 1 0 39360 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_406
timestamp 1621261055
transform 1 0 40128 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_410
timestamp 1621261055
transform 1 0 40512 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_412
timestamp 1621261055
transform 1 0 40704 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_414
timestamp 1621261055
transform 1 0 40896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_422
timestamp 1621261055
transform 1 0 41664 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_430
timestamp 1621261055
transform 1 0 42432 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_438
timestamp 1621261055
transform 1 0 43200 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_446
timestamp 1621261055
transform 1 0 43968 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_454
timestamp 1621261055
transform 1 0 44736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_462
timestamp 1621261055
transform 1 0 45504 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_707
timestamp 1621261055
transform 1 0 46080 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_466
timestamp 1621261055
transform 1 0 45888 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_469
timestamp 1621261055
transform 1 0 46176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_477
timestamp 1621261055
transform 1 0 46944 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_485
timestamp 1621261055
transform 1 0 47712 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_493
timestamp 1621261055
transform 1 0 48480 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_708
timestamp 1621261055
transform 1 0 51360 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_501
timestamp 1621261055
transform 1 0 49248 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_509
timestamp 1621261055
transform 1 0 50016 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_517
timestamp 1621261055
transform 1 0 50784 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_521
timestamp 1621261055
transform 1 0 51168 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_524
timestamp 1621261055
transform 1 0 51456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _182_
timestamp 1621261055
transform -1 0 55104 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_192
timestamp 1621261055
transform -1 0 54816 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_532
timestamp 1621261055
transform 1 0 52224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_540
timestamp 1621261055
transform 1 0 52992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_548
timestamp 1621261055
transform 1 0 53760 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_50_556
timestamp 1621261055
transform 1 0 54528 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_709
timestamp 1621261055
transform 1 0 56640 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_562
timestamp 1621261055
transform 1 0 55104 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_570
timestamp 1621261055
transform 1 0 55872 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_579
timestamp 1621261055
transform 1 0 56736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_587
timestamp 1621261055
transform 1 0 57504 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_101
timestamp 1621261055
transform -1 0 58848 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_595
timestamp 1621261055
transform 1 0 58272 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_102
timestamp 1621261055
transform 1 0 1152 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_4
timestamp 1621261055
transform 1 0 1536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_12
timestamp 1621261055
transform 1 0 2304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_20
timestamp 1621261055
transform 1 0 3072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_28
timestamp 1621261055
transform 1 0 3840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_710
timestamp 1621261055
transform 1 0 6432 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_36
timestamp 1621261055
transform 1 0 4608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_44
timestamp 1621261055
transform 1 0 5376 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_52
timestamp 1621261055
transform 1 0 6144 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_54
timestamp 1621261055
transform 1 0 6336 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_56
timestamp 1621261055
transform 1 0 6528 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_64
timestamp 1621261055
transform 1 0 7296 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_72
timestamp 1621261055
transform 1 0 8064 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_80
timestamp 1621261055
transform 1 0 8832 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_88
timestamp 1621261055
transform 1 0 9600 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_96
timestamp 1621261055
transform 1 0 10368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_711
timestamp 1621261055
transform 1 0 11712 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_104
timestamp 1621261055
transform 1 0 11136 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_108
timestamp 1621261055
transform 1 0 11520 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_111
timestamp 1621261055
transform 1 0 11808 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_119
timestamp 1621261055
transform 1 0 12576 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_127
timestamp 1621261055
transform 1 0 13344 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_712
timestamp 1621261055
transform 1 0 16992 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_135
timestamp 1621261055
transform 1 0 14112 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_143
timestamp 1621261055
transform 1 0 14880 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_151
timestamp 1621261055
transform 1 0 15648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_159
timestamp 1621261055
transform 1 0 16416 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_163
timestamp 1621261055
transform 1 0 16800 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_166
timestamp 1621261055
transform 1 0 17088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_174
timestamp 1621261055
transform 1 0 17856 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_182
timestamp 1621261055
transform 1 0 18624 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_190
timestamp 1621261055
transform 1 0 19392 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_198
timestamp 1621261055
transform 1 0 20160 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_713
timestamp 1621261055
transform 1 0 22272 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_206
timestamp 1621261055
transform 1 0 20928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_214
timestamp 1621261055
transform 1 0 21696 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_218
timestamp 1621261055
transform 1 0 22080 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_221
timestamp 1621261055
transform 1 0 22368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_229
timestamp 1621261055
transform 1 0 23136 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_237
timestamp 1621261055
transform 1 0 23904 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_245
timestamp 1621261055
transform 1 0 24672 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_253
timestamp 1621261055
transform 1 0 25440 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_261
timestamp 1621261055
transform 1 0 26208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_714
timestamp 1621261055
transform 1 0 27552 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_269
timestamp 1621261055
transform 1 0 26976 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_273
timestamp 1621261055
transform 1 0 27360 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_276
timestamp 1621261055
transform 1 0 27648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_284
timestamp 1621261055
transform 1 0 28416 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_292
timestamp 1621261055
transform 1 0 29184 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_715
timestamp 1621261055
transform 1 0 32832 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_300
timestamp 1621261055
transform 1 0 29952 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_308
timestamp 1621261055
transform 1 0 30720 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_316
timestamp 1621261055
transform 1 0 31488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_324
timestamp 1621261055
transform 1 0 32256 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_328
timestamp 1621261055
transform 1 0 32640 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_331
timestamp 1621261055
transform 1 0 32928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_339
timestamp 1621261055
transform 1 0 33696 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_347
timestamp 1621261055
transform 1 0 34464 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_355
timestamp 1621261055
transform 1 0 35232 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_363
timestamp 1621261055
transform 1 0 36000 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_716
timestamp 1621261055
transform 1 0 38112 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_371
timestamp 1621261055
transform 1 0 36768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_379
timestamp 1621261055
transform 1 0 37536 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_383
timestamp 1621261055
transform 1 0 37920 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_386
timestamp 1621261055
transform 1 0 38208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_394
timestamp 1621261055
transform 1 0 38976 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_402
timestamp 1621261055
transform 1 0 39744 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_410
timestamp 1621261055
transform 1 0 40512 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_418
timestamp 1621261055
transform 1 0 41280 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_426
timestamp 1621261055
transform 1 0 42048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_717
timestamp 1621261055
transform 1 0 43392 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_434
timestamp 1621261055
transform 1 0 42816 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_438
timestamp 1621261055
transform 1 0 43200 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_441
timestamp 1621261055
transform 1 0 43488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_449
timestamp 1621261055
transform 1 0 44256 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_457
timestamp 1621261055
transform 1 0 45024 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_718
timestamp 1621261055
transform 1 0 48672 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_465
timestamp 1621261055
transform 1 0 45792 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_473
timestamp 1621261055
transform 1 0 46560 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_481
timestamp 1621261055
transform 1 0 47328 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_489
timestamp 1621261055
transform 1 0 48096 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_493
timestamp 1621261055
transform 1 0 48480 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_496
timestamp 1621261055
transform 1 0 48768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_504
timestamp 1621261055
transform 1 0 49536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_512
timestamp 1621261055
transform 1 0 50304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_520
timestamp 1621261055
transform 1 0 51072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_528
timestamp 1621261055
transform 1 0 51840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_719
timestamp 1621261055
transform 1 0 53952 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_536
timestamp 1621261055
transform 1 0 52608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_544
timestamp 1621261055
transform 1 0 53376 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_548
timestamp 1621261055
transform 1 0 53760 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_551
timestamp 1621261055
transform 1 0 54048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_559
timestamp 1621261055
transform 1 0 54816 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_567
timestamp 1621261055
transform 1 0 55584 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_575
timestamp 1621261055
transform 1 0 56352 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_583
timestamp 1621261055
transform 1 0 57120 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_591
timestamp 1621261055
transform 1 0 57888 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_103
timestamp 1621261055
transform -1 0 58848 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_595
timestamp 1621261055
transform 1 0 58272 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_104
timestamp 1621261055
transform 1 0 1152 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_720
timestamp 1621261055
transform 1 0 3840 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_4
timestamp 1621261055
transform 1 0 1536 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_12
timestamp 1621261055
transform 1 0 2304 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_20
timestamp 1621261055
transform 1 0 3072 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_29
timestamp 1621261055
transform 1 0 3936 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_37
timestamp 1621261055
transform 1 0 4704 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_45
timestamp 1621261055
transform 1 0 5472 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_53
timestamp 1621261055
transform 1 0 6240 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_61
timestamp 1621261055
transform 1 0 7008 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_721
timestamp 1621261055
transform 1 0 9120 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_69
timestamp 1621261055
transform 1 0 7776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_77
timestamp 1621261055
transform 1 0 8544 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_81
timestamp 1621261055
transform 1 0 8928 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_84
timestamp 1621261055
transform 1 0 9216 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_92
timestamp 1621261055
transform 1 0 9984 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_100
timestamp 1621261055
transform 1 0 10752 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_108
timestamp 1621261055
transform 1 0 11520 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_116
timestamp 1621261055
transform 1 0 12288 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_124
timestamp 1621261055
transform 1 0 13056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_132
timestamp 1621261055
transform 1 0 13824 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _199_
timestamp 1621261055
transform -1 0 16704 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_722
timestamp 1621261055
transform 1 0 14400 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_200
timestamp 1621261055
transform -1 0 16416 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_136
timestamp 1621261055
transform 1 0 14208 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_139
timestamp 1621261055
transform 1 0 14496 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_147
timestamp 1621261055
transform 1 0 15264 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_155
timestamp 1621261055
transform 1 0 16032 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_162
timestamp 1621261055
transform 1 0 16704 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_723
timestamp 1621261055
transform 1 0 19680 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_170
timestamp 1621261055
transform 1 0 17472 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_178
timestamp 1621261055
transform 1 0 18240 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_186
timestamp 1621261055
transform 1 0 19008 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_190
timestamp 1621261055
transform 1 0 19392 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_192
timestamp 1621261055
transform 1 0 19584 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_194
timestamp 1621261055
transform 1 0 19776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_202
timestamp 1621261055
transform 1 0 20544 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_210
timestamp 1621261055
transform 1 0 21312 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_218
timestamp 1621261055
transform 1 0 22080 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_226
timestamp 1621261055
transform 1 0 22848 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_724
timestamp 1621261055
transform 1 0 24960 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_234
timestamp 1621261055
transform 1 0 23616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_242
timestamp 1621261055
transform 1 0 24384 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_246
timestamp 1621261055
transform 1 0 24768 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_249
timestamp 1621261055
transform 1 0 25056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_257
timestamp 1621261055
transform 1 0 25824 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_265
timestamp 1621261055
transform 1 0 26592 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_273
timestamp 1621261055
transform 1 0 27360 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_281
timestamp 1621261055
transform 1 0 28128 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_289
timestamp 1621261055
transform 1 0 28896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_297
timestamp 1621261055
transform 1 0 29664 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_725
timestamp 1621261055
transform 1 0 30240 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_301
timestamp 1621261055
transform 1 0 30048 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_304
timestamp 1621261055
transform 1 0 30336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_312
timestamp 1621261055
transform 1 0 31104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_320
timestamp 1621261055
transform 1 0 31872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_328
timestamp 1621261055
transform 1 0 32640 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_726
timestamp 1621261055
transform 1 0 35520 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_336
timestamp 1621261055
transform 1 0 33408 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_344
timestamp 1621261055
transform 1 0 34176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_352
timestamp 1621261055
transform 1 0 34944 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_356
timestamp 1621261055
transform 1 0 35328 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_359
timestamp 1621261055
transform 1 0 35616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_367
timestamp 1621261055
transform 1 0 36384 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_375
timestamp 1621261055
transform 1 0 37152 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_383
timestamp 1621261055
transform 1 0 37920 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_391
timestamp 1621261055
transform 1 0 38688 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _175_
timestamp 1621261055
transform 1 0 41568 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_727
timestamp 1621261055
transform 1 0 40800 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_93
timestamp 1621261055
transform 1 0 41376 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_399
timestamp 1621261055
transform 1 0 39456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_407
timestamp 1621261055
transform 1 0 40224 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_411
timestamp 1621261055
transform 1 0 40608 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_52_414
timestamp 1621261055
transform 1 0 40896 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_52_418
timestamp 1621261055
transform 1 0 41280 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_424
timestamp 1621261055
transform 1 0 41856 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _073_
timestamp 1621261055
transform -1 0 43488 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_111
timestamp 1621261055
transform -1 0 43200 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_52_432
timestamp 1621261055
transform 1 0 42624 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_441
timestamp 1621261055
transform 1 0 43488 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_449
timestamp 1621261055
transform 1 0 44256 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_457
timestamp 1621261055
transform 1 0 45024 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_728
timestamp 1621261055
transform 1 0 46080 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_465
timestamp 1621261055
transform 1 0 45792 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_467
timestamp 1621261055
transform 1 0 45984 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_469
timestamp 1621261055
transform 1 0 46176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_477
timestamp 1621261055
transform 1 0 46944 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_485
timestamp 1621261055
transform 1 0 47712 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_493
timestamp 1621261055
transform 1 0 48480 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_729
timestamp 1621261055
transform 1 0 51360 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_501
timestamp 1621261055
transform 1 0 49248 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_509
timestamp 1621261055
transform 1 0 50016 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_517
timestamp 1621261055
transform 1 0 50784 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_521
timestamp 1621261055
transform 1 0 51168 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_524
timestamp 1621261055
transform 1 0 51456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _196_
timestamp 1621261055
transform -1 0 54336 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_196
timestamp 1621261055
transform -1 0 54048 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_532
timestamp 1621261055
transform 1 0 52224 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_540
timestamp 1621261055
transform 1 0 52992 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_52_548
timestamp 1621261055
transform 1 0 53760 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_554
timestamp 1621261055
transform 1 0 54336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_730
timestamp 1621261055
transform 1 0 56640 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_562
timestamp 1621261055
transform 1 0 55104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_570
timestamp 1621261055
transform 1 0 55872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_579
timestamp 1621261055
transform 1 0 56736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_587
timestamp 1621261055
transform 1 0 57504 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_105
timestamp 1621261055
transform -1 0 58848 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_595
timestamp 1621261055
transform 1 0 58272 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_106
timestamp 1621261055
transform 1 0 1152 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_4
timestamp 1621261055
transform 1 0 1536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_12
timestamp 1621261055
transform 1 0 2304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_20
timestamp 1621261055
transform 1 0 3072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_28
timestamp 1621261055
transform 1 0 3840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_731
timestamp 1621261055
transform 1 0 6432 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_36
timestamp 1621261055
transform 1 0 4608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_44
timestamp 1621261055
transform 1 0 5376 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_52
timestamp 1621261055
transform 1 0 6144 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_54
timestamp 1621261055
transform 1 0 6336 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_56
timestamp 1621261055
transform 1 0 6528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_64
timestamp 1621261055
transform 1 0 7296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_72
timestamp 1621261055
transform 1 0 8064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_80
timestamp 1621261055
transform 1 0 8832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_88
timestamp 1621261055
transform 1 0 9600 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_96
timestamp 1621261055
transform 1 0 10368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_732
timestamp 1621261055
transform 1 0 11712 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_104
timestamp 1621261055
transform 1 0 11136 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_108
timestamp 1621261055
transform 1 0 11520 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_111
timestamp 1621261055
transform 1 0 11808 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_119
timestamp 1621261055
transform 1 0 12576 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_127
timestamp 1621261055
transform 1 0 13344 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _021_
timestamp 1621261055
transform 1 0 15936 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_733
timestamp 1621261055
transform 1 0 16992 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_135
timestamp 1621261055
transform 1 0 14112 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_143
timestamp 1621261055
transform 1 0 14880 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_151
timestamp 1621261055
transform 1 0 15648 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_153
timestamp 1621261055
transform 1 0 15840 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_157
timestamp 1621261055
transform 1 0 16224 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_166
timestamp 1621261055
transform 1 0 17088 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_174
timestamp 1621261055
transform 1 0 17856 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_182
timestamp 1621261055
transform 1 0 18624 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_190
timestamp 1621261055
transform 1 0 19392 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_198
timestamp 1621261055
transform 1 0 20160 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_734
timestamp 1621261055
transform 1 0 22272 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_206
timestamp 1621261055
transform 1 0 20928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_214
timestamp 1621261055
transform 1 0 21696 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_218
timestamp 1621261055
transform 1 0 22080 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_221
timestamp 1621261055
transform 1 0 22368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_229
timestamp 1621261055
transform 1 0 23136 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_237
timestamp 1621261055
transform 1 0 23904 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_245
timestamp 1621261055
transform 1 0 24672 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_253
timestamp 1621261055
transform 1 0 25440 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_261
timestamp 1621261055
transform 1 0 26208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_735
timestamp 1621261055
transform 1 0 27552 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_269
timestamp 1621261055
transform 1 0 26976 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_273
timestamp 1621261055
transform 1 0 27360 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_276
timestamp 1621261055
transform 1 0 27648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_284
timestamp 1621261055
transform 1 0 28416 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_292
timestamp 1621261055
transform 1 0 29184 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _118_
timestamp 1621261055
transform 1 0 30336 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_736
timestamp 1621261055
transform 1 0 32832 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_150
timestamp 1621261055
transform 1 0 30144 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_300
timestamp 1621261055
transform 1 0 29952 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_307
timestamp 1621261055
transform 1 0 30624 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_315
timestamp 1621261055
transform 1 0 31392 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_323
timestamp 1621261055
transform 1 0 32160 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_327
timestamp 1621261055
transform 1 0 32544 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_329
timestamp 1621261055
transform 1 0 32736 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_331
timestamp 1621261055
transform 1 0 32928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_339
timestamp 1621261055
transform 1 0 33696 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_347
timestamp 1621261055
transform 1 0 34464 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_355
timestamp 1621261055
transform 1 0 35232 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_363
timestamp 1621261055
transform 1 0 36000 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_737
timestamp 1621261055
transform 1 0 38112 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_371
timestamp 1621261055
transform 1 0 36768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_379
timestamp 1621261055
transform 1 0 37536 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_383
timestamp 1621261055
transform 1 0 37920 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_386
timestamp 1621261055
transform 1 0 38208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_394
timestamp 1621261055
transform 1 0 38976 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_402
timestamp 1621261055
transform 1 0 39744 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_410
timestamp 1621261055
transform 1 0 40512 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_418
timestamp 1621261055
transform 1 0 41280 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_426
timestamp 1621261055
transform 1 0 42048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_738
timestamp 1621261055
transform 1 0 43392 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_434
timestamp 1621261055
transform 1 0 42816 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_438
timestamp 1621261055
transform 1 0 43200 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_441
timestamp 1621261055
transform 1 0 43488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_449
timestamp 1621261055
transform 1 0 44256 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_457
timestamp 1621261055
transform 1 0 45024 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_739
timestamp 1621261055
transform 1 0 48672 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_465
timestamp 1621261055
transform 1 0 45792 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_473
timestamp 1621261055
transform 1 0 46560 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_481
timestamp 1621261055
transform 1 0 47328 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_489
timestamp 1621261055
transform 1 0 48096 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_493
timestamp 1621261055
transform 1 0 48480 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _027_
timestamp 1621261055
transform 1 0 51840 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_53_496
timestamp 1621261055
transform 1 0 48768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_504
timestamp 1621261055
transform 1 0 49536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_512
timestamp 1621261055
transform 1 0 50304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_520
timestamp 1621261055
transform 1 0 51072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_740
timestamp 1621261055
transform 1 0 53952 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_531
timestamp 1621261055
transform 1 0 52128 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_539
timestamp 1621261055
transform 1 0 52896 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_547
timestamp 1621261055
transform 1 0 53664 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_549
timestamp 1621261055
transform 1 0 53856 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_551
timestamp 1621261055
transform 1 0 54048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_559
timestamp 1621261055
transform 1 0 54816 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _083_
timestamp 1621261055
transform -1 0 58080 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_121
timestamp 1621261055
transform -1 0 57792 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_567
timestamp 1621261055
transform 1 0 55584 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_575
timestamp 1621261055
transform 1 0 56352 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_583
timestamp 1621261055
transform 1 0 57120 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_53_587
timestamp 1621261055
transform 1 0 57504 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_593
timestamp 1621261055
transform 1 0 58080 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_107
timestamp 1621261055
transform -1 0 58848 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_4
timestamp 1621261055
transform 1 0 1536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_4
timestamp 1621261055
transform 1 0 1536 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_110
timestamp 1621261055
transform 1 0 1152 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_108
timestamp 1621261055
transform 1 0 1152 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_12
timestamp 1621261055
transform 1 0 2304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_12
timestamp 1621261055
transform 1 0 2304 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_20
timestamp 1621261055
transform 1 0 3072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_20
timestamp 1621261055
transform 1 0 3072 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_28
timestamp 1621261055
transform 1 0 3840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_29
timestamp 1621261055
transform 1 0 3936 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_741
timestamp 1621261055
transform 1 0 3840 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_36
timestamp 1621261055
transform 1 0 4608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_37
timestamp 1621261055
transform 1 0 4704 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_44
timestamp 1621261055
transform 1 0 5376 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_50
timestamp 1621261055
transform 1 0 5952 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_45
timestamp 1621261055
transform 1 0 5472 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _028_
timestamp 1621261055
transform 1 0 5664 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_56
timestamp 1621261055
transform 1 0 6528 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_55_54
timestamp 1621261055
transform 1 0 6336 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_52
timestamp 1621261055
transform 1 0 6144 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_58
timestamp 1621261055
transform 1 0 6720 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_752
timestamp 1621261055
transform 1 0 6432 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_64
timestamp 1621261055
transform 1 0 7296 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_66
timestamp 1621261055
transform 1 0 7488 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_742
timestamp 1621261055
transform 1 0 9120 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_74
timestamp 1621261055
transform 1 0 8256 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_82
timestamp 1621261055
transform 1 0 9024 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_84
timestamp 1621261055
transform 1 0 9216 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_92
timestamp 1621261055
transform 1 0 9984 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_72
timestamp 1621261055
transform 1 0 8064 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_80
timestamp 1621261055
transform 1 0 8832 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_88
timestamp 1621261055
transform 1 0 9600 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_96
timestamp 1621261055
transform 1 0 10368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_104
timestamp 1621261055
transform 1 0 11136 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_100
timestamp 1621261055
transform 1 0 10752 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_111
timestamp 1621261055
transform 1 0 11808 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_108
timestamp 1621261055
transform 1 0 11520 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_116
timestamp 1621261055
transform 1 0 12288 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_108
timestamp 1621261055
transform 1 0 11520 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_178
timestamp 1621261055
transform 1 0 12000 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_753
timestamp 1621261055
transform 1 0 11712 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _142_
timestamp 1621261055
transform 1 0 12192 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_118
timestamp 1621261055
transform 1 0 12480 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_124
timestamp 1621261055
transform 1 0 13056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_126
timestamp 1621261055
transform 1 0 13248 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_132
timestamp 1621261055
transform 1 0 13824 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_134
timestamp 1621261055
transform 1 0 14016 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_139
timestamp 1621261055
transform 1 0 14496 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_136
timestamp 1621261055
transform 1 0 14208 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_743
timestamp 1621261055
transform 1 0 14400 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_142
timestamp 1621261055
transform 1 0 14784 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_147
timestamp 1621261055
transform 1 0 15264 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_158
timestamp 1621261055
transform 1 0 16320 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_150
timestamp 1621261055
transform 1 0 15552 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_155
timestamp 1621261055
transform 1 0 16032 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_55_164
timestamp 1621261055
transform 1 0 16896 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_162
timestamp 1621261055
transform 1 0 16704 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_163
timestamp 1621261055
transform 1 0 16800 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_754
timestamp 1621261055
transform 1 0 16992 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_166
timestamp 1621261055
transform 1 0 17088 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_171
timestamp 1621261055
transform 1 0 17568 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_182
timestamp 1621261055
transform 1 0 18624 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_174
timestamp 1621261055
transform 1 0 17856 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_179
timestamp 1621261055
transform 1 0 18336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_190
timestamp 1621261055
transform 1 0 19392 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_191
timestamp 1621261055
transform 1 0 19488 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_187
timestamp 1621261055
transform 1 0 19104 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_198
timestamp 1621261055
transform 1 0 20160 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_194
timestamp 1621261055
transform 1 0 19776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_744
timestamp 1621261055
transform 1 0 19680 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_206
timestamp 1621261055
transform 1 0 20928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_206
timestamp 1621261055
transform 1 0 20928 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_202
timestamp 1621261055
transform 1 0 20544 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_55_214
timestamp 1621261055
transform 1 0 21696 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_213
timestamp 1621261055
transform 1 0 21600 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_224
timestamp 1621261055
transform -1 0 21312 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _186_
timestamp 1621261055
transform -1 0 21600 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_221
timestamp 1621261055
transform 1 0 22368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_218
timestamp 1621261055
transform 1 0 22080 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_221
timestamp 1621261055
transform 1 0 22368 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_755
timestamp 1621261055
transform 1 0 22272 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_229
timestamp 1621261055
transform 1 0 23136 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_229
timestamp 1621261055
transform 1 0 23136 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_237
timestamp 1621261055
transform 1 0 23904 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_237
timestamp 1621261055
transform 1 0 23904 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_245
timestamp 1621261055
transform 1 0 24672 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_247
timestamp 1621261055
transform 1 0 24864 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_245
timestamp 1621261055
transform 1 0 24672 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_745
timestamp 1621261055
transform 1 0 24960 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_253
timestamp 1621261055
transform 1 0 25440 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_257
timestamp 1621261055
transform 1 0 25824 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_249
timestamp 1621261055
transform 1 0 25056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_261
timestamp 1621261055
transform 1 0 26208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_269
timestamp 1621261055
transform 1 0 26976 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_272
timestamp 1621261055
transform 1 0 27264 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_265
timestamp 1621261055
transform 1 0 26592 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_158
timestamp 1621261055
transform 1 0 26784 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _124_
timestamp 1621261055
transform 1 0 26976 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_276
timestamp 1621261055
transform 1 0 27648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_273
timestamp 1621261055
transform 1 0 27360 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_280
timestamp 1621261055
transform 1 0 28032 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_756
timestamp 1621261055
transform 1 0 27552 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_284
timestamp 1621261055
transform 1 0 28416 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_288
timestamp 1621261055
transform 1 0 28800 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_292
timestamp 1621261055
transform 1 0 29184 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_296
timestamp 1621261055
transform 1 0 29568 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_300
timestamp 1621261055
transform 1 0 29952 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_304
timestamp 1621261055
transform 1 0 30336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_302
timestamp 1621261055
transform 1 0 30144 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_300
timestamp 1621261055
transform 1 0 29952 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_746
timestamp 1621261055
transform 1 0 30240 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_308
timestamp 1621261055
transform 1 0 30720 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_312
timestamp 1621261055
transform 1 0 31104 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_316
timestamp 1621261055
transform 1 0 31488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_320
timestamp 1621261055
transform 1 0 31872 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_328
timestamp 1621261055
transform 1 0 32640 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_324
timestamp 1621261055
transform 1 0 32256 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_328
timestamp 1621261055
transform 1 0 32640 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_757
timestamp 1621261055
transform 1 0 32832 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_331
timestamp 1621261055
transform 1 0 32928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_336
timestamp 1621261055
transform 1 0 33408 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_347
timestamp 1621261055
transform 1 0 34464 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_339
timestamp 1621261055
transform 1 0 33696 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_344
timestamp 1621261055
transform 1 0 34176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_355
timestamp 1621261055
transform 1 0 35232 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_356
timestamp 1621261055
transform 1 0 35328 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_352
timestamp 1621261055
transform 1 0 34944 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_363
timestamp 1621261055
transform 1 0 36000 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_359
timestamp 1621261055
transform 1 0 35616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_747
timestamp 1621261055
transform 1 0 35520 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_371
timestamp 1621261055
transform 1 0 36768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_367
timestamp 1621261055
transform 1 0 36384 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_379
timestamp 1621261055
transform 1 0 37536 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_375
timestamp 1621261055
transform 1 0 37152 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_386
timestamp 1621261055
transform 1 0 38208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_383
timestamp 1621261055
transform 1 0 37920 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_383
timestamp 1621261055
transform 1 0 37920 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_758
timestamp 1621261055
transform 1 0 38112 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_394
timestamp 1621261055
transform 1 0 38976 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_391
timestamp 1621261055
transform 1 0 38688 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_402
timestamp 1621261055
transform 1 0 39744 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_399
timestamp 1621261055
transform 1 0 39456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_410
timestamp 1621261055
transform 1 0 40512 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_411
timestamp 1621261055
transform 1 0 40608 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_407
timestamp 1621261055
transform 1 0 40224 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_748
timestamp 1621261055
transform 1 0 40800 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_418
timestamp 1621261055
transform 1 0 41280 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_422
timestamp 1621261055
transform 1 0 41664 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_414
timestamp 1621261055
transform 1 0 40896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_426
timestamp 1621261055
transform 1 0 42048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_434
timestamp 1621261055
transform 1 0 42816 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_430
timestamp 1621261055
transform 1 0 42432 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_441
timestamp 1621261055
transform 1 0 43488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_438
timestamp 1621261055
transform 1 0 43200 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_446
timestamp 1621261055
transform 1 0 43968 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_438
timestamp 1621261055
transform 1 0 43200 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_759
timestamp 1621261055
transform 1 0 43392 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_449
timestamp 1621261055
transform 1 0 44256 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_454
timestamp 1621261055
transform 1 0 44736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_457
timestamp 1621261055
transform 1 0 45024 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_462
timestamp 1621261055
transform 1 0 45504 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_473
timestamp 1621261055
transform 1 0 46560 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_465
timestamp 1621261055
transform 1 0 45792 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_469
timestamp 1621261055
transform 1 0 46176 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_466
timestamp 1621261055
transform 1 0 45888 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_127
timestamp 1621261055
transform 1 0 46368 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_749
timestamp 1621261055
transform 1 0 46080 0 -1 39294
box -38 -49 134 715
use NAND3X1  NAND3X1
timestamp 1623610208
transform 1 0 46560 0 -1 39294
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_8  FILLER_55_481
timestamp 1621261055
transform 1 0 47328 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_485
timestamp 1621261055
transform 1 0 47712 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_493
timestamp 1621261055
transform 1 0 48480 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_489
timestamp 1621261055
transform 1 0 48096 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_493
timestamp 1621261055
transform 1 0 48480 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_760
timestamp 1621261055
transform 1 0 48672 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_496
timestamp 1621261055
transform 1 0 48768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_501
timestamp 1621261055
transform 1 0 49248 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_512
timestamp 1621261055
transform 1 0 50304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_504
timestamp 1621261055
transform 1 0 49536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_509
timestamp 1621261055
transform 1 0 50016 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_520
timestamp 1621261055
transform 1 0 51072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_521
timestamp 1621261055
transform 1 0 51168 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_517
timestamp 1621261055
transform 1 0 50784 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_528
timestamp 1621261055
transform 1 0 51840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_524
timestamp 1621261055
transform 1 0 51456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_750
timestamp 1621261055
transform 1 0 51360 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_536
timestamp 1621261055
transform 1 0 52608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_532
timestamp 1621261055
transform 1 0 52224 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_544
timestamp 1621261055
transform 1 0 53376 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_540
timestamp 1621261055
transform 1 0 52992 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_551
timestamp 1621261055
transform 1 0 54048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_548
timestamp 1621261055
transform 1 0 53760 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_548
timestamp 1621261055
transform 1 0 53760 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_761
timestamp 1621261055
transform 1 0 53952 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_559
timestamp 1621261055
transform 1 0 54816 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_556
timestamp 1621261055
transform 1 0 54528 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_567
timestamp 1621261055
transform 1 0 55584 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_564
timestamp 1621261055
transform 1 0 55296 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_575
timestamp 1621261055
transform 1 0 56352 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_576
timestamp 1621261055
transform 1 0 56448 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_572
timestamp 1621261055
transform 1 0 56064 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_751
timestamp 1621261055
transform 1 0 56640 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_583
timestamp 1621261055
transform 1 0 57120 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_587
timestamp 1621261055
transform 1 0 57504 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_579
timestamp 1621261055
transform 1 0 56736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_591
timestamp 1621261055
transform 1 0 57888 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_109
timestamp 1621261055
transform -1 0 58848 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_111
timestamp 1621261055
transform -1 0 58848 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_595
timestamp 1621261055
transform 1 0 58272 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_595
timestamp 1621261055
transform 1 0 58272 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_112
timestamp 1621261055
transform 1 0 1152 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_762
timestamp 1621261055
transform 1 0 3840 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_4
timestamp 1621261055
transform 1 0 1536 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_12
timestamp 1621261055
transform 1 0 2304 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_20
timestamp 1621261055
transform 1 0 3072 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_29
timestamp 1621261055
transform 1 0 3936 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_37
timestamp 1621261055
transform 1 0 4704 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_45
timestamp 1621261055
transform 1 0 5472 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_53
timestamp 1621261055
transform 1 0 6240 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_61
timestamp 1621261055
transform 1 0 7008 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_763
timestamp 1621261055
transform 1 0 9120 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_69
timestamp 1621261055
transform 1 0 7776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_77
timestamp 1621261055
transform 1 0 8544 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_81
timestamp 1621261055
transform 1 0 8928 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_84
timestamp 1621261055
transform 1 0 9216 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_92
timestamp 1621261055
transform 1 0 9984 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_100
timestamp 1621261055
transform 1 0 10752 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_108
timestamp 1621261055
transform 1 0 11520 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_116
timestamp 1621261055
transform 1 0 12288 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_124
timestamp 1621261055
transform 1 0 13056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_132
timestamp 1621261055
transform 1 0 13824 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _043_
timestamp 1621261055
transform 1 0 16512 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_764
timestamp 1621261055
transform 1 0 14400 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_136
timestamp 1621261055
transform 1 0 14208 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_139
timestamp 1621261055
transform 1 0 14496 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_147
timestamp 1621261055
transform 1 0 15264 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_155
timestamp 1621261055
transform 1 0 16032 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_56_159
timestamp 1621261055
transform 1 0 16416 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_163
timestamp 1621261055
transform 1 0 16800 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_765
timestamp 1621261055
transform 1 0 19680 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_171
timestamp 1621261055
transform 1 0 17568 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_179
timestamp 1621261055
transform 1 0 18336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_187
timestamp 1621261055
transform 1 0 19104 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_191
timestamp 1621261055
transform 1 0 19488 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_194
timestamp 1621261055
transform 1 0 19776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_202
timestamp 1621261055
transform 1 0 20544 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_210
timestamp 1621261055
transform 1 0 21312 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_218
timestamp 1621261055
transform 1 0 22080 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_226
timestamp 1621261055
transform 1 0 22848 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_766
timestamp 1621261055
transform 1 0 24960 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_234
timestamp 1621261055
transform 1 0 23616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_242
timestamp 1621261055
transform 1 0 24384 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_246
timestamp 1621261055
transform 1 0 24768 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_249
timestamp 1621261055
transform 1 0 25056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_257
timestamp 1621261055
transform 1 0 25824 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_265
timestamp 1621261055
transform 1 0 26592 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_273
timestamp 1621261055
transform 1 0 27360 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_281
timestamp 1621261055
transform 1 0 28128 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_289
timestamp 1621261055
transform 1 0 28896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_297
timestamp 1621261055
transform 1 0 29664 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_767
timestamp 1621261055
transform 1 0 30240 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_301
timestamp 1621261055
transform 1 0 30048 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_304
timestamp 1621261055
transform 1 0 30336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_312
timestamp 1621261055
transform 1 0 31104 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_320
timestamp 1621261055
transform 1 0 31872 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_328
timestamp 1621261055
transform 1 0 32640 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_768
timestamp 1621261055
transform 1 0 35520 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_336
timestamp 1621261055
transform 1 0 33408 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_344
timestamp 1621261055
transform 1 0 34176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_352
timestamp 1621261055
transform 1 0 34944 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_356
timestamp 1621261055
transform 1 0 35328 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_359
timestamp 1621261055
transform 1 0 35616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_367
timestamp 1621261055
transform 1 0 36384 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_375
timestamp 1621261055
transform 1 0 37152 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_383
timestamp 1621261055
transform 1 0 37920 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_391
timestamp 1621261055
transform 1 0 38688 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_769
timestamp 1621261055
transform 1 0 40800 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_399
timestamp 1621261055
transform 1 0 39456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_407
timestamp 1621261055
transform 1 0 40224 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_411
timestamp 1621261055
transform 1 0 40608 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_414
timestamp 1621261055
transform 1 0 40896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_422
timestamp 1621261055
transform 1 0 41664 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_430
timestamp 1621261055
transform 1 0 42432 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_438
timestamp 1621261055
transform 1 0 43200 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_446
timestamp 1621261055
transform 1 0 43968 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_454
timestamp 1621261055
transform 1 0 44736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_462
timestamp 1621261055
transform 1 0 45504 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_770
timestamp 1621261055
transform 1 0 46080 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_466
timestamp 1621261055
transform 1 0 45888 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_469
timestamp 1621261055
transform 1 0 46176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_477
timestamp 1621261055
transform 1 0 46944 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_485
timestamp 1621261055
transform 1 0 47712 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_493
timestamp 1621261055
transform 1 0 48480 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _018_
timestamp 1621261055
transform 1 0 49536 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _055_
timestamp 1621261055
transform 1 0 51840 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_771
timestamp 1621261055
transform 1 0 51360 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_501
timestamp 1621261055
transform 1 0 49248 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_503
timestamp 1621261055
transform 1 0 49440 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_507
timestamp 1621261055
transform 1 0 49824 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_515
timestamp 1621261055
transform 1 0 50592 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_524
timestamp 1621261055
transform 1 0 51456 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_56_531
timestamp 1621261055
transform 1 0 52128 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_539
timestamp 1621261055
transform 1 0 52896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_547
timestamp 1621261055
transform 1 0 53664 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_555
timestamp 1621261055
transform 1 0 54432 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_772
timestamp 1621261055
transform 1 0 56640 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_563
timestamp 1621261055
transform 1 0 55200 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_571
timestamp 1621261055
transform 1 0 55968 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_575
timestamp 1621261055
transform 1 0 56352 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_577
timestamp 1621261055
transform 1 0 56544 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_579
timestamp 1621261055
transform 1 0 56736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_587
timestamp 1621261055
transform 1 0 57504 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_113
timestamp 1621261055
transform -1 0 58848 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_595
timestamp 1621261055
transform 1 0 58272 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_114
timestamp 1621261055
transform 1 0 1152 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_57_4
timestamp 1621261055
transform 1 0 1536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_12
timestamp 1621261055
transform 1 0 2304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_20
timestamp 1621261055
transform 1 0 3072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_28
timestamp 1621261055
transform 1 0 3840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_773
timestamp 1621261055
transform 1 0 6432 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_36
timestamp 1621261055
transform 1 0 4608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_44
timestamp 1621261055
transform 1 0 5376 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_52
timestamp 1621261055
transform 1 0 6144 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_54
timestamp 1621261055
transform 1 0 6336 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_56
timestamp 1621261055
transform 1 0 6528 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_64
timestamp 1621261055
transform 1 0 7296 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_72
timestamp 1621261055
transform 1 0 8064 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_80
timestamp 1621261055
transform 1 0 8832 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_88
timestamp 1621261055
transform 1 0 9600 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_96
timestamp 1621261055
transform 1 0 10368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_774
timestamp 1621261055
transform 1 0 11712 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_104
timestamp 1621261055
transform 1 0 11136 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_108
timestamp 1621261055
transform 1 0 11520 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_111
timestamp 1621261055
transform 1 0 11808 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_119
timestamp 1621261055
transform 1 0 12576 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_127
timestamp 1621261055
transform 1 0 13344 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_775
timestamp 1621261055
transform 1 0 16992 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_135
timestamp 1621261055
transform 1 0 14112 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_143
timestamp 1621261055
transform 1 0 14880 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_151
timestamp 1621261055
transform 1 0 15648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_159
timestamp 1621261055
transform 1 0 16416 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_163
timestamp 1621261055
transform 1 0 16800 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_166
timestamp 1621261055
transform 1 0 17088 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_174
timestamp 1621261055
transform 1 0 17856 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_182
timestamp 1621261055
transform 1 0 18624 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_190
timestamp 1621261055
transform 1 0 19392 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_198
timestamp 1621261055
transform 1 0 20160 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _133_
timestamp 1621261055
transform 1 0 23136 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_776
timestamp 1621261055
transform 1 0 22272 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_168
timestamp 1621261055
transform 1 0 22944 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_206
timestamp 1621261055
transform 1 0 20928 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_214
timestamp 1621261055
transform 1 0 21696 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_218
timestamp 1621261055
transform 1 0 22080 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_57_221
timestamp 1621261055
transform 1 0 22368 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_225
timestamp 1621261055
transform 1 0 22752 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_232
timestamp 1621261055
transform 1 0 23424 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_240
timestamp 1621261055
transform 1 0 24192 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_248
timestamp 1621261055
transform 1 0 24960 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_256
timestamp 1621261055
transform 1 0 25728 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_264
timestamp 1621261055
transform 1 0 26496 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_777
timestamp 1621261055
transform 1 0 27552 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_272
timestamp 1621261055
transform 1 0 27264 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_274
timestamp 1621261055
transform 1 0 27456 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_276
timestamp 1621261055
transform 1 0 27648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_284
timestamp 1621261055
transform 1 0 28416 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_292
timestamp 1621261055
transform 1 0 29184 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _062_
timestamp 1621261055
transform 1 0 29952 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_778
timestamp 1621261055
transform 1 0 32832 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_303
timestamp 1621261055
transform 1 0 30240 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_311
timestamp 1621261055
transform 1 0 31008 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_319
timestamp 1621261055
transform 1 0 31776 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_327
timestamp 1621261055
transform 1 0 32544 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_329
timestamp 1621261055
transform 1 0 32736 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_331
timestamp 1621261055
transform 1 0 32928 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_339
timestamp 1621261055
transform 1 0 33696 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_347
timestamp 1621261055
transform 1 0 34464 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_355
timestamp 1621261055
transform 1 0 35232 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_363
timestamp 1621261055
transform 1 0 36000 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_779
timestamp 1621261055
transform 1 0 38112 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_371
timestamp 1621261055
transform 1 0 36768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_379
timestamp 1621261055
transform 1 0 37536 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_383
timestamp 1621261055
transform 1 0 37920 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_386
timestamp 1621261055
transform 1 0 38208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_394
timestamp 1621261055
transform 1 0 38976 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_402
timestamp 1621261055
transform 1 0 39744 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_410
timestamp 1621261055
transform 1 0 40512 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_418
timestamp 1621261055
transform 1 0 41280 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_426
timestamp 1621261055
transform 1 0 42048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _215_
timestamp 1621261055
transform 1 0 45504 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_780
timestamp 1621261055
transform 1 0 43392 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_434
timestamp 1621261055
transform 1 0 42816 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_438
timestamp 1621261055
transform 1 0 43200 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_441
timestamp 1621261055
transform 1 0 43488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_449
timestamp 1621261055
transform 1 0 44256 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_457
timestamp 1621261055
transform 1 0 45024 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_57_461
timestamp 1621261055
transform 1 0 45408 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_781
timestamp 1621261055
transform 1 0 48672 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_465
timestamp 1621261055
transform 1 0 45792 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_473
timestamp 1621261055
transform 1 0 46560 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_481
timestamp 1621261055
transform 1 0 47328 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_489
timestamp 1621261055
transform 1 0 48096 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_493
timestamp 1621261055
transform 1 0 48480 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_496
timestamp 1621261055
transform 1 0 48768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_504
timestamp 1621261055
transform 1 0 49536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_512
timestamp 1621261055
transform 1 0 50304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_520
timestamp 1621261055
transform 1 0 51072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_528
timestamp 1621261055
transform 1 0 51840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_782
timestamp 1621261055
transform 1 0 53952 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_536
timestamp 1621261055
transform 1 0 52608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_544
timestamp 1621261055
transform 1 0 53376 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_548
timestamp 1621261055
transform 1 0 53760 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_551
timestamp 1621261055
transform 1 0 54048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_559
timestamp 1621261055
transform 1 0 54816 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_567
timestamp 1621261055
transform 1 0 55584 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_575
timestamp 1621261055
transform 1 0 56352 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_583
timestamp 1621261055
transform 1 0 57120 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_591
timestamp 1621261055
transform 1 0 57888 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_115
timestamp 1621261055
transform -1 0 58848 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_595
timestamp 1621261055
transform 1 0 58272 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_116
timestamp 1621261055
transform 1 0 1152 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_783
timestamp 1621261055
transform 1 0 3840 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_4
timestamp 1621261055
transform 1 0 1536 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_12
timestamp 1621261055
transform 1 0 2304 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_20
timestamp 1621261055
transform 1 0 3072 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_29
timestamp 1621261055
transform 1 0 3936 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_37
timestamp 1621261055
transform 1 0 4704 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_45
timestamp 1621261055
transform 1 0 5472 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_53
timestamp 1621261055
transform 1 0 6240 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_61
timestamp 1621261055
transform 1 0 7008 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_784
timestamp 1621261055
transform 1 0 9120 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_69
timestamp 1621261055
transform 1 0 7776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_77
timestamp 1621261055
transform 1 0 8544 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_81
timestamp 1621261055
transform 1 0 8928 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_84
timestamp 1621261055
transform 1 0 9216 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_92
timestamp 1621261055
transform 1 0 9984 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_100
timestamp 1621261055
transform 1 0 10752 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_108
timestamp 1621261055
transform 1 0 11520 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_116
timestamp 1621261055
transform 1 0 12288 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_124
timestamp 1621261055
transform 1 0 13056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_132
timestamp 1621261055
transform 1 0 13824 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_785
timestamp 1621261055
transform 1 0 14400 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_136
timestamp 1621261055
transform 1 0 14208 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_139
timestamp 1621261055
transform 1 0 14496 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_147
timestamp 1621261055
transform 1 0 15264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_155
timestamp 1621261055
transform 1 0 16032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_163
timestamp 1621261055
transform 1 0 16800 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_786
timestamp 1621261055
transform 1 0 19680 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_171
timestamp 1621261055
transform 1 0 17568 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_179
timestamp 1621261055
transform 1 0 18336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_187
timestamp 1621261055
transform 1 0 19104 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_191
timestamp 1621261055
transform 1 0 19488 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_194
timestamp 1621261055
transform 1 0 19776 0 -1 41958
box -38 -49 806 715
use AND2X2  AND2X2
timestamp 1623610208
transform 1 0 21888 0 -1 41958
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_8  FILLER_58_202
timestamp 1621261055
transform 1 0 20544 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_210
timestamp 1621261055
transform 1 0 21312 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_214
timestamp 1621261055
transform 1 0 21696 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_228
timestamp 1621261055
transform 1 0 23040 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_787
timestamp 1621261055
transform 1 0 24960 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_236
timestamp 1621261055
transform 1 0 23808 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_244
timestamp 1621261055
transform 1 0 24576 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_58_249
timestamp 1621261055
transform 1 0 25056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_257
timestamp 1621261055
transform 1 0 25824 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_265
timestamp 1621261055
transform 1 0 26592 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_273
timestamp 1621261055
transform 1 0 27360 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_281
timestamp 1621261055
transform 1 0 28128 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_289
timestamp 1621261055
transform 1 0 28896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_297
timestamp 1621261055
transform 1 0 29664 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_788
timestamp 1621261055
transform 1 0 30240 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_301
timestamp 1621261055
transform 1 0 30048 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_304
timestamp 1621261055
transform 1 0 30336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_312
timestamp 1621261055
transform 1 0 31104 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_320
timestamp 1621261055
transform 1 0 31872 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_328
timestamp 1621261055
transform 1 0 32640 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_789
timestamp 1621261055
transform 1 0 35520 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_336
timestamp 1621261055
transform 1 0 33408 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_344
timestamp 1621261055
transform 1 0 34176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_352
timestamp 1621261055
transform 1 0 34944 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_356
timestamp 1621261055
transform 1 0 35328 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_359
timestamp 1621261055
transform 1 0 35616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_367
timestamp 1621261055
transform 1 0 36384 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_375
timestamp 1621261055
transform 1 0 37152 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_383
timestamp 1621261055
transform 1 0 37920 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_391
timestamp 1621261055
transform 1 0 38688 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_790
timestamp 1621261055
transform 1 0 40800 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_222
timestamp 1621261055
transform -1 0 42432 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_399
timestamp 1621261055
transform 1 0 39456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_407
timestamp 1621261055
transform 1 0 40224 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_411
timestamp 1621261055
transform 1 0 40608 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_414
timestamp 1621261055
transform 1 0 40896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_422
timestamp 1621261055
transform 1 0 41664 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_426
timestamp 1621261055
transform 1 0 42048 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _185_
timestamp 1621261055
transform -1 0 42720 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_58_433
timestamp 1621261055
transform 1 0 42720 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_441
timestamp 1621261055
transform 1 0 43488 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_449
timestamp 1621261055
transform 1 0 44256 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_457
timestamp 1621261055
transform 1 0 45024 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_791
timestamp 1621261055
transform 1 0 46080 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_465
timestamp 1621261055
transform 1 0 45792 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_467
timestamp 1621261055
transform 1 0 45984 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_469
timestamp 1621261055
transform 1 0 46176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_477
timestamp 1621261055
transform 1 0 46944 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_485
timestamp 1621261055
transform 1 0 47712 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_493
timestamp 1621261055
transform 1 0 48480 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_792
timestamp 1621261055
transform 1 0 51360 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_501
timestamp 1621261055
transform 1 0 49248 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_509
timestamp 1621261055
transform 1 0 50016 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_517
timestamp 1621261055
transform 1 0 50784 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_521
timestamp 1621261055
transform 1 0 51168 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_524
timestamp 1621261055
transform 1 0 51456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_532
timestamp 1621261055
transform 1 0 52224 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_540
timestamp 1621261055
transform 1 0 52992 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_548
timestamp 1621261055
transform 1 0 53760 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_556
timestamp 1621261055
transform 1 0 54528 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _190_
timestamp 1621261055
transform -1 0 57504 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_793
timestamp 1621261055
transform 1 0 56640 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_228
timestamp 1621261055
transform -1 0 57216 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_564
timestamp 1621261055
transform 1 0 55296 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_572
timestamp 1621261055
transform 1 0 56064 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_576
timestamp 1621261055
transform 1 0 56448 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_579
timestamp 1621261055
transform 1 0 56736 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_581
timestamp 1621261055
transform 1 0 56928 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_587
timestamp 1621261055
transform 1 0 57504 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_117
timestamp 1621261055
transform -1 0 58848 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_595
timestamp 1621261055
transform 1 0 58272 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_118
timestamp 1621261055
transform 1 0 1152 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_4
timestamp 1621261055
transform 1 0 1536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_12
timestamp 1621261055
transform 1 0 2304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_20
timestamp 1621261055
transform 1 0 3072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_28
timestamp 1621261055
transform 1 0 3840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_794
timestamp 1621261055
transform 1 0 6432 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_36
timestamp 1621261055
transform 1 0 4608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_44
timestamp 1621261055
transform 1 0 5376 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_52
timestamp 1621261055
transform 1 0 6144 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_54
timestamp 1621261055
transform 1 0 6336 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_56
timestamp 1621261055
transform 1 0 6528 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_64
timestamp 1621261055
transform 1 0 7296 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_72
timestamp 1621261055
transform 1 0 8064 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_80
timestamp 1621261055
transform 1 0 8832 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_88
timestamp 1621261055
transform 1 0 9600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_96
timestamp 1621261055
transform 1 0 10368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_795
timestamp 1621261055
transform 1 0 11712 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_104
timestamp 1621261055
transform 1 0 11136 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_108
timestamp 1621261055
transform 1 0 11520 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_111
timestamp 1621261055
transform 1 0 11808 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_119
timestamp 1621261055
transform 1 0 12576 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_127
timestamp 1621261055
transform 1 0 13344 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_796
timestamp 1621261055
transform 1 0 16992 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_135
timestamp 1621261055
transform 1 0 14112 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_143
timestamp 1621261055
transform 1 0 14880 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_151
timestamp 1621261055
transform 1 0 15648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_159
timestamp 1621261055
transform 1 0 16416 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_163
timestamp 1621261055
transform 1 0 16800 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_166
timestamp 1621261055
transform 1 0 17088 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_174
timestamp 1621261055
transform 1 0 17856 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_182
timestamp 1621261055
transform 1 0 18624 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_190
timestamp 1621261055
transform 1 0 19392 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_198
timestamp 1621261055
transform 1 0 20160 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_797
timestamp 1621261055
transform 1 0 22272 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_206
timestamp 1621261055
transform 1 0 20928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_214
timestamp 1621261055
transform 1 0 21696 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_218
timestamp 1621261055
transform 1 0 22080 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_221
timestamp 1621261055
transform 1 0 22368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_229
timestamp 1621261055
transform 1 0 23136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_237
timestamp 1621261055
transform 1 0 23904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_245
timestamp 1621261055
transform 1 0 24672 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_253
timestamp 1621261055
transform 1 0 25440 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_261
timestamp 1621261055
transform 1 0 26208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _006_
timestamp 1621261055
transform 1 0 28032 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_798
timestamp 1621261055
transform 1 0 27552 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_269
timestamp 1621261055
transform 1 0 26976 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_273
timestamp 1621261055
transform 1 0 27360 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_59_276
timestamp 1621261055
transform 1 0 27648 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_283
timestamp 1621261055
transform 1 0 28320 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_291
timestamp 1621261055
transform 1 0 29088 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _206_
timestamp 1621261055
transform -1 0 30432 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_799
timestamp 1621261055
transform 1 0 32832 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_210
timestamp 1621261055
transform -1 0 30144 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_299
timestamp 1621261055
transform 1 0 29856 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_305
timestamp 1621261055
transform 1 0 30432 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_313
timestamp 1621261055
transform 1 0 31200 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_321
timestamp 1621261055
transform 1 0 31968 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_59_329
timestamp 1621261055
transform 1 0 32736 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_331
timestamp 1621261055
transform 1 0 32928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_339
timestamp 1621261055
transform 1 0 33696 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_347
timestamp 1621261055
transform 1 0 34464 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_355
timestamp 1621261055
transform 1 0 35232 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_363
timestamp 1621261055
transform 1 0 36000 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_800
timestamp 1621261055
transform 1 0 38112 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_371
timestamp 1621261055
transform 1 0 36768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_379
timestamp 1621261055
transform 1 0 37536 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_383
timestamp 1621261055
transform 1 0 37920 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_386
timestamp 1621261055
transform 1 0 38208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_394
timestamp 1621261055
transform 1 0 38976 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_402
timestamp 1621261055
transform 1 0 39744 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_410
timestamp 1621261055
transform 1 0 40512 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_418
timestamp 1621261055
transform 1 0 41280 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_426
timestamp 1621261055
transform 1 0 42048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_801
timestamp 1621261055
transform 1 0 43392 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_434
timestamp 1621261055
transform 1 0 42816 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_438
timestamp 1621261055
transform 1 0 43200 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_441
timestamp 1621261055
transform 1 0 43488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_449
timestamp 1621261055
transform 1 0 44256 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_457
timestamp 1621261055
transform 1 0 45024 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_802
timestamp 1621261055
transform 1 0 48672 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_465
timestamp 1621261055
transform 1 0 45792 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_473
timestamp 1621261055
transform 1 0 46560 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_481
timestamp 1621261055
transform 1 0 47328 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_489
timestamp 1621261055
transform 1 0 48096 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_493
timestamp 1621261055
transform 1 0 48480 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_496
timestamp 1621261055
transform 1 0 48768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_504
timestamp 1621261055
transform 1 0 49536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_512
timestamp 1621261055
transform 1 0 50304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_520
timestamp 1621261055
transform 1 0 51072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_528
timestamp 1621261055
transform 1 0 51840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_803
timestamp 1621261055
transform 1 0 53952 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_172
timestamp 1621261055
transform -1 0 55104 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_536
timestamp 1621261055
transform 1 0 52608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_544
timestamp 1621261055
transform 1 0 53376 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_548
timestamp 1621261055
transform 1 0 53760 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_551
timestamp 1621261055
transform 1 0 54048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_59_559
timestamp 1621261055
transform 1 0 54816 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _135_
timestamp 1621261055
transform -1 0 55392 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_59_565
timestamp 1621261055
transform 1 0 55392 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_573
timestamp 1621261055
transform 1 0 56160 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_581
timestamp 1621261055
transform 1 0 56928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_589
timestamp 1621261055
transform 1 0 57696 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_119
timestamp 1621261055
transform -1 0 58848 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_120
timestamp 1621261055
transform 1 0 1152 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_804
timestamp 1621261055
transform 1 0 3840 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_4
timestamp 1621261055
transform 1 0 1536 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_12
timestamp 1621261055
transform 1 0 2304 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_20
timestamp 1621261055
transform 1 0 3072 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_29
timestamp 1621261055
transform 1 0 3936 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_37
timestamp 1621261055
transform 1 0 4704 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_45
timestamp 1621261055
transform 1 0 5472 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_53
timestamp 1621261055
transform 1 0 6240 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_61
timestamp 1621261055
transform 1 0 7008 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_805
timestamp 1621261055
transform 1 0 9120 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_69
timestamp 1621261055
transform 1 0 7776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_77
timestamp 1621261055
transform 1 0 8544 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_81
timestamp 1621261055
transform 1 0 8928 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_84
timestamp 1621261055
transform 1 0 9216 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_92
timestamp 1621261055
transform 1 0 9984 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_100
timestamp 1621261055
transform 1 0 10752 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_108
timestamp 1621261055
transform 1 0 11520 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_116
timestamp 1621261055
transform 1 0 12288 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_124
timestamp 1621261055
transform 1 0 13056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_132
timestamp 1621261055
transform 1 0 13824 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _123_
timestamp 1621261055
transform 1 0 14880 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_806
timestamp 1621261055
transform 1 0 14400 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_156
timestamp 1621261055
transform 1 0 14688 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_136
timestamp 1621261055
transform 1 0 14208 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_139
timestamp 1621261055
transform 1 0 14496 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_146
timestamp 1621261055
transform 1 0 15168 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_154
timestamp 1621261055
transform 1 0 15936 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_162
timestamp 1621261055
transform 1 0 16704 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_807
timestamp 1621261055
transform 1 0 19680 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_170
timestamp 1621261055
transform 1 0 17472 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_178
timestamp 1621261055
transform 1 0 18240 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_186
timestamp 1621261055
transform 1 0 19008 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_190
timestamp 1621261055
transform 1 0 19392 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_192
timestamp 1621261055
transform 1 0 19584 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_194
timestamp 1621261055
transform 1 0 19776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_202
timestamp 1621261055
transform 1 0 20544 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_210
timestamp 1621261055
transform 1 0 21312 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_218
timestamp 1621261055
transform 1 0 22080 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_226
timestamp 1621261055
transform 1 0 22848 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_808
timestamp 1621261055
transform 1 0 24960 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_234
timestamp 1621261055
transform 1 0 23616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_242
timestamp 1621261055
transform 1 0 24384 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_246
timestamp 1621261055
transform 1 0 24768 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_249
timestamp 1621261055
transform 1 0 25056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_257
timestamp 1621261055
transform 1 0 25824 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_265
timestamp 1621261055
transform 1 0 26592 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_273
timestamp 1621261055
transform 1 0 27360 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_281
timestamp 1621261055
transform 1 0 28128 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_289
timestamp 1621261055
transform 1 0 28896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_297
timestamp 1621261055
transform 1 0 29664 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_809
timestamp 1621261055
transform 1 0 30240 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_301
timestamp 1621261055
transform 1 0 30048 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_304
timestamp 1621261055
transform 1 0 30336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_312
timestamp 1621261055
transform 1 0 31104 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_320
timestamp 1621261055
transform 1 0 31872 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_328
timestamp 1621261055
transform 1 0 32640 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _208_
timestamp 1621261055
transform -1 0 35136 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_810
timestamp 1621261055
transform 1 0 35520 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_212
timestamp 1621261055
transform -1 0 34848 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_336
timestamp 1621261055
transform 1 0 33408 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_344
timestamp 1621261055
transform 1 0 34176 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_60_348
timestamp 1621261055
transform 1 0 34560 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_354
timestamp 1621261055
transform 1 0 35136 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_60_359
timestamp 1621261055
transform 1 0 35616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_367
timestamp 1621261055
transform 1 0 36384 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_375
timestamp 1621261055
transform 1 0 37152 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_383
timestamp 1621261055
transform 1 0 37920 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_391
timestamp 1621261055
transform 1 0 38688 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_811
timestamp 1621261055
transform 1 0 40800 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_399
timestamp 1621261055
transform 1 0 39456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_407
timestamp 1621261055
transform 1 0 40224 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_411
timestamp 1621261055
transform 1 0 40608 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_414
timestamp 1621261055
transform 1 0 40896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_422
timestamp 1621261055
transform 1 0 41664 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_430
timestamp 1621261055
transform 1 0 42432 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_438
timestamp 1621261055
transform 1 0 43200 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_446
timestamp 1621261055
transform 1 0 43968 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_454
timestamp 1621261055
transform 1 0 44736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_462
timestamp 1621261055
transform 1 0 45504 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_812
timestamp 1621261055
transform 1 0 46080 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_466
timestamp 1621261055
transform 1 0 45888 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_469
timestamp 1621261055
transform 1 0 46176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_477
timestamp 1621261055
transform 1 0 46944 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_485
timestamp 1621261055
transform 1 0 47712 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_493
timestamp 1621261055
transform 1 0 48480 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _058_
timestamp 1621261055
transform 1 0 50304 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_813
timestamp 1621261055
transform 1 0 51360 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_501
timestamp 1621261055
transform 1 0 49248 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_509
timestamp 1621261055
transform 1 0 50016 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_511
timestamp 1621261055
transform 1 0 50208 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_515
timestamp 1621261055
transform 1 0 50592 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_524
timestamp 1621261055
transform 1 0 51456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _111_
timestamp 1621261055
transform -1 0 52992 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_141
timestamp 1621261055
transform -1 0 52704 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_532
timestamp 1621261055
transform 1 0 52224 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_534
timestamp 1621261055
transform 1 0 52416 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_540
timestamp 1621261055
transform 1 0 52992 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_548
timestamp 1621261055
transform 1 0 53760 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_556
timestamp 1621261055
transform 1 0 54528 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_814
timestamp 1621261055
transform 1 0 56640 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_564
timestamp 1621261055
transform 1 0 55296 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_572
timestamp 1621261055
transform 1 0 56064 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_576
timestamp 1621261055
transform 1 0 56448 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_579
timestamp 1621261055
transform 1 0 56736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_587
timestamp 1621261055
transform 1 0 57504 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_121
timestamp 1621261055
transform -1 0 58848 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_595
timestamp 1621261055
transform 1 0 58272 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_4
timestamp 1621261055
transform 1 0 1536 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_4
timestamp 1621261055
transform 1 0 1536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_124
timestamp 1621261055
transform 1 0 1152 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_122
timestamp 1621261055
transform 1 0 1152 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_12
timestamp 1621261055
transform 1 0 2304 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_12
timestamp 1621261055
transform 1 0 2304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_20
timestamp 1621261055
transform 1 0 3072 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_20
timestamp 1621261055
transform 1 0 3072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_29
timestamp 1621261055
transform 1 0 3936 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_28
timestamp 1621261055
transform 1 0 3840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_825
timestamp 1621261055
transform 1 0 3840 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_37
timestamp 1621261055
transform 1 0 4704 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_36
timestamp 1621261055
transform 1 0 4608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_45
timestamp 1621261055
transform 1 0 5472 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_44
timestamp 1621261055
transform 1 0 5376 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_53
timestamp 1621261055
transform 1 0 6240 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_56
timestamp 1621261055
transform 1 0 6528 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_54
timestamp 1621261055
transform 1 0 6336 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_52
timestamp 1621261055
transform 1 0 6144 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_815
timestamp 1621261055
transform 1 0 6432 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_61
timestamp 1621261055
transform 1 0 7008 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_64
timestamp 1621261055
transform 1 0 7296 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_69
timestamp 1621261055
transform 1 0 7776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_72
timestamp 1621261055
transform 1 0 8064 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_81
timestamp 1621261055
transform 1 0 8928 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_77
timestamp 1621261055
transform 1 0 8544 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_80
timestamp 1621261055
transform 1 0 8832 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_826
timestamp 1621261055
transform 1 0 9120 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_92
timestamp 1621261055
transform 1 0 9984 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_84
timestamp 1621261055
transform 1 0 9216 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_88
timestamp 1621261055
transform 1 0 9600 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_96
timestamp 1621261055
transform 1 0 10368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_100
timestamp 1621261055
transform 1 0 10752 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_104
timestamp 1621261055
transform 1 0 11136 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_116
timestamp 1621261055
transform 1 0 12288 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_108
timestamp 1621261055
transform 1 0 11520 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_111
timestamp 1621261055
transform 1 0 11808 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_108
timestamp 1621261055
transform 1 0 11520 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_816
timestamp 1621261055
transform 1 0 11712 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_124
timestamp 1621261055
transform 1 0 13056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_119
timestamp 1621261055
transform 1 0 12576 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_132
timestamp 1621261055
transform 1 0 13824 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_127
timestamp 1621261055
transform 1 0 13344 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_139
timestamp 1621261055
transform 1 0 14496 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_136
timestamp 1621261055
transform 1 0 14208 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_135
timestamp 1621261055
transform 1 0 14112 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_827
timestamp 1621261055
transform 1 0 14400 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_147
timestamp 1621261055
transform 1 0 15264 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_143
timestamp 1621261055
transform 1 0 14880 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_155
timestamp 1621261055
transform 1 0 16032 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_151
timestamp 1621261055
transform 1 0 15648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_163
timestamp 1621261055
transform 1 0 16800 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_163
timestamp 1621261055
transform 1 0 16800 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_159
timestamp 1621261055
transform 1 0 16416 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_817
timestamp 1621261055
transform 1 0 16992 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_171
timestamp 1621261055
transform 1 0 17568 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_166
timestamp 1621261055
transform 1 0 17088 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_179
timestamp 1621261055
transform 1 0 18336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_182
timestamp 1621261055
transform 1 0 18624 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_174
timestamp 1621261055
transform 1 0 17856 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_191
timestamp 1621261055
transform 1 0 19488 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_187
timestamp 1621261055
transform 1 0 19104 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_190
timestamp 1621261055
transform 1 0 19392 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_194
timestamp 1621261055
transform 1 0 19776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_198
timestamp 1621261055
transform 1 0 20160 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_828
timestamp 1621261055
transform 1 0 19680 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_202
timestamp 1621261055
transform 1 0 20544 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_206
timestamp 1621261055
transform 1 0 20928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_210
timestamp 1621261055
transform 1 0 21312 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_214
timestamp 1621261055
transform 1 0 21696 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_218
timestamp 1621261055
transform 1 0 22080 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_221
timestamp 1621261055
transform 1 0 22368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_218
timestamp 1621261055
transform 1 0 22080 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_818
timestamp 1621261055
transform 1 0 22272 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_226
timestamp 1621261055
transform 1 0 22848 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_229
timestamp 1621261055
transform 1 0 23136 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_234
timestamp 1621261055
transform 1 0 23616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_237
timestamp 1621261055
transform 1 0 23904 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_246
timestamp 1621261055
transform 1 0 24768 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_242
timestamp 1621261055
transform 1 0 24384 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_245
timestamp 1621261055
transform 1 0 24672 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_829
timestamp 1621261055
transform 1 0 24960 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_257
timestamp 1621261055
transform 1 0 25824 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_249
timestamp 1621261055
transform 1 0 25056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_253
timestamp 1621261055
transform 1 0 25440 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_261
timestamp 1621261055
transform 1 0 26208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_265
timestamp 1621261055
transform 1 0 26592 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_61_269
timestamp 1621261055
transform 1 0 26976 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_84
timestamp 1621261055
transform 1 0 26976 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _168_
timestamp 1621261055
transform 1 0 27168 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_274
timestamp 1621261055
transform 1 0 27456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_280
timestamp 1621261055
transform 1 0 28032 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_276
timestamp 1621261055
transform 1 0 27648 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_273
timestamp 1621261055
transform 1 0 27360 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_119
timestamp 1621261055
transform -1 0 28320 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_819
timestamp 1621261055
transform 1 0 27552 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_290
timestamp 1621261055
transform 1 0 28992 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_282
timestamp 1621261055
transform 1 0 28224 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_286
timestamp 1621261055
transform 1 0 28608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _080_
timestamp 1621261055
transform -1 0 28608 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_61_294
timestamp 1621261055
transform 1 0 29376 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_304
timestamp 1621261055
transform 1 0 30336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_62_302
timestamp 1621261055
transform 1 0 30144 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_62_298
timestamp 1621261055
transform 1 0 29760 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_302
timestamp 1621261055
transform 1 0 30144 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_830
timestamp 1621261055
transform 1 0 30240 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_312
timestamp 1621261055
transform 1 0 31104 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_310
timestamp 1621261055
transform 1 0 30912 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_320
timestamp 1621261055
transform 1 0 31872 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_318
timestamp 1621261055
transform 1 0 31680 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_330
timestamp 1621261055
transform 1 0 32832 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_62_324
timestamp 1621261055
transform 1 0 32256 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_326
timestamp 1621261055
transform 1 0 32448 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_186
timestamp 1621261055
transform 1 0 32352 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_820
timestamp 1621261055
transform 1 0 32832 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _151_
timestamp 1621261055
transform 1 0 32544 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_338
timestamp 1621261055
transform 1 0 33600 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_62_332
timestamp 1621261055
transform 1 0 33024 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_331
timestamp 1621261055
transform 1 0 32928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_198
timestamp 1621261055
transform -1 0 33312 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _198_
timestamp 1621261055
transform -1 0 33600 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_346
timestamp 1621261055
transform 1 0 34368 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_347
timestamp 1621261055
transform 1 0 34464 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_339
timestamp 1621261055
transform 1 0 33696 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_354
timestamp 1621261055
transform 1 0 35136 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_62_348
timestamp 1621261055
transform 1 0 34560 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_355
timestamp 1621261055
transform 1 0 35232 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_208
timestamp 1621261055
transform -1 0 34848 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _204_
timestamp 1621261055
transform -1 0 35136 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_359
timestamp 1621261055
transform 1 0 35616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_363
timestamp 1621261055
transform 1 0 36000 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_831
timestamp 1621261055
transform 1 0 35520 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_367
timestamp 1621261055
transform 1 0 36384 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_371
timestamp 1621261055
transform 1 0 36768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_375
timestamp 1621261055
transform 1 0 37152 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_379
timestamp 1621261055
transform 1 0 37536 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_383
timestamp 1621261055
transform 1 0 37920 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_386
timestamp 1621261055
transform 1 0 38208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_383
timestamp 1621261055
transform 1 0 37920 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_821
timestamp 1621261055
transform 1 0 38112 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_391
timestamp 1621261055
transform 1 0 38688 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_394
timestamp 1621261055
transform 1 0 38976 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_399
timestamp 1621261055
transform 1 0 39456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_402
timestamp 1621261055
transform 1 0 39744 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_411
timestamp 1621261055
transform 1 0 40608 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_407
timestamp 1621261055
transform 1 0 40224 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_410
timestamp 1621261055
transform 1 0 40512 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_832
timestamp 1621261055
transform 1 0 40800 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_422
timestamp 1621261055
transform 1 0 41664 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_414
timestamp 1621261055
transform 1 0 40896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_418
timestamp 1621261055
transform 1 0 41280 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_426
timestamp 1621261055
transform 1 0 42048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_430
timestamp 1621261055
transform 1 0 42432 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_434
timestamp 1621261055
transform 1 0 42816 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_446
timestamp 1621261055
transform 1 0 43968 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_438
timestamp 1621261055
transform 1 0 43200 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_441
timestamp 1621261055
transform 1 0 43488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_438
timestamp 1621261055
transform 1 0 43200 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_822
timestamp 1621261055
transform 1 0 43392 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_62_454
timestamp 1621261055
transform 1 0 44736 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_449
timestamp 1621261055
transform 1 0 44256 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_62_460
timestamp 1621261055
transform 1 0 45312 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_458
timestamp 1621261055
transform 1 0 45120 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_457
timestamp 1621261055
transform 1 0 45024 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _037_
timestamp 1621261055
transform 1 0 45408 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_469
timestamp 1621261055
transform 1 0 46176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_464
timestamp 1621261055
transform 1 0 45696 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_470
timestamp 1621261055
transform 1 0 46272 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_91
timestamp 1621261055
transform 1 0 45792 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_833
timestamp 1621261055
transform 1 0 46080 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _174_
timestamp 1621261055
transform 1 0 45984 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_477
timestamp 1621261055
transform 1 0 46944 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_478
timestamp 1621261055
transform 1 0 47040 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_485
timestamp 1621261055
transform 1 0 47712 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_486
timestamp 1621261055
transform 1 0 47808 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_493
timestamp 1621261055
transform 1 0 48480 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_494
timestamp 1621261055
transform 1 0 48576 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_823
timestamp 1621261055
transform 1 0 48672 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_501
timestamp 1621261055
transform 1 0 49248 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_496
timestamp 1621261055
transform 1 0 48768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_509
timestamp 1621261055
transform 1 0 50016 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_512
timestamp 1621261055
transform 1 0 50304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_504
timestamp 1621261055
transform 1 0 49536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_521
timestamp 1621261055
transform 1 0 51168 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_517
timestamp 1621261055
transform 1 0 50784 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_520
timestamp 1621261055
transform 1 0 51072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_524
timestamp 1621261055
transform 1 0 51456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_528
timestamp 1621261055
transform 1 0 51840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_834
timestamp 1621261055
transform 1 0 51360 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_532
timestamp 1621261055
transform 1 0 52224 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_536
timestamp 1621261055
transform 1 0 52608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_540
timestamp 1621261055
transform 1 0 52992 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_544
timestamp 1621261055
transform 1 0 53376 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_548
timestamp 1621261055
transform 1 0 53760 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_551
timestamp 1621261055
transform 1 0 54048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_548
timestamp 1621261055
transform 1 0 53760 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_824
timestamp 1621261055
transform 1 0 53952 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_62_556
timestamp 1621261055
transform 1 0 54528 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_559
timestamp 1621261055
transform 1 0 54816 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_89
timestamp 1621261055
transform 1 0 54912 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_565
timestamp 1621261055
transform 1 0 55392 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_567
timestamp 1621261055
transform 1 0 55584 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _173_
timestamp 1621261055
transform 1 0 55104 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_62_577
timestamp 1621261055
transform 1 0 56544 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_62_573
timestamp 1621261055
transform 1 0 56160 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_575
timestamp 1621261055
transform 1 0 56352 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_835
timestamp 1621261055
transform 1 0 56640 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_587
timestamp 1621261055
transform 1 0 57504 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_579
timestamp 1621261055
transform 1 0 56736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_583
timestamp 1621261055
transform 1 0 57120 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_591
timestamp 1621261055
transform 1 0 57888 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_123
timestamp 1621261055
transform -1 0 58848 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_125
timestamp 1621261055
transform -1 0 58848 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_595
timestamp 1621261055
transform 1 0 58272 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_595
timestamp 1621261055
transform 1 0 58272 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_126
timestamp 1621261055
transform 1 0 1152 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_4
timestamp 1621261055
transform 1 0 1536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_12
timestamp 1621261055
transform 1 0 2304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_20
timestamp 1621261055
transform 1 0 3072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_28
timestamp 1621261055
transform 1 0 3840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_836
timestamp 1621261055
transform 1 0 6432 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_36
timestamp 1621261055
transform 1 0 4608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_44
timestamp 1621261055
transform 1 0 5376 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_52
timestamp 1621261055
transform 1 0 6144 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_54
timestamp 1621261055
transform 1 0 6336 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_56
timestamp 1621261055
transform 1 0 6528 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_64
timestamp 1621261055
transform 1 0 7296 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_72
timestamp 1621261055
transform 1 0 8064 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_80
timestamp 1621261055
transform 1 0 8832 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_88
timestamp 1621261055
transform 1 0 9600 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_96
timestamp 1621261055
transform 1 0 10368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_837
timestamp 1621261055
transform 1 0 11712 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_104
timestamp 1621261055
transform 1 0 11136 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_108
timestamp 1621261055
transform 1 0 11520 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_111
timestamp 1621261055
transform 1 0 11808 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_119
timestamp 1621261055
transform 1 0 12576 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_127
timestamp 1621261055
transform 1 0 13344 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_838
timestamp 1621261055
transform 1 0 16992 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_135
timestamp 1621261055
transform 1 0 14112 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_143
timestamp 1621261055
transform 1 0 14880 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_151
timestamp 1621261055
transform 1 0 15648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_159
timestamp 1621261055
transform 1 0 16416 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_163
timestamp 1621261055
transform 1 0 16800 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_166
timestamp 1621261055
transform 1 0 17088 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_174
timestamp 1621261055
transform 1 0 17856 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_182
timestamp 1621261055
transform 1 0 18624 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_190
timestamp 1621261055
transform 1 0 19392 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_198
timestamp 1621261055
transform 1 0 20160 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_839
timestamp 1621261055
transform 1 0 22272 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_206
timestamp 1621261055
transform 1 0 20928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_214
timestamp 1621261055
transform 1 0 21696 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_218
timestamp 1621261055
transform 1 0 22080 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_221
timestamp 1621261055
transform 1 0 22368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_229
timestamp 1621261055
transform 1 0 23136 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _137_
timestamp 1621261055
transform 1 0 26400 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_174
timestamp 1621261055
transform 1 0 26208 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_237
timestamp 1621261055
transform 1 0 23904 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_245
timestamp 1621261055
transform 1 0 24672 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_253
timestamp 1621261055
transform 1 0 25440 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_840
timestamp 1621261055
transform 1 0 27552 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_266
timestamp 1621261055
transform 1 0 26688 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_63_274
timestamp 1621261055
transform 1 0 27456 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_276
timestamp 1621261055
transform 1 0 27648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_284
timestamp 1621261055
transform 1 0 28416 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_292
timestamp 1621261055
transform 1 0 29184 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_841
timestamp 1621261055
transform 1 0 32832 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_300
timestamp 1621261055
transform 1 0 29952 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_308
timestamp 1621261055
transform 1 0 30720 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_316
timestamp 1621261055
transform 1 0 31488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_324
timestamp 1621261055
transform 1 0 32256 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_328
timestamp 1621261055
transform 1 0 32640 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_331
timestamp 1621261055
transform 1 0 32928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_339
timestamp 1621261055
transform 1 0 33696 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_347
timestamp 1621261055
transform 1 0 34464 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_355
timestamp 1621261055
transform 1 0 35232 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_363
timestamp 1621261055
transform 1 0 36000 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_842
timestamp 1621261055
transform 1 0 38112 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_371
timestamp 1621261055
transform 1 0 36768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_379
timestamp 1621261055
transform 1 0 37536 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_383
timestamp 1621261055
transform 1 0 37920 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_386
timestamp 1621261055
transform 1 0 38208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_394
timestamp 1621261055
transform 1 0 38976 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_402
timestamp 1621261055
transform 1 0 39744 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_410
timestamp 1621261055
transform 1 0 40512 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_418
timestamp 1621261055
transform 1 0 41280 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_426
timestamp 1621261055
transform 1 0 42048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_843
timestamp 1621261055
transform 1 0 43392 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_434
timestamp 1621261055
transform 1 0 42816 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_438
timestamp 1621261055
transform 1 0 43200 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_441
timestamp 1621261055
transform 1 0 43488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_449
timestamp 1621261055
transform 1 0 44256 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_457
timestamp 1621261055
transform 1 0 45024 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_844
timestamp 1621261055
transform 1 0 48672 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_465
timestamp 1621261055
transform 1 0 45792 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_473
timestamp 1621261055
transform 1 0 46560 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_481
timestamp 1621261055
transform 1 0 47328 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_489
timestamp 1621261055
transform 1 0 48096 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_493
timestamp 1621261055
transform 1 0 48480 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_496
timestamp 1621261055
transform 1 0 48768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_504
timestamp 1621261055
transform 1 0 49536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_512
timestamp 1621261055
transform 1 0 50304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_520
timestamp 1621261055
transform 1 0 51072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_528
timestamp 1621261055
transform 1 0 51840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_845
timestamp 1621261055
transform 1 0 53952 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_536
timestamp 1621261055
transform 1 0 52608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_544
timestamp 1621261055
transform 1 0 53376 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_548
timestamp 1621261055
transform 1 0 53760 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_551
timestamp 1621261055
transform 1 0 54048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_559
timestamp 1621261055
transform 1 0 54816 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_567
timestamp 1621261055
transform 1 0 55584 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_575
timestamp 1621261055
transform 1 0 56352 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_583
timestamp 1621261055
transform 1 0 57120 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_591
timestamp 1621261055
transform 1 0 57888 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_127
timestamp 1621261055
transform -1 0 58848 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_595
timestamp 1621261055
transform 1 0 58272 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_128
timestamp 1621261055
transform 1 0 1152 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_846
timestamp 1621261055
transform 1 0 3840 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_4
timestamp 1621261055
transform 1 0 1536 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_12
timestamp 1621261055
transform 1 0 2304 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_20
timestamp 1621261055
transform 1 0 3072 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_29
timestamp 1621261055
transform 1 0 3936 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_37
timestamp 1621261055
transform 1 0 4704 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_45
timestamp 1621261055
transform 1 0 5472 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_53
timestamp 1621261055
transform 1 0 6240 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_61
timestamp 1621261055
transform 1 0 7008 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_847
timestamp 1621261055
transform 1 0 9120 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_69
timestamp 1621261055
transform 1 0 7776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_77
timestamp 1621261055
transform 1 0 8544 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_81
timestamp 1621261055
transform 1 0 8928 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_84
timestamp 1621261055
transform 1 0 9216 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_92
timestamp 1621261055
transform 1 0 9984 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_100
timestamp 1621261055
transform 1 0 10752 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_108
timestamp 1621261055
transform 1 0 11520 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_116
timestamp 1621261055
transform 1 0 12288 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_124
timestamp 1621261055
transform 1 0 13056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_132
timestamp 1621261055
transform 1 0 13824 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_848
timestamp 1621261055
transform 1 0 14400 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_136
timestamp 1621261055
transform 1 0 14208 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_139
timestamp 1621261055
transform 1 0 14496 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_147
timestamp 1621261055
transform 1 0 15264 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_155
timestamp 1621261055
transform 1 0 16032 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_163
timestamp 1621261055
transform 1 0 16800 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_849
timestamp 1621261055
transform 1 0 19680 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_171
timestamp 1621261055
transform 1 0 17568 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_179
timestamp 1621261055
transform 1 0 18336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_187
timestamp 1621261055
transform 1 0 19104 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_191
timestamp 1621261055
transform 1 0 19488 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_194
timestamp 1621261055
transform 1 0 19776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_202
timestamp 1621261055
transform 1 0 20544 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_210
timestamp 1621261055
transform 1 0 21312 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_218
timestamp 1621261055
transform 1 0 22080 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_226
timestamp 1621261055
transform 1 0 22848 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_850
timestamp 1621261055
transform 1 0 24960 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_234
timestamp 1621261055
transform 1 0 23616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_242
timestamp 1621261055
transform 1 0 24384 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_246
timestamp 1621261055
transform 1 0 24768 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_249
timestamp 1621261055
transform 1 0 25056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_257
timestamp 1621261055
transform 1 0 25824 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _149_
timestamp 1621261055
transform 1 0 28032 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_184
timestamp 1621261055
transform 1 0 27840 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_265
timestamp 1621261055
transform 1 0 26592 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_273
timestamp 1621261055
transform 1 0 27360 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_64_277
timestamp 1621261055
transform 1 0 27744 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_283
timestamp 1621261055
transform 1 0 28320 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_291
timestamp 1621261055
transform 1 0 29088 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_851
timestamp 1621261055
transform 1 0 30240 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_299
timestamp 1621261055
transform 1 0 29856 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_64_304
timestamp 1621261055
transform 1 0 30336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_312
timestamp 1621261055
transform 1 0 31104 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_320
timestamp 1621261055
transform 1 0 31872 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_328
timestamp 1621261055
transform 1 0 32640 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_852
timestamp 1621261055
transform 1 0 35520 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_336
timestamp 1621261055
transform 1 0 33408 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_344
timestamp 1621261055
transform 1 0 34176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_352
timestamp 1621261055
transform 1 0 34944 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_356
timestamp 1621261055
transform 1 0 35328 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_359
timestamp 1621261055
transform 1 0 35616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _098_
timestamp 1621261055
transform -1 0 39360 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_135
timestamp 1621261055
transform -1 0 39072 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_367
timestamp 1621261055
transform 1 0 36384 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_375
timestamp 1621261055
transform 1 0 37152 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_383
timestamp 1621261055
transform 1 0 37920 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_391
timestamp 1621261055
transform 1 0 38688 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_853
timestamp 1621261055
transform 1 0 40800 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_398
timestamp 1621261055
transform 1 0 39360 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_406
timestamp 1621261055
transform 1 0 40128 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_410
timestamp 1621261055
transform 1 0 40512 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_412
timestamp 1621261055
transform 1 0 40704 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_414
timestamp 1621261055
transform 1 0 40896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_422
timestamp 1621261055
transform 1 0 41664 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_430
timestamp 1621261055
transform 1 0 42432 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_438
timestamp 1621261055
transform 1 0 43200 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_446
timestamp 1621261055
transform 1 0 43968 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_454
timestamp 1621261055
transform 1 0 44736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_462
timestamp 1621261055
transform 1 0 45504 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_854
timestamp 1621261055
transform 1 0 46080 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_466
timestamp 1621261055
transform 1 0 45888 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_469
timestamp 1621261055
transform 1 0 46176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_477
timestamp 1621261055
transform 1 0 46944 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_485
timestamp 1621261055
transform 1 0 47712 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_493
timestamp 1621261055
transform 1 0 48480 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _051_
timestamp 1621261055
transform 1 0 48864 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_855
timestamp 1621261055
transform 1 0 51360 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_500
timestamp 1621261055
transform 1 0 49152 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_508
timestamp 1621261055
transform 1 0 49920 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_516
timestamp 1621261055
transform 1 0 50688 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_520
timestamp 1621261055
transform 1 0 51072 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_522
timestamp 1621261055
transform 1 0 51264 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_524
timestamp 1621261055
transform 1 0 51456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_532
timestamp 1621261055
transform 1 0 52224 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_540
timestamp 1621261055
transform 1 0 52992 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_548
timestamp 1621261055
transform 1 0 53760 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_556
timestamp 1621261055
transform 1 0 54528 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_856
timestamp 1621261055
transform 1 0 56640 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_564
timestamp 1621261055
transform 1 0 55296 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_572
timestamp 1621261055
transform 1 0 56064 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_576
timestamp 1621261055
transform 1 0 56448 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_579
timestamp 1621261055
transform 1 0 56736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_587
timestamp 1621261055
transform 1 0 57504 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_129
timestamp 1621261055
transform -1 0 58848 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_595
timestamp 1621261055
transform 1 0 58272 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_130
timestamp 1621261055
transform 1 0 1152 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_4
timestamp 1621261055
transform 1 0 1536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_12
timestamp 1621261055
transform 1 0 2304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_20
timestamp 1621261055
transform 1 0 3072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_28
timestamp 1621261055
transform 1 0 3840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_857
timestamp 1621261055
transform 1 0 6432 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_36
timestamp 1621261055
transform 1 0 4608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_44
timestamp 1621261055
transform 1 0 5376 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_52
timestamp 1621261055
transform 1 0 6144 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_54
timestamp 1621261055
transform 1 0 6336 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_56
timestamp 1621261055
transform 1 0 6528 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_64
timestamp 1621261055
transform 1 0 7296 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_72
timestamp 1621261055
transform 1 0 8064 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_80
timestamp 1621261055
transform 1 0 8832 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_88
timestamp 1621261055
transform 1 0 9600 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_96
timestamp 1621261055
transform 1 0 10368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_104
timestamp 1621261055
transform 1 0 11136 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_115
timestamp 1621261055
transform 1 0 12192 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_65_111
timestamp 1621261055
transform 1 0 11808 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_108
timestamp 1621261055
transform 1 0 11520 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_858
timestamp 1621261055
transform 1 0 11712 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_123
timestamp 1621261055
transform 1 0 12960 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_65_117
timestamp 1621261055
transform 1 0 12384 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_216
timestamp 1621261055
transform 1 0 12480 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _211_
timestamp 1621261055
transform 1 0 12672 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_214
timestamp 1621261055
transform -1 0 13920 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _209_
timestamp 1621261055
transform -1 0 14208 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_859
timestamp 1621261055
transform 1 0 16992 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_136
timestamp 1621261055
transform 1 0 14208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_144
timestamp 1621261055
transform 1 0 14976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_152
timestamp 1621261055
transform 1 0 15744 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_160
timestamp 1621261055
transform 1 0 16512 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_65_164
timestamp 1621261055
transform 1 0 16896 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_166
timestamp 1621261055
transform 1 0 17088 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_174
timestamp 1621261055
transform 1 0 17856 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_182
timestamp 1621261055
transform 1 0 18624 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_190
timestamp 1621261055
transform 1 0 19392 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_198
timestamp 1621261055
transform 1 0 20160 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _130_
timestamp 1621261055
transform 1 0 23232 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_860
timestamp 1621261055
transform 1 0 22272 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_162
timestamp 1621261055
transform 1 0 23040 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_206
timestamp 1621261055
transform 1 0 20928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_214
timestamp 1621261055
transform 1 0 21696 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_218
timestamp 1621261055
transform 1 0 22080 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_65_221
timestamp 1621261055
transform 1 0 22368 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_225
timestamp 1621261055
transform 1 0 22752 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_227
timestamp 1621261055
transform 1 0 22944 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _102_
timestamp 1621261055
transform 1 0 26112 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_137
timestamp 1621261055
transform 1 0 25920 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_233
timestamp 1621261055
transform 1 0 23520 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_241
timestamp 1621261055
transform 1 0 24288 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_249
timestamp 1621261055
transform 1 0 25056 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_65_257
timestamp 1621261055
transform 1 0 25824 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_263
timestamp 1621261055
transform 1 0 26400 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_861
timestamp 1621261055
transform 1 0 27552 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_271
timestamp 1621261055
transform 1 0 27168 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_276
timestamp 1621261055
transform 1 0 27648 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_284
timestamp 1621261055
transform 1 0 28416 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_292
timestamp 1621261055
transform 1 0 29184 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_862
timestamp 1621261055
transform 1 0 32832 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_300
timestamp 1621261055
transform 1 0 29952 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_308
timestamp 1621261055
transform 1 0 30720 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_316
timestamp 1621261055
transform 1 0 31488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_324
timestamp 1621261055
transform 1 0 32256 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_328
timestamp 1621261055
transform 1 0 32640 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _002_
timestamp 1621261055
transform 1 0 35616 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_65_331
timestamp 1621261055
transform 1 0 32928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_339
timestamp 1621261055
transform 1 0 33696 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_347
timestamp 1621261055
transform 1 0 34464 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_355
timestamp 1621261055
transform 1 0 35232 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_362
timestamp 1621261055
transform 1 0 35904 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_863
timestamp 1621261055
transform 1 0 38112 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_370
timestamp 1621261055
transform 1 0 36672 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_378
timestamp 1621261055
transform 1 0 37440 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_382
timestamp 1621261055
transform 1 0 37824 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_384
timestamp 1621261055
transform 1 0 38016 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_386
timestamp 1621261055
transform 1 0 38208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_394
timestamp 1621261055
transform 1 0 38976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_402
timestamp 1621261055
transform 1 0 39744 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_410
timestamp 1621261055
transform 1 0 40512 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_418
timestamp 1621261055
transform 1 0 41280 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_426
timestamp 1621261055
transform 1 0 42048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_864
timestamp 1621261055
transform 1 0 43392 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_434
timestamp 1621261055
transform 1 0 42816 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_438
timestamp 1621261055
transform 1 0 43200 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_441
timestamp 1621261055
transform 1 0 43488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_449
timestamp 1621261055
transform 1 0 44256 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_457
timestamp 1621261055
transform 1 0 45024 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_865
timestamp 1621261055
transform 1 0 48672 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_465
timestamp 1621261055
transform 1 0 45792 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_473
timestamp 1621261055
transform 1 0 46560 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_481
timestamp 1621261055
transform 1 0 47328 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_489
timestamp 1621261055
transform 1 0 48096 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_493
timestamp 1621261055
transform 1 0 48480 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _012_
timestamp 1621261055
transform 1 0 50016 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _044_
timestamp 1621261055
transform 1 0 50688 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_65_496
timestamp 1621261055
transform 1 0 48768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_504
timestamp 1621261055
transform 1 0 49536 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_65_508
timestamp 1621261055
transform 1 0 49920 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_512
timestamp 1621261055
transform 1 0 50304 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_519
timestamp 1621261055
transform 1 0 50976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_527
timestamp 1621261055
transform 1 0 51744 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_866
timestamp 1621261055
transform 1 0 53952 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_535
timestamp 1621261055
transform 1 0 52512 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_543
timestamp 1621261055
transform 1 0 53280 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_547
timestamp 1621261055
transform 1 0 53664 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_549
timestamp 1621261055
transform 1 0 53856 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_551
timestamp 1621261055
transform 1 0 54048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_559
timestamp 1621261055
transform 1 0 54816 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_567
timestamp 1621261055
transform 1 0 55584 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_575
timestamp 1621261055
transform 1 0 56352 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_583
timestamp 1621261055
transform 1 0 57120 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_591
timestamp 1621261055
transform 1 0 57888 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_131
timestamp 1621261055
transform -1 0 58848 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_595
timestamp 1621261055
transform 1 0 58272 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_132
timestamp 1621261055
transform 1 0 1152 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_867
timestamp 1621261055
transform 1 0 3840 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_4
timestamp 1621261055
transform 1 0 1536 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_12
timestamp 1621261055
transform 1 0 2304 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_20
timestamp 1621261055
transform 1 0 3072 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_29
timestamp 1621261055
transform 1 0 3936 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_37
timestamp 1621261055
transform 1 0 4704 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_45
timestamp 1621261055
transform 1 0 5472 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_53
timestamp 1621261055
transform 1 0 6240 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_61
timestamp 1621261055
transform 1 0 7008 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_868
timestamp 1621261055
transform 1 0 9120 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_69
timestamp 1621261055
transform 1 0 7776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_77
timestamp 1621261055
transform 1 0 8544 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_81
timestamp 1621261055
transform 1 0 8928 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_84
timestamp 1621261055
transform 1 0 9216 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_92
timestamp 1621261055
transform 1 0 9984 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_100
timestamp 1621261055
transform 1 0 10752 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_108
timestamp 1621261055
transform 1 0 11520 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_116
timestamp 1621261055
transform 1 0 12288 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_124
timestamp 1621261055
transform 1 0 13056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_132
timestamp 1621261055
transform 1 0 13824 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_869
timestamp 1621261055
transform 1 0 14400 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_136
timestamp 1621261055
transform 1 0 14208 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_139
timestamp 1621261055
transform 1 0 14496 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_147
timestamp 1621261055
transform 1 0 15264 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_155
timestamp 1621261055
transform 1 0 16032 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_163
timestamp 1621261055
transform 1 0 16800 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_870
timestamp 1621261055
transform 1 0 19680 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_171
timestamp 1621261055
transform 1 0 17568 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_179
timestamp 1621261055
transform 1 0 18336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_187
timestamp 1621261055
transform 1 0 19104 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_191
timestamp 1621261055
transform 1 0 19488 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_194
timestamp 1621261055
transform 1 0 19776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_202
timestamp 1621261055
transform 1 0 20544 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_210
timestamp 1621261055
transform 1 0 21312 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_218
timestamp 1621261055
transform 1 0 22080 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_226
timestamp 1621261055
transform 1 0 22848 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_871
timestamp 1621261055
transform 1 0 24960 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_234
timestamp 1621261055
transform 1 0 23616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_242
timestamp 1621261055
transform 1 0 24384 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_246
timestamp 1621261055
transform 1 0 24768 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_249
timestamp 1621261055
transform 1 0 25056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_257
timestamp 1621261055
transform 1 0 25824 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_265
timestamp 1621261055
transform 1 0 26592 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_273
timestamp 1621261055
transform 1 0 27360 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_281
timestamp 1621261055
transform 1 0 28128 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_289
timestamp 1621261055
transform 1 0 28896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_297
timestamp 1621261055
transform 1 0 29664 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_872
timestamp 1621261055
transform 1 0 30240 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_301
timestamp 1621261055
transform 1 0 30048 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_304
timestamp 1621261055
transform 1 0 30336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_312
timestamp 1621261055
transform 1 0 31104 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_320
timestamp 1621261055
transform 1 0 31872 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_328
timestamp 1621261055
transform 1 0 32640 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_873
timestamp 1621261055
transform 1 0 35520 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_336
timestamp 1621261055
transform 1 0 33408 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_344
timestamp 1621261055
transform 1 0 34176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_352
timestamp 1621261055
transform 1 0 34944 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_356
timestamp 1621261055
transform 1 0 35328 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_359
timestamp 1621261055
transform 1 0 35616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_367
timestamp 1621261055
transform 1 0 36384 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_375
timestamp 1621261055
transform 1 0 37152 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_383
timestamp 1621261055
transform 1 0 37920 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_391
timestamp 1621261055
transform 1 0 38688 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_874
timestamp 1621261055
transform 1 0 40800 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_399
timestamp 1621261055
transform 1 0 39456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_407
timestamp 1621261055
transform 1 0 40224 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_411
timestamp 1621261055
transform 1 0 40608 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_414
timestamp 1621261055
transform 1 0 40896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_422
timestamp 1621261055
transform 1 0 41664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_430
timestamp 1621261055
transform 1 0 42432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_438
timestamp 1621261055
transform 1 0 43200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_446
timestamp 1621261055
transform 1 0 43968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_454
timestamp 1621261055
transform 1 0 44736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_462
timestamp 1621261055
transform 1 0 45504 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_875
timestamp 1621261055
transform 1 0 46080 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_466
timestamp 1621261055
transform 1 0 45888 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_469
timestamp 1621261055
transform 1 0 46176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_477
timestamp 1621261055
transform 1 0 46944 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_485
timestamp 1621261055
transform 1 0 47712 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_493
timestamp 1621261055
transform 1 0 48480 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _131_
timestamp 1621261055
transform -1 0 52128 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_876
timestamp 1621261055
transform 1 0 51360 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_164
timestamp 1621261055
transform -1 0 51840 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_501
timestamp 1621261055
transform 1 0 49248 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_509
timestamp 1621261055
transform 1 0 50016 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_517
timestamp 1621261055
transform 1 0 50784 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_521
timestamp 1621261055
transform 1 0 51168 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_524
timestamp 1621261055
transform 1 0 51456 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_531
timestamp 1621261055
transform 1 0 52128 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_539
timestamp 1621261055
transform 1 0 52896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_547
timestamp 1621261055
transform 1 0 53664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_555
timestamp 1621261055
transform 1 0 54432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_877
timestamp 1621261055
transform 1 0 56640 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_563
timestamp 1621261055
transform 1 0 55200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_571
timestamp 1621261055
transform 1 0 55968 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_575
timestamp 1621261055
transform 1 0 56352 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_66_577
timestamp 1621261055
transform 1 0 56544 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_579
timestamp 1621261055
transform 1 0 56736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_587
timestamp 1621261055
transform 1 0 57504 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_133
timestamp 1621261055
transform -1 0 58848 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_595
timestamp 1621261055
transform 1 0 58272 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_134
timestamp 1621261055
transform 1 0 1152 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_4
timestamp 1621261055
transform 1 0 1536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_12
timestamp 1621261055
transform 1 0 2304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_20
timestamp 1621261055
transform 1 0 3072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_28
timestamp 1621261055
transform 1 0 3840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_878
timestamp 1621261055
transform 1 0 6432 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_36
timestamp 1621261055
transform 1 0 4608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_44
timestamp 1621261055
transform 1 0 5376 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_52
timestamp 1621261055
transform 1 0 6144 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_54
timestamp 1621261055
transform 1 0 6336 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_56
timestamp 1621261055
transform 1 0 6528 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_64
timestamp 1621261055
transform 1 0 7296 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_72
timestamp 1621261055
transform 1 0 8064 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_80
timestamp 1621261055
transform 1 0 8832 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_88
timestamp 1621261055
transform 1 0 9600 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_96
timestamp 1621261055
transform 1 0 10368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_879
timestamp 1621261055
transform 1 0 11712 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_104
timestamp 1621261055
transform 1 0 11136 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_108
timestamp 1621261055
transform 1 0 11520 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_111
timestamp 1621261055
transform 1 0 11808 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_119
timestamp 1621261055
transform 1 0 12576 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_127
timestamp 1621261055
transform 1 0 13344 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_880
timestamp 1621261055
transform 1 0 16992 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_135
timestamp 1621261055
transform 1 0 14112 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_143
timestamp 1621261055
transform 1 0 14880 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_151
timestamp 1621261055
transform 1 0 15648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_159
timestamp 1621261055
transform 1 0 16416 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_163
timestamp 1621261055
transform 1 0 16800 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_166
timestamp 1621261055
transform 1 0 17088 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_174
timestamp 1621261055
transform 1 0 17856 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_182
timestamp 1621261055
transform 1 0 18624 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_190
timestamp 1621261055
transform 1 0 19392 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_198
timestamp 1621261055
transform 1 0 20160 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_881
timestamp 1621261055
transform 1 0 22272 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_206
timestamp 1621261055
transform 1 0 20928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_214
timestamp 1621261055
transform 1 0 21696 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_218
timestamp 1621261055
transform 1 0 22080 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_221
timestamp 1621261055
transform 1 0 22368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_229
timestamp 1621261055
transform 1 0 23136 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_237
timestamp 1621261055
transform 1 0 23904 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_245
timestamp 1621261055
transform 1 0 24672 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_253
timestamp 1621261055
transform 1 0 25440 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_261
timestamp 1621261055
transform 1 0 26208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_882
timestamp 1621261055
transform 1 0 27552 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_269
timestamp 1621261055
transform 1 0 26976 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_273
timestamp 1621261055
transform 1 0 27360 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_276
timestamp 1621261055
transform 1 0 27648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_284
timestamp 1621261055
transform 1 0 28416 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_292
timestamp 1621261055
transform 1 0 29184 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _094_
timestamp 1621261055
transform -1 0 32448 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_883
timestamp 1621261055
transform 1 0 32832 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_131
timestamp 1621261055
transform -1 0 32160 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_300
timestamp 1621261055
transform 1 0 29952 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_308
timestamp 1621261055
transform 1 0 30720 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_316
timestamp 1621261055
transform 1 0 31488 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_67_320
timestamp 1621261055
transform 1 0 31872 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_326
timestamp 1621261055
transform 1 0 32448 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_331
timestamp 1621261055
transform 1 0 32928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_339
timestamp 1621261055
transform 1 0 33696 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_347
timestamp 1621261055
transform 1 0 34464 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_355
timestamp 1621261055
transform 1 0 35232 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_363
timestamp 1621261055
transform 1 0 36000 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_884
timestamp 1621261055
transform 1 0 38112 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_371
timestamp 1621261055
transform 1 0 36768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_379
timestamp 1621261055
transform 1 0 37536 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_383
timestamp 1621261055
transform 1 0 37920 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_386
timestamp 1621261055
transform 1 0 38208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_394
timestamp 1621261055
transform 1 0 38976 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_402
timestamp 1621261055
transform 1 0 39744 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_410
timestamp 1621261055
transform 1 0 40512 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_418
timestamp 1621261055
transform 1 0 41280 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_426
timestamp 1621261055
transform 1 0 42048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_885
timestamp 1621261055
transform 1 0 43392 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_434
timestamp 1621261055
transform 1 0 42816 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_438
timestamp 1621261055
transform 1 0 43200 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_441
timestamp 1621261055
transform 1 0 43488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_449
timestamp 1621261055
transform 1 0 44256 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_457
timestamp 1621261055
transform 1 0 45024 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_886
timestamp 1621261055
transform 1 0 48672 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_465
timestamp 1621261055
transform 1 0 45792 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_473
timestamp 1621261055
transform 1 0 46560 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_481
timestamp 1621261055
transform 1 0 47328 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_489
timestamp 1621261055
transform 1 0 48096 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_493
timestamp 1621261055
transform 1 0 48480 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_496
timestamp 1621261055
transform 1 0 48768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_504
timestamp 1621261055
transform 1 0 49536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_512
timestamp 1621261055
transform 1 0 50304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_520
timestamp 1621261055
transform 1 0 51072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_528
timestamp 1621261055
transform 1 0 51840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_887
timestamp 1621261055
transform 1 0 53952 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_536
timestamp 1621261055
transform 1 0 52608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_544
timestamp 1621261055
transform 1 0 53376 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_548
timestamp 1621261055
transform 1 0 53760 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_551
timestamp 1621261055
transform 1 0 54048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_559
timestamp 1621261055
transform 1 0 54816 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_567
timestamp 1621261055
transform 1 0 55584 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_575
timestamp 1621261055
transform 1 0 56352 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_583
timestamp 1621261055
transform 1 0 57120 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_591
timestamp 1621261055
transform 1 0 57888 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_135
timestamp 1621261055
transform -1 0 58848 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_595
timestamp 1621261055
transform 1 0 58272 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_136
timestamp 1621261055
transform 1 0 1152 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_888
timestamp 1621261055
transform 1 0 3840 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_4
timestamp 1621261055
transform 1 0 1536 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_12
timestamp 1621261055
transform 1 0 2304 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_20
timestamp 1621261055
transform 1 0 3072 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_29
timestamp 1621261055
transform 1 0 3936 0 -1 48618
box -38 -49 806 715
use AND2X1  AND2X1
timestamp 1623610208
transform 1 0 5280 0 -1 48618
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_4  FILLER_68_37
timestamp 1621261055
transform 1 0 4704 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_41
timestamp 1621261055
transform 1 0 5088 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_55
timestamp 1621261055
transform 1 0 6432 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_63
timestamp 1621261055
transform 1 0 7200 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_889
timestamp 1621261055
transform 1 0 9120 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_71
timestamp 1621261055
transform 1 0 7968 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_79
timestamp 1621261055
transform 1 0 8736 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_84
timestamp 1621261055
transform 1 0 9216 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_92
timestamp 1621261055
transform 1 0 9984 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_100
timestamp 1621261055
transform 1 0 10752 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_108
timestamp 1621261055
transform 1 0 11520 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_116
timestamp 1621261055
transform 1 0 12288 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_124
timestamp 1621261055
transform 1 0 13056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_132
timestamp 1621261055
transform 1 0 13824 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_890
timestamp 1621261055
transform 1 0 14400 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_136
timestamp 1621261055
transform 1 0 14208 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_139
timestamp 1621261055
transform 1 0 14496 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_147
timestamp 1621261055
transform 1 0 15264 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_155
timestamp 1621261055
transform 1 0 16032 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_163
timestamp 1621261055
transform 1 0 16800 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_891
timestamp 1621261055
transform 1 0 19680 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_171
timestamp 1621261055
transform 1 0 17568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_179
timestamp 1621261055
transform 1 0 18336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_187
timestamp 1621261055
transform 1 0 19104 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_191
timestamp 1621261055
transform 1 0 19488 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_194
timestamp 1621261055
transform 1 0 19776 0 -1 48618
box -38 -49 806 715
use BUFX2  BUFX2
timestamp 1623610208
transform 1 0 21696 0 -1 48618
box 0 -48 864 714
use sky130_fd_sc_ls__decap_8  FILLER_68_202
timestamp 1621261055
transform 1 0 20544 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_210
timestamp 1621261055
transform 1 0 21312 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_223
timestamp 1621261055
transform 1 0 22560 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_231
timestamp 1621261055
transform 1 0 23328 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_892
timestamp 1621261055
transform 1 0 24960 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_239
timestamp 1621261055
transform 1 0 24096 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_68_247
timestamp 1621261055
transform 1 0 24864 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_249
timestamp 1621261055
transform 1 0 25056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_257
timestamp 1621261055
transform 1 0 25824 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_265
timestamp 1621261055
transform 1 0 26592 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_273
timestamp 1621261055
transform 1 0 27360 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_281
timestamp 1621261055
transform 1 0 28128 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_289
timestamp 1621261055
transform 1 0 28896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_297
timestamp 1621261055
transform 1 0 29664 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_893
timestamp 1621261055
transform 1 0 30240 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_301
timestamp 1621261055
transform 1 0 30048 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_304
timestamp 1621261055
transform 1 0 30336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_312
timestamp 1621261055
transform 1 0 31104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_320
timestamp 1621261055
transform 1 0 31872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_328
timestamp 1621261055
transform 1 0 32640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_894
timestamp 1621261055
transform 1 0 35520 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_336
timestamp 1621261055
transform 1 0 33408 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_344
timestamp 1621261055
transform 1 0 34176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_352
timestamp 1621261055
transform 1 0 34944 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_356
timestamp 1621261055
transform 1 0 35328 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_359
timestamp 1621261055
transform 1 0 35616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_367
timestamp 1621261055
transform 1 0 36384 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_375
timestamp 1621261055
transform 1 0 37152 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_383
timestamp 1621261055
transform 1 0 37920 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_391
timestamp 1621261055
transform 1 0 38688 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_895
timestamp 1621261055
transform 1 0 40800 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_399
timestamp 1621261055
transform 1 0 39456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_407
timestamp 1621261055
transform 1 0 40224 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_411
timestamp 1621261055
transform 1 0 40608 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_414
timestamp 1621261055
transform 1 0 40896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_422
timestamp 1621261055
transform 1 0 41664 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_430
timestamp 1621261055
transform 1 0 42432 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_438
timestamp 1621261055
transform 1 0 43200 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_446
timestamp 1621261055
transform 1 0 43968 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_454
timestamp 1621261055
transform 1 0 44736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_462
timestamp 1621261055
transform 1 0 45504 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_896
timestamp 1621261055
transform 1 0 46080 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_466
timestamp 1621261055
transform 1 0 45888 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_469
timestamp 1621261055
transform 1 0 46176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_477
timestamp 1621261055
transform 1 0 46944 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_485
timestamp 1621261055
transform 1 0 47712 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_493
timestamp 1621261055
transform 1 0 48480 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_897
timestamp 1621261055
transform 1 0 51360 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_501
timestamp 1621261055
transform 1 0 49248 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_509
timestamp 1621261055
transform 1 0 50016 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_517
timestamp 1621261055
transform 1 0 50784 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_521
timestamp 1621261055
transform 1 0 51168 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_524
timestamp 1621261055
transform 1 0 51456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_532
timestamp 1621261055
transform 1 0 52224 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_540
timestamp 1621261055
transform 1 0 52992 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_548
timestamp 1621261055
transform 1 0 53760 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_556
timestamp 1621261055
transform 1 0 54528 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_898
timestamp 1621261055
transform 1 0 56640 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_564
timestamp 1621261055
transform 1 0 55296 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_572
timestamp 1621261055
transform 1 0 56064 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_576
timestamp 1621261055
transform 1 0 56448 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_579
timestamp 1621261055
transform 1 0 56736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_587
timestamp 1621261055
transform 1 0 57504 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_137
timestamp 1621261055
transform -1 0 58848 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_595
timestamp 1621261055
transform 1 0 58272 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_4
timestamp 1621261055
transform 1 0 1536 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_4
timestamp 1621261055
transform 1 0 1536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_140
timestamp 1621261055
transform 1 0 1152 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_138
timestamp 1621261055
transform 1 0 1152 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_12
timestamp 1621261055
transform 1 0 2304 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_12
timestamp 1621261055
transform 1 0 2304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_20
timestamp 1621261055
transform 1 0 3072 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_20
timestamp 1621261055
transform 1 0 3072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_29
timestamp 1621261055
transform 1 0 3936 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_28
timestamp 1621261055
transform 1 0 3840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_909
timestamp 1621261055
transform 1 0 3840 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_37
timestamp 1621261055
transform 1 0 4704 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_36
timestamp 1621261055
transform 1 0 4608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_45
timestamp 1621261055
transform 1 0 5472 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_44
timestamp 1621261055
transform 1 0 5376 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_53
timestamp 1621261055
transform 1 0 6240 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_56
timestamp 1621261055
transform 1 0 6528 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_69_54
timestamp 1621261055
transform 1 0 6336 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_52
timestamp 1621261055
transform 1 0 6144 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_218
timestamp 1621261055
transform -1 0 6912 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_899
timestamp 1621261055
transform 1 0 6432 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_61
timestamp 1621261055
transform 1 0 7008 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_63
timestamp 1621261055
transform 1 0 7200 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _184_
timestamp 1621261055
transform -1 0 7200 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_69
timestamp 1621261055
transform 1 0 7776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_71
timestamp 1621261055
transform 1 0 7968 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_81
timestamp 1621261055
transform 1 0 8928 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_77
timestamp 1621261055
transform 1 0 8544 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_79
timestamp 1621261055
transform 1 0 8736 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_910
timestamp 1621261055
transform 1 0 9120 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_92
timestamp 1621261055
transform 1 0 9984 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_84
timestamp 1621261055
transform 1 0 9216 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_87
timestamp 1621261055
transform 1 0 9504 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_95
timestamp 1621261055
transform 1 0 10272 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_100
timestamp 1621261055
transform 1 0 10752 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_107
timestamp 1621261055
transform 1 0 11424 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_103
timestamp 1621261055
transform 1 0 11040 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_70_114
timestamp 1621261055
transform 1 0 12096 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_112
timestamp 1621261055
transform 1 0 11904 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_108
timestamp 1621261055
transform 1 0 11520 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_111
timestamp 1621261055
transform 1 0 11808 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_109
timestamp 1621261055
transform 1 0 11616 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_194
timestamp 1621261055
transform -1 0 12384 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_900
timestamp 1621261055
transform 1 0 11712 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_120
timestamp 1621261055
transform 1 0 12672 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_123
timestamp 1621261055
transform 1 0 12960 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_119
timestamp 1621261055
transform 1 0 12576 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _194_
timestamp 1621261055
transform -1 0 12672 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _010_
timestamp 1621261055
transform 1 0 12672 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_128
timestamp 1621261055
transform 1 0 13440 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_131
timestamp 1621261055
transform 1 0 13728 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_139
timestamp 1621261055
transform 1 0 14496 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_136
timestamp 1621261055
transform 1 0 14208 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_139
timestamp 1621261055
transform 1 0 14496 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_911
timestamp 1621261055
transform 1 0 14400 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_147
timestamp 1621261055
transform 1 0 15264 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_147
timestamp 1621261055
transform 1 0 15264 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_155
timestamp 1621261055
transform 1 0 16032 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_155
timestamp 1621261055
transform 1 0 16032 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_163
timestamp 1621261055
transform 1 0 16800 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_163
timestamp 1621261055
transform 1 0 16800 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_901
timestamp 1621261055
transform 1 0 16992 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_171
timestamp 1621261055
transform 1 0 17568 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_166
timestamp 1621261055
transform 1 0 17088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_179
timestamp 1621261055
transform 1 0 18336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_182
timestamp 1621261055
transform 1 0 18624 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_174
timestamp 1621261055
transform 1 0 17856 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_191
timestamp 1621261055
transform 1 0 19488 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_187
timestamp 1621261055
transform 1 0 19104 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_190
timestamp 1621261055
transform 1 0 19392 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_194
timestamp 1621261055
transform 1 0 19776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_198
timestamp 1621261055
transform 1 0 20160 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_912
timestamp 1621261055
transform 1 0 19680 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_202
timestamp 1621261055
transform 1 0 20544 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_206
timestamp 1621261055
transform 1 0 20928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_210
timestamp 1621261055
transform 1 0 21312 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_214
timestamp 1621261055
transform 1 0 21696 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_218
timestamp 1621261055
transform 1 0 22080 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_221
timestamp 1621261055
transform 1 0 22368 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_218
timestamp 1621261055
transform 1 0 22080 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_902
timestamp 1621261055
transform 1 0 22272 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_70_226
timestamp 1621261055
transform 1 0 22848 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_230
timestamp 1621261055
transform 1 0 23232 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_225
timestamp 1621261055
transform 1 0 22752 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_226
timestamp 1621261055
transform -1 0 23136 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _189_
timestamp 1621261055
transform -1 0 23424 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _025_
timestamp 1621261055
transform 1 0 22944 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_240
timestamp 1621261055
transform 1 0 24192 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_232
timestamp 1621261055
transform 1 0 23424 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_238
timestamp 1621261055
transform 1 0 24000 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_249
timestamp 1621261055
transform 1 0 25056 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_246
timestamp 1621261055
transform 1 0 24768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_913
timestamp 1621261055
transform 1 0 24960 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_254
timestamp 1621261055
transform 1 0 25536 0 1 48618
box -38 -49 806 715
use NAND2X1  NAND2X1
timestamp 1623610208
transform 1 0 25440 0 -1 49950
box 0 -48 864 714
use sky130_fd_sc_ls__decap_4  FILLER_70_262
timestamp 1621261055
transform 1 0 26304 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_262
timestamp 1621261055
transform 1 0 26304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_269
timestamp 1621261055
transform 1 0 26976 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_270
timestamp 1621261055
transform 1 0 27072 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _009_
timestamp 1621261055
transform 1 0 26688 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_277
timestamp 1621261055
transform 1 0 27744 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_276
timestamp 1621261055
transform 1 0 27648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_274
timestamp 1621261055
transform 1 0 27456 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_903
timestamp 1621261055
transform 1 0 27552 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_285
timestamp 1621261055
transform 1 0 28512 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_284
timestamp 1621261055
transform 1 0 28416 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_293
timestamp 1621261055
transform 1 0 29280 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_292
timestamp 1621261055
transform 1 0 29184 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_304
timestamp 1621261055
transform 1 0 30336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_301
timestamp 1621261055
transform 1 0 30048 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_300
timestamp 1621261055
transform 1 0 29952 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_914
timestamp 1621261055
transform 1 0 30240 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_312
timestamp 1621261055
transform 1 0 31104 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_308
timestamp 1621261055
transform 1 0 30720 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_316
timestamp 1621261055
transform 1 0 31488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_115
timestamp 1621261055
transform -1 0 32064 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _076_
timestamp 1621261055
transform -1 0 32352 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_325
timestamp 1621261055
transform 1 0 32352 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_328
timestamp 1621261055
transform 1 0 32640 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_324
timestamp 1621261055
transform 1 0 32256 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_904
timestamp 1621261055
transform 1 0 32832 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_333
timestamp 1621261055
transform 1 0 33120 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_331
timestamp 1621261055
transform 1 0 32928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_341
timestamp 1621261055
transform 1 0 33888 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_347
timestamp 1621261055
transform 1 0 34464 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_339
timestamp 1621261055
transform 1 0 33696 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_349
timestamp 1621261055
transform 1 0 34656 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_355
timestamp 1621261055
transform 1 0 35232 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_359
timestamp 1621261055
transform 1 0 35616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_70_357
timestamp 1621261055
transform 1 0 35424 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_363
timestamp 1621261055
transform 1 0 36000 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_915
timestamp 1621261055
transform 1 0 35520 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_367
timestamp 1621261055
transform 1 0 36384 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_371
timestamp 1621261055
transform 1 0 36768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_375
timestamp 1621261055
transform 1 0 37152 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_379
timestamp 1621261055
transform 1 0 37536 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_383
timestamp 1621261055
transform 1 0 37920 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_386
timestamp 1621261055
transform 1 0 38208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_383
timestamp 1621261055
transform 1 0 37920 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_905
timestamp 1621261055
transform 1 0 38112 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_391
timestamp 1621261055
transform 1 0 38688 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_394
timestamp 1621261055
transform 1 0 38976 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_399
timestamp 1621261055
transform 1 0 39456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_402
timestamp 1621261055
transform 1 0 39744 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_411
timestamp 1621261055
transform 1 0 40608 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_407
timestamp 1621261055
transform 1 0 40224 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_410
timestamp 1621261055
transform 1 0 40512 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_916
timestamp 1621261055
transform 1 0 40800 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_422
timestamp 1621261055
transform 1 0 41664 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_414
timestamp 1621261055
transform 1 0 40896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_418
timestamp 1621261055
transform 1 0 41280 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_426
timestamp 1621261055
transform 1 0 42048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_430
timestamp 1621261055
transform 1 0 42432 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_434
timestamp 1621261055
transform 1 0 42816 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_446
timestamp 1621261055
transform 1 0 43968 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_438
timestamp 1621261055
transform 1 0 43200 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_441
timestamp 1621261055
transform 1 0 43488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_438
timestamp 1621261055
transform 1 0 43200 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_906
timestamp 1621261055
transform 1 0 43392 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_454
timestamp 1621261055
transform 1 0 44736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_449
timestamp 1621261055
transform 1 0 44256 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_462
timestamp 1621261055
transform 1 0 45504 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_457
timestamp 1621261055
transform 1 0 45024 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_469
timestamp 1621261055
transform 1 0 46176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_466
timestamp 1621261055
transform 1 0 45888 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_465
timestamp 1621261055
transform 1 0 45792 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_917
timestamp 1621261055
transform 1 0 46080 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_477
timestamp 1621261055
transform 1 0 46944 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_473
timestamp 1621261055
transform 1 0 46560 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_485
timestamp 1621261055
transform 1 0 47712 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_481
timestamp 1621261055
transform 1 0 47328 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_493
timestamp 1621261055
transform 1 0 48480 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_493
timestamp 1621261055
transform 1 0 48480 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_489
timestamp 1621261055
transform 1 0 48096 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_907
timestamp 1621261055
transform 1 0 48672 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_501
timestamp 1621261055
transform 1 0 49248 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_496
timestamp 1621261055
transform 1 0 48768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_509
timestamp 1621261055
transform 1 0 50016 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_512
timestamp 1621261055
transform 1 0 50304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_504
timestamp 1621261055
transform 1 0 49536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_521
timestamp 1621261055
transform 1 0 51168 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_517
timestamp 1621261055
transform 1 0 50784 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_520
timestamp 1621261055
transform 1 0 51072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_524
timestamp 1621261055
transform 1 0 51456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_528
timestamp 1621261055
transform 1 0 51840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_918
timestamp 1621261055
transform 1 0 51360 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_532
timestamp 1621261055
transform 1 0 52224 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_536
timestamp 1621261055
transform 1 0 52608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_540
timestamp 1621261055
transform 1 0 52992 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_544
timestamp 1621261055
transform 1 0 53376 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_548
timestamp 1621261055
transform 1 0 53760 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_551
timestamp 1621261055
transform 1 0 54048 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_548
timestamp 1621261055
transform 1 0 53760 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_87
timestamp 1621261055
transform 1 0 54240 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_908
timestamp 1621261055
transform 1 0 53952 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_556
timestamp 1621261055
transform 1 0 54528 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_558
timestamp 1621261055
transform 1 0 54720 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _170_
timestamp 1621261055
transform 1 0 54432 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_564
timestamp 1621261055
transform 1 0 55296 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_566
timestamp 1621261055
transform 1 0 55488 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _057_
timestamp 1621261055
transform 1 0 55584 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_576
timestamp 1621261055
transform 1 0 56448 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_572
timestamp 1621261055
transform 1 0 56064 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_578
timestamp 1621261055
transform 1 0 56640 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_570
timestamp 1621261055
transform 1 0 55872 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_919
timestamp 1621261055
transform 1 0 56640 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_587
timestamp 1621261055
transform 1 0 57504 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_579
timestamp 1621261055
transform 1 0 56736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_586
timestamp 1621261055
transform 1 0 57408 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_594
timestamp 1621261055
transform 1 0 58176 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_139
timestamp 1621261055
transform -1 0 58848 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_141
timestamp 1621261055
transform -1 0 58848 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_69_596
timestamp 1621261055
transform 1 0 58368 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_595
timestamp 1621261055
transform 1 0 58272 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_142
timestamp 1621261055
transform 1 0 1152 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_4
timestamp 1621261055
transform 1 0 1536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_12
timestamp 1621261055
transform 1 0 2304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_20
timestamp 1621261055
transform 1 0 3072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_28
timestamp 1621261055
transform 1 0 3840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _003_
timestamp 1621261055
transform 1 0 6912 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_920
timestamp 1621261055
transform 1 0 6432 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_36
timestamp 1621261055
transform 1 0 4608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_44
timestamp 1621261055
transform 1 0 5376 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_52
timestamp 1621261055
transform 1 0 6144 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_54
timestamp 1621261055
transform 1 0 6336 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_56
timestamp 1621261055
transform 1 0 6528 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_63
timestamp 1621261055
transform 1 0 7200 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_71
timestamp 1621261055
transform 1 0 7968 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_79
timestamp 1621261055
transform 1 0 8736 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_87
timestamp 1621261055
transform 1 0 9504 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_95
timestamp 1621261055
transform 1 0 10272 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_921
timestamp 1621261055
transform 1 0 11712 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_103
timestamp 1621261055
transform 1 0 11040 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_107
timestamp 1621261055
transform 1 0 11424 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_109
timestamp 1621261055
transform 1 0 11616 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_111
timestamp 1621261055
transform 1 0 11808 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_119
timestamp 1621261055
transform 1 0 12576 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_127
timestamp 1621261055
transform 1 0 13344 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_922
timestamp 1621261055
transform 1 0 16992 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_135
timestamp 1621261055
transform 1 0 14112 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_143
timestamp 1621261055
transform 1 0 14880 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_151
timestamp 1621261055
transform 1 0 15648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_159
timestamp 1621261055
transform 1 0 16416 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_163
timestamp 1621261055
transform 1 0 16800 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_166
timestamp 1621261055
transform 1 0 17088 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_174
timestamp 1621261055
transform 1 0 17856 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_182
timestamp 1621261055
transform 1 0 18624 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_190
timestamp 1621261055
transform 1 0 19392 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_198
timestamp 1621261055
transform 1 0 20160 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _017_
timestamp 1621261055
transform 1 0 23328 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_923
timestamp 1621261055
transform 1 0 22272 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_206
timestamp 1621261055
transform 1 0 20928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_214
timestamp 1621261055
transform 1 0 21696 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_218
timestamp 1621261055
transform 1 0 22080 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_221
timestamp 1621261055
transform 1 0 22368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_229
timestamp 1621261055
transform 1 0 23136 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _159_
timestamp 1621261055
transform 1 0 26400 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_75
timestamp 1621261055
transform 1 0 26208 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_234
timestamp 1621261055
transform 1 0 23616 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_242
timestamp 1621261055
transform 1 0 24384 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_250
timestamp 1621261055
transform 1 0 25152 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_258
timestamp 1621261055
transform 1 0 25920 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_260
timestamp 1621261055
transform 1 0 26112 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _013_
timestamp 1621261055
transform 1 0 29280 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_924
timestamp 1621261055
transform 1 0 27552 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_266
timestamp 1621261055
transform 1 0 26688 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_71_274
timestamp 1621261055
transform 1 0 27456 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_276
timestamp 1621261055
transform 1 0 27648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_284
timestamp 1621261055
transform 1 0 28416 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_71_292
timestamp 1621261055
transform 1 0 29184 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_296
timestamp 1621261055
transform 1 0 29568 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _007_
timestamp 1621261055
transform 1 0 29952 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_925
timestamp 1621261055
transform 1 0 32832 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_303
timestamp 1621261055
transform 1 0 30240 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_311
timestamp 1621261055
transform 1 0 31008 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_319
timestamp 1621261055
transform 1 0 31776 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_327
timestamp 1621261055
transform 1 0 32544 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_329
timestamp 1621261055
transform 1 0 32736 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_331
timestamp 1621261055
transform 1 0 32928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_339
timestamp 1621261055
transform 1 0 33696 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_347
timestamp 1621261055
transform 1 0 34464 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_355
timestamp 1621261055
transform 1 0 35232 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_363
timestamp 1621261055
transform 1 0 36000 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_926
timestamp 1621261055
transform 1 0 38112 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_371
timestamp 1621261055
transform 1 0 36768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_379
timestamp 1621261055
transform 1 0 37536 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_383
timestamp 1621261055
transform 1 0 37920 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_386
timestamp 1621261055
transform 1 0 38208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_394
timestamp 1621261055
transform 1 0 38976 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_402
timestamp 1621261055
transform 1 0 39744 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_410
timestamp 1621261055
transform 1 0 40512 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_418
timestamp 1621261055
transform 1 0 41280 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_426
timestamp 1621261055
transform 1 0 42048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_927
timestamp 1621261055
transform 1 0 43392 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_434
timestamp 1621261055
transform 1 0 42816 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_438
timestamp 1621261055
transform 1 0 43200 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_441
timestamp 1621261055
transform 1 0 43488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_449
timestamp 1621261055
transform 1 0 44256 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_457
timestamp 1621261055
transform 1 0 45024 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _201_
timestamp 1621261055
transform -1 0 47808 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_928
timestamp 1621261055
transform 1 0 48672 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_204
timestamp 1621261055
transform -1 0 47520 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_465
timestamp 1621261055
transform 1 0 45792 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_473
timestamp 1621261055
transform 1 0 46560 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_486
timestamp 1621261055
transform 1 0 47808 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_71_494
timestamp 1621261055
transform 1 0 48576 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_496
timestamp 1621261055
transform 1 0 48768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_504
timestamp 1621261055
transform 1 0 49536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_512
timestamp 1621261055
transform 1 0 50304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_520
timestamp 1621261055
transform 1 0 51072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_528
timestamp 1621261055
transform 1 0 51840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _120_
timestamp 1621261055
transform -1 0 54720 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_929
timestamp 1621261055
transform 1 0 53952 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_152
timestamp 1621261055
transform -1 0 54432 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_536
timestamp 1621261055
transform 1 0 52608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_544
timestamp 1621261055
transform 1 0 53376 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_548
timestamp 1621261055
transform 1 0 53760 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_551
timestamp 1621261055
transform 1 0 54048 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_558
timestamp 1621261055
transform 1 0 54720 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_566
timestamp 1621261055
transform 1 0 55488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_574
timestamp 1621261055
transform 1 0 56256 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_582
timestamp 1621261055
transform 1 0 57024 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_590
timestamp 1621261055
transform 1 0 57792 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_594
timestamp 1621261055
transform 1 0 58176 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_143
timestamp 1621261055
transform -1 0 58848 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_71_596
timestamp 1621261055
transform 1 0 58368 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_144
timestamp 1621261055
transform 1 0 1152 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_930
timestamp 1621261055
transform 1 0 3840 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_4
timestamp 1621261055
transform 1 0 1536 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_12
timestamp 1621261055
transform 1 0 2304 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_20
timestamp 1621261055
transform 1 0 3072 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_29
timestamp 1621261055
transform 1 0 3936 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_37
timestamp 1621261055
transform 1 0 4704 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_45
timestamp 1621261055
transform 1 0 5472 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_53
timestamp 1621261055
transform 1 0 6240 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_61
timestamp 1621261055
transform 1 0 7008 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_931
timestamp 1621261055
transform 1 0 9120 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_154
timestamp 1621261055
transform 1 0 10560 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_69
timestamp 1621261055
transform 1 0 7776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_77
timestamp 1621261055
transform 1 0 8544 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_81
timestamp 1621261055
transform 1 0 8928 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_84
timestamp 1621261055
transform 1 0 9216 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_92
timestamp 1621261055
transform 1 0 9984 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_96
timestamp 1621261055
transform 1 0 10368 0 -1 51282
box -38 -49 230 715
use NOR2X1  NOR2X1
timestamp 1623610208
transform 1 0 10752 0 -1 51282
box 0 -48 864 714
use sky130_fd_sc_ls__decap_8  FILLER_72_109
timestamp 1621261055
transform 1 0 11616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_117
timestamp 1621261055
transform 1 0 12384 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_125
timestamp 1621261055
transform 1 0 13152 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_932
timestamp 1621261055
transform 1 0 14400 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_133
timestamp 1621261055
transform 1 0 13920 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_72_137
timestamp 1621261055
transform 1 0 14304 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_139
timestamp 1621261055
transform 1 0 14496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_147
timestamp 1621261055
transform 1 0 15264 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_155
timestamp 1621261055
transform 1 0 16032 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_163
timestamp 1621261055
transform 1 0 16800 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_933
timestamp 1621261055
transform 1 0 19680 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_171
timestamp 1621261055
transform 1 0 17568 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_179
timestamp 1621261055
transform 1 0 18336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_187
timestamp 1621261055
transform 1 0 19104 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_191
timestamp 1621261055
transform 1 0 19488 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_194
timestamp 1621261055
transform 1 0 19776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _001_
timestamp 1621261055
transform 1 0 20736 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_202
timestamp 1621261055
transform 1 0 20544 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_207
timestamp 1621261055
transform 1 0 21024 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_215
timestamp 1621261055
transform 1 0 21792 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_223
timestamp 1621261055
transform 1 0 22560 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_231
timestamp 1621261055
transform 1 0 23328 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_934
timestamp 1621261055
transform 1 0 24960 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_239
timestamp 1621261055
transform 1 0 24096 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_72_247
timestamp 1621261055
transform 1 0 24864 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_249
timestamp 1621261055
transform 1 0 25056 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_257
timestamp 1621261055
transform 1 0 25824 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _177_
timestamp 1621261055
transform 1 0 27264 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_95
timestamp 1621261055
transform 1 0 27072 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_72_265
timestamp 1621261055
transform 1 0 26592 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_72_269
timestamp 1621261055
transform 1 0 26976 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_275
timestamp 1621261055
transform 1 0 27552 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_283
timestamp 1621261055
transform 1 0 28320 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_291
timestamp 1621261055
transform 1 0 29088 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_935
timestamp 1621261055
transform 1 0 30240 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_299
timestamp 1621261055
transform 1 0 29856 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_72_304
timestamp 1621261055
transform 1 0 30336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_312
timestamp 1621261055
transform 1 0 31104 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_320
timestamp 1621261055
transform 1 0 31872 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_328
timestamp 1621261055
transform 1 0 32640 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_936
timestamp 1621261055
transform 1 0 35520 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_336
timestamp 1621261055
transform 1 0 33408 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_344
timestamp 1621261055
transform 1 0 34176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_352
timestamp 1621261055
transform 1 0 34944 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_356
timestamp 1621261055
transform 1 0 35328 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_359
timestamp 1621261055
transform 1 0 35616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_367
timestamp 1621261055
transform 1 0 36384 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_375
timestamp 1621261055
transform 1 0 37152 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_383
timestamp 1621261055
transform 1 0 37920 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_391
timestamp 1621261055
transform 1 0 38688 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_937
timestamp 1621261055
transform 1 0 40800 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_399
timestamp 1621261055
transform 1 0 39456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_407
timestamp 1621261055
transform 1 0 40224 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_411
timestamp 1621261055
transform 1 0 40608 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_414
timestamp 1621261055
transform 1 0 40896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_422
timestamp 1621261055
transform 1 0 41664 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_430
timestamp 1621261055
transform 1 0 42432 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_438
timestamp 1621261055
transform 1 0 43200 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_446
timestamp 1621261055
transform 1 0 43968 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_454
timestamp 1621261055
transform 1 0 44736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_462
timestamp 1621261055
transform 1 0 45504 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_938
timestamp 1621261055
transform 1 0 46080 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_466
timestamp 1621261055
transform 1 0 45888 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_469
timestamp 1621261055
transform 1 0 46176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_477
timestamp 1621261055
transform 1 0 46944 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_485
timestamp 1621261055
transform 1 0 47712 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_493
timestamp 1621261055
transform 1 0 48480 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_939
timestamp 1621261055
transform 1 0 51360 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_501
timestamp 1621261055
transform 1 0 49248 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_509
timestamp 1621261055
transform 1 0 50016 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_517
timestamp 1621261055
transform 1 0 50784 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_521
timestamp 1621261055
transform 1 0 51168 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_524
timestamp 1621261055
transform 1 0 51456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_532
timestamp 1621261055
transform 1 0 52224 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_540
timestamp 1621261055
transform 1 0 52992 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_548
timestamp 1621261055
transform 1 0 53760 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_556
timestamp 1621261055
transform 1 0 54528 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_940
timestamp 1621261055
transform 1 0 56640 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_564
timestamp 1621261055
transform 1 0 55296 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_572
timestamp 1621261055
transform 1 0 56064 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_576
timestamp 1621261055
transform 1 0 56448 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_579
timestamp 1621261055
transform 1 0 56736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_587
timestamp 1621261055
transform 1 0 57504 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_145
timestamp 1621261055
transform -1 0 58848 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_595
timestamp 1621261055
transform 1 0 58272 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _056_
timestamp 1621261055
transform 1 0 4320 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_146
timestamp 1621261055
transform 1 0 1152 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_73_4
timestamp 1621261055
transform 1 0 1536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_12
timestamp 1621261055
transform 1 0 2304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_20
timestamp 1621261055
transform 1 0 3072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_28
timestamp 1621261055
transform 1 0 3840 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_73_32
timestamp 1621261055
transform 1 0 4224 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_941
timestamp 1621261055
transform 1 0 6432 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_36
timestamp 1621261055
transform 1 0 4608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_44
timestamp 1621261055
transform 1 0 5376 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_52
timestamp 1621261055
transform 1 0 6144 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_54
timestamp 1621261055
transform 1 0 6336 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_56
timestamp 1621261055
transform 1 0 6528 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_64
timestamp 1621261055
transform 1 0 7296 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_72
timestamp 1621261055
transform 1 0 8064 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_80
timestamp 1621261055
transform 1 0 8832 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_88
timestamp 1621261055
transform 1 0 9600 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_96
timestamp 1621261055
transform 1 0 10368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _026_
timestamp 1621261055
transform 1 0 13248 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_942
timestamp 1621261055
transform 1 0 11712 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_104
timestamp 1621261055
transform 1 0 11136 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_108
timestamp 1621261055
transform 1 0 11520 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_111
timestamp 1621261055
transform 1 0 11808 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_119
timestamp 1621261055
transform 1 0 12576 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_123
timestamp 1621261055
transform 1 0 12960 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_125
timestamp 1621261055
transform 1 0 13152 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_129
timestamp 1621261055
transform 1 0 13536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _161_
timestamp 1621261055
transform 1 0 15936 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_943
timestamp 1621261055
transform 1 0 16992 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_77
timestamp 1621261055
transform 1 0 15744 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_137
timestamp 1621261055
transform 1 0 14304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_145
timestamp 1621261055
transform 1 0 15072 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_149
timestamp 1621261055
transform 1 0 15456 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_151
timestamp 1621261055
transform 1 0 15648 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_157
timestamp 1621261055
transform 1 0 16224 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_166
timestamp 1621261055
transform 1 0 17088 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_174
timestamp 1621261055
transform 1 0 17856 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_182
timestamp 1621261055
transform 1 0 18624 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_190
timestamp 1621261055
transform 1 0 19392 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_198
timestamp 1621261055
transform 1 0 20160 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_944
timestamp 1621261055
transform 1 0 22272 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_107
timestamp 1621261055
transform -1 0 23424 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_206
timestamp 1621261055
transform 1 0 20928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_214
timestamp 1621261055
transform 1 0 21696 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_218
timestamp 1621261055
transform 1 0 22080 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_221
timestamp 1621261055
transform 1 0 22368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_73_229
timestamp 1621261055
transform 1 0 23136 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _072_
timestamp 1621261055
transform -1 0 23712 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_73_235
timestamp 1621261055
transform 1 0 23712 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_243
timestamp 1621261055
transform 1 0 24480 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_251
timestamp 1621261055
transform 1 0 25248 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_259
timestamp 1621261055
transform 1 0 26016 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_945
timestamp 1621261055
transform 1 0 27552 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_267
timestamp 1621261055
transform 1 0 26784 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_276
timestamp 1621261055
transform 1 0 27648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_284
timestamp 1621261055
transform 1 0 28416 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_292
timestamp 1621261055
transform 1 0 29184 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_946
timestamp 1621261055
transform 1 0 32832 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_300
timestamp 1621261055
transform 1 0 29952 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_308
timestamp 1621261055
transform 1 0 30720 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_316
timestamp 1621261055
transform 1 0 31488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_324
timestamp 1621261055
transform 1 0 32256 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_328
timestamp 1621261055
transform 1 0 32640 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_331
timestamp 1621261055
transform 1 0 32928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_339
timestamp 1621261055
transform 1 0 33696 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_347
timestamp 1621261055
transform 1 0 34464 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_355
timestamp 1621261055
transform 1 0 35232 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_363
timestamp 1621261055
transform 1 0 36000 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_947
timestamp 1621261055
transform 1 0 38112 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_371
timestamp 1621261055
transform 1 0 36768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_379
timestamp 1621261055
transform 1 0 37536 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_383
timestamp 1621261055
transform 1 0 37920 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_386
timestamp 1621261055
transform 1 0 38208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_394
timestamp 1621261055
transform 1 0 38976 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_402
timestamp 1621261055
transform 1 0 39744 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_410
timestamp 1621261055
transform 1 0 40512 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_418
timestamp 1621261055
transform 1 0 41280 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_426
timestamp 1621261055
transform 1 0 42048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_948
timestamp 1621261055
transform 1 0 43392 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_434
timestamp 1621261055
transform 1 0 42816 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_438
timestamp 1621261055
transform 1 0 43200 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_441
timestamp 1621261055
transform 1 0 43488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_449
timestamp 1621261055
transform 1 0 44256 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_457
timestamp 1621261055
transform 1 0 45024 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_949
timestamp 1621261055
transform 1 0 48672 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_465
timestamp 1621261055
transform 1 0 45792 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_473
timestamp 1621261055
transform 1 0 46560 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_481
timestamp 1621261055
transform 1 0 47328 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_489
timestamp 1621261055
transform 1 0 48096 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_493
timestamp 1621261055
transform 1 0 48480 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_496
timestamp 1621261055
transform 1 0 48768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_504
timestamp 1621261055
transform 1 0 49536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_512
timestamp 1621261055
transform 1 0 50304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_520
timestamp 1621261055
transform 1 0 51072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_528
timestamp 1621261055
transform 1 0 51840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_950
timestamp 1621261055
transform 1 0 53952 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_536
timestamp 1621261055
transform 1 0 52608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_544
timestamp 1621261055
transform 1 0 53376 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_548
timestamp 1621261055
transform 1 0 53760 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_551
timestamp 1621261055
transform 1 0 54048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_559
timestamp 1621261055
transform 1 0 54816 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_567
timestamp 1621261055
transform 1 0 55584 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_575
timestamp 1621261055
transform 1 0 56352 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_583
timestamp 1621261055
transform 1 0 57120 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_591
timestamp 1621261055
transform 1 0 57888 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_147
timestamp 1621261055
transform -1 0 58848 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_595
timestamp 1621261055
transform 1 0 58272 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_148
timestamp 1621261055
transform 1 0 1152 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_951
timestamp 1621261055
transform 1 0 3840 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_4
timestamp 1621261055
transform 1 0 1536 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_12
timestamp 1621261055
transform 1 0 2304 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_20
timestamp 1621261055
transform 1 0 3072 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_29
timestamp 1621261055
transform 1 0 3936 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_37
timestamp 1621261055
transform 1 0 4704 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_45
timestamp 1621261055
transform 1 0 5472 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_53
timestamp 1621261055
transform 1 0 6240 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_61
timestamp 1621261055
transform 1 0 7008 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_952
timestamp 1621261055
transform 1 0 9120 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_69
timestamp 1621261055
transform 1 0 7776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_77
timestamp 1621261055
transform 1 0 8544 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_81
timestamp 1621261055
transform 1 0 8928 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_84
timestamp 1621261055
transform 1 0 9216 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_92
timestamp 1621261055
transform 1 0 9984 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_100
timestamp 1621261055
transform 1 0 10752 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_108
timestamp 1621261055
transform 1 0 11520 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_116
timestamp 1621261055
transform 1 0 12288 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_124
timestamp 1621261055
transform 1 0 13056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_132
timestamp 1621261055
transform 1 0 13824 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_953
timestamp 1621261055
transform 1 0 14400 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_136
timestamp 1621261055
transform 1 0 14208 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_139
timestamp 1621261055
transform 1 0 14496 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_147
timestamp 1621261055
transform 1 0 15264 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_155
timestamp 1621261055
transform 1 0 16032 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_163
timestamp 1621261055
transform 1 0 16800 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _077_
timestamp 1621261055
transform 1 0 17760 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _183_
timestamp 1621261055
transform -1 0 20448 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_954
timestamp 1621261055
transform 1 0 19680 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_117
timestamp 1621261055
transform 1 0 17568 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_206
timestamp 1621261055
transform -1 0 20160 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_176
timestamp 1621261055
transform 1 0 18048 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_184
timestamp 1621261055
transform 1 0 18816 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_74_192
timestamp 1621261055
transform 1 0 19584 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_194
timestamp 1621261055
transform 1 0 19776 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_201
timestamp 1621261055
transform 1 0 20448 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_209
timestamp 1621261055
transform 1 0 21216 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_217
timestamp 1621261055
transform 1 0 21984 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_225
timestamp 1621261055
transform 1 0 22752 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_955
timestamp 1621261055
transform 1 0 24960 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_233
timestamp 1621261055
transform 1 0 23520 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_241
timestamp 1621261055
transform 1 0 24288 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_245
timestamp 1621261055
transform 1 0 24672 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_74_247
timestamp 1621261055
transform 1 0 24864 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_249
timestamp 1621261055
transform 1 0 25056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_257
timestamp 1621261055
transform 1 0 25824 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_265
timestamp 1621261055
transform 1 0 26592 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_273
timestamp 1621261055
transform 1 0 27360 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_281
timestamp 1621261055
transform 1 0 28128 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_289
timestamp 1621261055
transform 1 0 28896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_297
timestamp 1621261055
transform 1 0 29664 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _167_
timestamp 1621261055
transform 1 0 32448 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_956
timestamp 1621261055
transform 1 0 30240 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_82
timestamp 1621261055
transform 1 0 32256 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_301
timestamp 1621261055
transform 1 0 30048 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_304
timestamp 1621261055
transform 1 0 30336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_312
timestamp 1621261055
transform 1 0 31104 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_320
timestamp 1621261055
transform 1 0 31872 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_329
timestamp 1621261055
transform 1 0 32736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_957
timestamp 1621261055
transform 1 0 35520 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_337
timestamp 1621261055
transform 1 0 33504 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_345
timestamp 1621261055
transform 1 0 34272 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_353
timestamp 1621261055
transform 1 0 35040 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_74_357
timestamp 1621261055
transform 1 0 35424 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_359
timestamp 1621261055
transform 1 0 35616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_367
timestamp 1621261055
transform 1 0 36384 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_375
timestamp 1621261055
transform 1 0 37152 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_383
timestamp 1621261055
transform 1 0 37920 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_391
timestamp 1621261055
transform 1 0 38688 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_958
timestamp 1621261055
transform 1 0 40800 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_399
timestamp 1621261055
transform 1 0 39456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_407
timestamp 1621261055
transform 1 0 40224 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_411
timestamp 1621261055
transform 1 0 40608 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_414
timestamp 1621261055
transform 1 0 40896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_422
timestamp 1621261055
transform 1 0 41664 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_430
timestamp 1621261055
transform 1 0 42432 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_438
timestamp 1621261055
transform 1 0 43200 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_446
timestamp 1621261055
transform 1 0 43968 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_454
timestamp 1621261055
transform 1 0 44736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_462
timestamp 1621261055
transform 1 0 45504 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_959
timestamp 1621261055
transform 1 0 46080 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_466
timestamp 1621261055
transform 1 0 45888 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_469
timestamp 1621261055
transform 1 0 46176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_477
timestamp 1621261055
transform 1 0 46944 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_485
timestamp 1621261055
transform 1 0 47712 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_493
timestamp 1621261055
transform 1 0 48480 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_960
timestamp 1621261055
transform 1 0 51360 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_501
timestamp 1621261055
transform 1 0 49248 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_509
timestamp 1621261055
transform 1 0 50016 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_517
timestamp 1621261055
transform 1 0 50784 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_521
timestamp 1621261055
transform 1 0 51168 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_524
timestamp 1621261055
transform 1 0 51456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_532
timestamp 1621261055
transform 1 0 52224 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_540
timestamp 1621261055
transform 1 0 52992 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_548
timestamp 1621261055
transform 1 0 53760 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_556
timestamp 1621261055
transform 1 0 54528 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_961
timestamp 1621261055
transform 1 0 56640 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_564
timestamp 1621261055
transform 1 0 55296 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_572
timestamp 1621261055
transform 1 0 56064 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_576
timestamp 1621261055
transform 1 0 56448 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_579
timestamp 1621261055
transform 1 0 56736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_587
timestamp 1621261055
transform 1 0 57504 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_149
timestamp 1621261055
transform -1 0 58848 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_595
timestamp 1621261055
transform 1 0 58272 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_150
timestamp 1621261055
transform 1 0 1152 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_75_4
timestamp 1621261055
transform 1 0 1536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_12
timestamp 1621261055
transform 1 0 2304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_20
timestamp 1621261055
transform 1 0 3072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_28
timestamp 1621261055
transform 1 0 3840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_962
timestamp 1621261055
transform 1 0 6432 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_36
timestamp 1621261055
transform 1 0 4608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_44
timestamp 1621261055
transform 1 0 5376 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_52
timestamp 1621261055
transform 1 0 6144 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_54
timestamp 1621261055
transform 1 0 6336 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_56
timestamp 1621261055
transform 1 0 6528 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_64
timestamp 1621261055
transform 1 0 7296 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_72
timestamp 1621261055
transform 1 0 8064 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_80
timestamp 1621261055
transform 1 0 8832 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_88
timestamp 1621261055
transform 1 0 9600 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_96
timestamp 1621261055
transform 1 0 10368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_963
timestamp 1621261055
transform 1 0 11712 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_104
timestamp 1621261055
transform 1 0 11136 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_108
timestamp 1621261055
transform 1 0 11520 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_111
timestamp 1621261055
transform 1 0 11808 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_119
timestamp 1621261055
transform 1 0 12576 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_127
timestamp 1621261055
transform 1 0 13344 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_964
timestamp 1621261055
transform 1 0 16992 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_135
timestamp 1621261055
transform 1 0 14112 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_143
timestamp 1621261055
transform 1 0 14880 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_151
timestamp 1621261055
transform 1 0 15648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_159
timestamp 1621261055
transform 1 0 16416 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_163
timestamp 1621261055
transform 1 0 16800 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_166
timestamp 1621261055
transform 1 0 17088 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_174
timestamp 1621261055
transform 1 0 17856 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_182
timestamp 1621261055
transform 1 0 18624 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_190
timestamp 1621261055
transform 1 0 19392 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_198
timestamp 1621261055
transform 1 0 20160 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_965
timestamp 1621261055
transform 1 0 22272 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_206
timestamp 1621261055
transform 1 0 20928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_214
timestamp 1621261055
transform 1 0 21696 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_218
timestamp 1621261055
transform 1 0 22080 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_221
timestamp 1621261055
transform 1 0 22368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_229
timestamp 1621261055
transform 1 0 23136 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_237
timestamp 1621261055
transform 1 0 23904 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_245
timestamp 1621261055
transform 1 0 24672 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_253
timestamp 1621261055
transform 1 0 25440 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_261
timestamp 1621261055
transform 1 0 26208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _064_
timestamp 1621261055
transform -1 0 29952 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_966
timestamp 1621261055
transform 1 0 27552 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_166
timestamp 1621261055
transform -1 0 29664 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_75_269
timestamp 1621261055
transform 1 0 26976 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_273
timestamp 1621261055
transform 1 0 27360 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_276
timestamp 1621261055
transform 1 0 27648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_284
timestamp 1621261055
transform 1 0 28416 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_292
timestamp 1621261055
transform 1 0 29184 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_294
timestamp 1621261055
transform 1 0 29376 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_967
timestamp 1621261055
transform 1 0 32832 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_300
timestamp 1621261055
transform 1 0 29952 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_308
timestamp 1621261055
transform 1 0 30720 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_316
timestamp 1621261055
transform 1 0 31488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_324
timestamp 1621261055
transform 1 0 32256 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_328
timestamp 1621261055
transform 1 0 32640 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_331
timestamp 1621261055
transform 1 0 32928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_339
timestamp 1621261055
transform 1 0 33696 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_347
timestamp 1621261055
transform 1 0 34464 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_355
timestamp 1621261055
transform 1 0 35232 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_363
timestamp 1621261055
transform 1 0 36000 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_968
timestamp 1621261055
transform 1 0 38112 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_371
timestamp 1621261055
transform 1 0 36768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_379
timestamp 1621261055
transform 1 0 37536 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_383
timestamp 1621261055
transform 1 0 37920 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_386
timestamp 1621261055
transform 1 0 38208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_394
timestamp 1621261055
transform 1 0 38976 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_402
timestamp 1621261055
transform 1 0 39744 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_410
timestamp 1621261055
transform 1 0 40512 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_418
timestamp 1621261055
transform 1 0 41280 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_426
timestamp 1621261055
transform 1 0 42048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_969
timestamp 1621261055
transform 1 0 43392 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_434
timestamp 1621261055
transform 1 0 42816 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_438
timestamp 1621261055
transform 1 0 43200 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_441
timestamp 1621261055
transform 1 0 43488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_449
timestamp 1621261055
transform 1 0 44256 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_457
timestamp 1621261055
transform 1 0 45024 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_970
timestamp 1621261055
transform 1 0 48672 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_465
timestamp 1621261055
transform 1 0 45792 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_473
timestamp 1621261055
transform 1 0 46560 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_481
timestamp 1621261055
transform 1 0 47328 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_489
timestamp 1621261055
transform 1 0 48096 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_493
timestamp 1621261055
transform 1 0 48480 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_496
timestamp 1621261055
transform 1 0 48768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_504
timestamp 1621261055
transform 1 0 49536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_512
timestamp 1621261055
transform 1 0 50304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_520
timestamp 1621261055
transform 1 0 51072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_528
timestamp 1621261055
transform 1 0 51840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_971
timestamp 1621261055
transform 1 0 53952 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_536
timestamp 1621261055
transform 1 0 52608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_544
timestamp 1621261055
transform 1 0 53376 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_548
timestamp 1621261055
transform 1 0 53760 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_551
timestamp 1621261055
transform 1 0 54048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_559
timestamp 1621261055
transform 1 0 54816 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _066_
timestamp 1621261055
transform -1 0 56544 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_188
timestamp 1621261055
transform -1 0 56256 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_75_567
timestamp 1621261055
transform 1 0 55584 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_75_571
timestamp 1621261055
transform 1 0 55968 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_577
timestamp 1621261055
transform 1 0 56544 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_585
timestamp 1621261055
transform 1 0 57312 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_593
timestamp 1621261055
transform 1 0 58080 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_151
timestamp 1621261055
transform -1 0 58848 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_152
timestamp 1621261055
transform 1 0 1152 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_972
timestamp 1621261055
transform 1 0 3840 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_4
timestamp 1621261055
transform 1 0 1536 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_12
timestamp 1621261055
transform 1 0 2304 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_20
timestamp 1621261055
transform 1 0 3072 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_29
timestamp 1621261055
transform 1 0 3936 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_37
timestamp 1621261055
transform 1 0 4704 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_45
timestamp 1621261055
transform 1 0 5472 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_53
timestamp 1621261055
transform 1 0 6240 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_61
timestamp 1621261055
transform 1 0 7008 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_973
timestamp 1621261055
transform 1 0 9120 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_69
timestamp 1621261055
transform 1 0 7776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_77
timestamp 1621261055
transform 1 0 8544 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_81
timestamp 1621261055
transform 1 0 8928 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_84
timestamp 1621261055
transform 1 0 9216 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_92
timestamp 1621261055
transform 1 0 9984 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_100
timestamp 1621261055
transform 1 0 10752 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_108
timestamp 1621261055
transform 1 0 11520 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_116
timestamp 1621261055
transform 1 0 12288 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_124
timestamp 1621261055
transform 1 0 13056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_132
timestamp 1621261055
transform 1 0 13824 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_974
timestamp 1621261055
transform 1 0 14400 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_136
timestamp 1621261055
transform 1 0 14208 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_139
timestamp 1621261055
transform 1 0 14496 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_147
timestamp 1621261055
transform 1 0 15264 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_155
timestamp 1621261055
transform 1 0 16032 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_163
timestamp 1621261055
transform 1 0 16800 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_975
timestamp 1621261055
transform 1 0 19680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_171
timestamp 1621261055
transform 1 0 17568 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_179
timestamp 1621261055
transform 1 0 18336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_187
timestamp 1621261055
transform 1 0 19104 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_191
timestamp 1621261055
transform 1 0 19488 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_194
timestamp 1621261055
transform 1 0 19776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _089_
timestamp 1621261055
transform 1 0 22368 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_123
timestamp 1621261055
transform 1 0 22176 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_202
timestamp 1621261055
transform 1 0 20544 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_210
timestamp 1621261055
transform 1 0 21312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_76_218
timestamp 1621261055
transform 1 0 22080 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_224
timestamp 1621261055
transform 1 0 22656 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_976
timestamp 1621261055
transform 1 0 24960 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_232
timestamp 1621261055
transform 1 0 23424 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_240
timestamp 1621261055
transform 1 0 24192 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_249
timestamp 1621261055
transform 1 0 25056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_257
timestamp 1621261055
transform 1 0 25824 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_265
timestamp 1621261055
transform 1 0 26592 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_273
timestamp 1621261055
transform 1 0 27360 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_281
timestamp 1621261055
transform 1 0 28128 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_289
timestamp 1621261055
transform 1 0 28896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_297
timestamp 1621261055
transform 1 0 29664 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_977
timestamp 1621261055
transform 1 0 30240 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_301
timestamp 1621261055
transform 1 0 30048 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_304
timestamp 1621261055
transform 1 0 30336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_312
timestamp 1621261055
transform 1 0 31104 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_320
timestamp 1621261055
transform 1 0 31872 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_328
timestamp 1621261055
transform 1 0 32640 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_978
timestamp 1621261055
transform 1 0 35520 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_336
timestamp 1621261055
transform 1 0 33408 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_344
timestamp 1621261055
transform 1 0 34176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_352
timestamp 1621261055
transform 1 0 34944 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_356
timestamp 1621261055
transform 1 0 35328 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_359
timestamp 1621261055
transform 1 0 35616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_367
timestamp 1621261055
transform 1 0 36384 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_375
timestamp 1621261055
transform 1 0 37152 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_383
timestamp 1621261055
transform 1 0 37920 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_391
timestamp 1621261055
transform 1 0 38688 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_979
timestamp 1621261055
transform 1 0 40800 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_399
timestamp 1621261055
transform 1 0 39456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_407
timestamp 1621261055
transform 1 0 40224 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_411
timestamp 1621261055
transform 1 0 40608 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_414
timestamp 1621261055
transform 1 0 40896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_422
timestamp 1621261055
transform 1 0 41664 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _153_
timestamp 1621261055
transform 1 0 45024 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_73
timestamp 1621261055
transform 1 0 44832 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_430
timestamp 1621261055
transform 1 0 42432 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_438
timestamp 1621261055
transform 1 0 43200 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_446
timestamp 1621261055
transform 1 0 43968 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_76_454
timestamp 1621261055
transform 1 0 44736 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_460
timestamp 1621261055
transform 1 0 45312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_980
timestamp 1621261055
transform 1 0 46080 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_469
timestamp 1621261055
transform 1 0 46176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_477
timestamp 1621261055
transform 1 0 46944 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_485
timestamp 1621261055
transform 1 0 47712 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_493
timestamp 1621261055
transform 1 0 48480 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_981
timestamp 1621261055
transform 1 0 51360 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_501
timestamp 1621261055
transform 1 0 49248 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_509
timestamp 1621261055
transform 1 0 50016 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_517
timestamp 1621261055
transform 1 0 50784 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_521
timestamp 1621261055
transform 1 0 51168 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_524
timestamp 1621261055
transform 1 0 51456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_532
timestamp 1621261055
transform 1 0 52224 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_540
timestamp 1621261055
transform 1 0 52992 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_548
timestamp 1621261055
transform 1 0 53760 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_556
timestamp 1621261055
transform 1 0 54528 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_982
timestamp 1621261055
transform 1 0 56640 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output436
timestamp 1621261055
transform -1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_66
timestamp 1621261055
transform -1 0 57696 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_564
timestamp 1621261055
transform 1 0 55296 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_572
timestamp 1621261055
transform 1 0 56064 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_576
timestamp 1621261055
transform 1 0 56448 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_579
timestamp 1621261055
transform 1 0 56736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_593
timestamp 1621261055
transform 1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_153
timestamp 1621261055
transform -1 0 58848 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_4
timestamp 1621261055
transform 1 0 1536 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_4
timestamp 1621261055
transform 1 0 1536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_156
timestamp 1621261055
transform 1 0 1152 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_154
timestamp 1621261055
transform 1 0 1152 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_12
timestamp 1621261055
transform 1 0 2304 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_12
timestamp 1621261055
transform 1 0 2304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_20
timestamp 1621261055
transform 1 0 3072 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_20
timestamp 1621261055
transform 1 0 3072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_29
timestamp 1621261055
transform 1 0 3936 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_28
timestamp 1621261055
transform 1 0 3840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_993
timestamp 1621261055
transform 1 0 3840 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_37
timestamp 1621261055
transform 1 0 4704 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_36
timestamp 1621261055
transform 1 0 4608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_45
timestamp 1621261055
transform 1 0 5472 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_44
timestamp 1621261055
transform 1 0 5376 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_53
timestamp 1621261055
transform 1 0 6240 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_56
timestamp 1621261055
transform 1 0 6528 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_54
timestamp 1621261055
transform 1 0 6336 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_52
timestamp 1621261055
transform 1 0 6144 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_983
timestamp 1621261055
transform 1 0 6432 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_61
timestamp 1621261055
transform 1 0 7008 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_64
timestamp 1621261055
transform 1 0 7296 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_69
timestamp 1621261055
transform 1 0 7776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_72
timestamp 1621261055
transform 1 0 8064 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_81
timestamp 1621261055
transform 1 0 8928 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_77
timestamp 1621261055
transform 1 0 8544 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_80
timestamp 1621261055
transform 1 0 8832 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_994
timestamp 1621261055
transform 1 0 9120 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_92
timestamp 1621261055
transform 1 0 9984 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_84
timestamp 1621261055
transform 1 0 9216 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_88
timestamp 1621261055
transform 1 0 9600 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_96
timestamp 1621261055
transform 1 0 10368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_100
timestamp 1621261055
transform 1 0 10752 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_104
timestamp 1621261055
transform 1 0 11136 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_116
timestamp 1621261055
transform 1 0 12288 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_108
timestamp 1621261055
transform 1 0 11520 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_111
timestamp 1621261055
transform 1 0 11808 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_108
timestamp 1621261055
transform 1 0 11520 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_984
timestamp 1621261055
transform 1 0 11712 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_124
timestamp 1621261055
transform 1 0 13056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_119
timestamp 1621261055
transform 1 0 12576 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_132
timestamp 1621261055
transform 1 0 13824 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_127
timestamp 1621261055
transform 1 0 13344 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_139
timestamp 1621261055
transform 1 0 14496 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_136
timestamp 1621261055
transform 1 0 14208 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_135
timestamp 1621261055
transform 1 0 14112 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_995
timestamp 1621261055
transform 1 0 14400 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_147
timestamp 1621261055
transform 1 0 15264 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_143
timestamp 1621261055
transform 1 0 14880 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_155
timestamp 1621261055
transform 1 0 16032 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_151
timestamp 1621261055
transform 1 0 15648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_163
timestamp 1621261055
transform 1 0 16800 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_163
timestamp 1621261055
transform 1 0 16800 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_159
timestamp 1621261055
transform 1 0 16416 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_985
timestamp 1621261055
transform 1 0 16992 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_171
timestamp 1621261055
transform 1 0 17568 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_166
timestamp 1621261055
transform 1 0 17088 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_179
timestamp 1621261055
transform 1 0 18336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_182
timestamp 1621261055
transform 1 0 18624 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_174
timestamp 1621261055
transform 1 0 17856 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_191
timestamp 1621261055
transform 1 0 19488 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_187
timestamp 1621261055
transform 1 0 19104 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_190
timestamp 1621261055
transform 1 0 19392 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_194
timestamp 1621261055
transform 1 0 19776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_198
timestamp 1621261055
transform 1 0 20160 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_996
timestamp 1621261055
transform 1 0 19680 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_202
timestamp 1621261055
transform 1 0 20544 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_206
timestamp 1621261055
transform 1 0 20928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_210
timestamp 1621261055
transform 1 0 21312 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_214
timestamp 1621261055
transform 1 0 21696 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_218
timestamp 1621261055
transform 1 0 22080 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_221
timestamp 1621261055
transform 1 0 22368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_218
timestamp 1621261055
transform 1 0 22080 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_986
timestamp 1621261055
transform 1 0 22272 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_226
timestamp 1621261055
transform 1 0 22848 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_229
timestamp 1621261055
transform 1 0 23136 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_234
timestamp 1621261055
transform 1 0 23616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_237
timestamp 1621261055
transform 1 0 23904 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_246
timestamp 1621261055
transform 1 0 24768 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_242
timestamp 1621261055
transform 1 0 24384 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_245
timestamp 1621261055
transform 1 0 24672 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_997
timestamp 1621261055
transform 1 0 24960 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_257
timestamp 1621261055
transform 1 0 25824 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_249
timestamp 1621261055
transform 1 0 25056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_253
timestamp 1621261055
transform 1 0 25440 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_261
timestamp 1621261055
transform 1 0 26208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_265
timestamp 1621261055
transform 1 0 26592 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_269
timestamp 1621261055
transform 1 0 26976 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_281
timestamp 1621261055
transform 1 0 28128 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_273
timestamp 1621261055
transform 1 0 27360 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_276
timestamp 1621261055
transform 1 0 27648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_273
timestamp 1621261055
transform 1 0 27360 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_987
timestamp 1621261055
transform 1 0 27552 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_289
timestamp 1621261055
transform 1 0 28896 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_284
timestamp 1621261055
transform 1 0 28416 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_297
timestamp 1621261055
transform 1 0 29664 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_292
timestamp 1621261055
transform 1 0 29184 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_304
timestamp 1621261055
transform 1 0 30336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_301
timestamp 1621261055
transform 1 0 30048 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_300
timestamp 1621261055
transform 1 0 29952 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_998
timestamp 1621261055
transform 1 0 30240 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_312
timestamp 1621261055
transform 1 0 31104 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_308
timestamp 1621261055
transform 1 0 30720 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_320
timestamp 1621261055
transform 1 0 31872 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_316
timestamp 1621261055
transform 1 0 31488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_328
timestamp 1621261055
transform 1 0 32640 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_328
timestamp 1621261055
transform 1 0 32640 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_324
timestamp 1621261055
transform 1 0 32256 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_988
timestamp 1621261055
transform 1 0 32832 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_344
timestamp 1621261055
transform 1 0 34176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_336
timestamp 1621261055
transform 1 0 33408 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_339
timestamp 1621261055
transform 1 0 33696 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_331
timestamp 1621261055
transform 1 0 32928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_113
timestamp 1621261055
transform 1 0 33888 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_359
timestamp 1621261055
transform 1 0 35616 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_356
timestamp 1621261055
transform 1 0 35328 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_352
timestamp 1621261055
transform 1 0 34944 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_125
timestamp 1621261055
transform -1 0 36000 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_999
timestamp 1621261055
transform 1 0 35520 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _092_
timestamp 1621261055
transform -1 0 36288 0 -1 55278
box -38 -49 326 715
use XNOR2X1  XNOR2X1
timestamp 1623610208
transform 1 0 34080 0 1 53946
box 0 -48 2016 714
use sky130_fd_sc_ls__decap_8  FILLER_78_366
timestamp 1621261055
transform 1 0 36288 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_371
timestamp 1621261055
transform 1 0 36768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_364
timestamp 1621261055
transform 1 0 36096 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_220
timestamp 1621261055
transform -1 0 36480 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _213_
timestamp 1621261055
transform -1 0 36768 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_374
timestamp 1621261055
transform 1 0 37056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_379
timestamp 1621261055
transform 1 0 37536 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_382
timestamp 1621261055
transform 1 0 37824 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_386
timestamp 1621261055
transform 1 0 38208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_383
timestamp 1621261055
transform 1 0 37920 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_989
timestamp 1621261055
transform 1 0 38112 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_78_394
timestamp 1621261055
transform 1 0 38976 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_390
timestamp 1621261055
transform 1 0 38592 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_394
timestamp 1621261055
transform 1 0 38976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output422
timestamp 1621261055
transform 1 0 39072 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_399
timestamp 1621261055
transform 1 0 39456 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_402
timestamp 1621261055
transform 1 0 39744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_103
timestamp 1621261055
transform -1 0 39840 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _070_
timestamp 1621261055
transform -1 0 40128 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_78_412
timestamp 1621261055
transform 1 0 40704 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_410
timestamp 1621261055
transform 1 0 40512 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_406
timestamp 1621261055
transform 1 0 40128 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_410
timestamp 1621261055
transform 1 0 40512 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1000
timestamp 1621261055
transform 1 0 40800 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_422
timestamp 1621261055
transform 1 0 41664 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_414
timestamp 1621261055
transform 1 0 40896 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_418
timestamp 1621261055
transform 1 0 41280 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_426
timestamp 1621261055
transform 1 0 42048 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_430
timestamp 1621261055
transform 1 0 42432 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_437
timestamp 1621261055
transform 1 0 43104 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_433
timestamp 1621261055
transform 1 0 42720 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _039_
timestamp 1621261055
transform 1 0 42432 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_446
timestamp 1621261055
transform 1 0 43968 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_438
timestamp 1621261055
transform 1 0 43200 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_441
timestamp 1621261055
transform 1 0 43488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_439
timestamp 1621261055
transform 1 0 43296 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_990
timestamp 1621261055
transform 1 0 43392 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_454
timestamp 1621261055
transform 1 0 44736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_449
timestamp 1621261055
transform 1 0 44256 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_462
timestamp 1621261055
transform 1 0 45504 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_457
timestamp 1621261055
transform 1 0 45024 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_469
timestamp 1621261055
transform 1 0 46176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_466
timestamp 1621261055
transform 1 0 45888 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_465
timestamp 1621261055
transform 1 0 45792 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1001
timestamp 1621261055
transform 1 0 46080 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_477
timestamp 1621261055
transform 1 0 46944 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_473
timestamp 1621261055
transform 1 0 46560 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_485
timestamp 1621261055
transform 1 0 47712 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_481
timestamp 1621261055
transform 1 0 47328 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_493
timestamp 1621261055
transform 1 0 48480 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_493
timestamp 1621261055
transform 1 0 48480 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_489
timestamp 1621261055
transform 1 0 48096 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_991
timestamp 1621261055
transform 1 0 48672 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_501
timestamp 1621261055
transform 1 0 49248 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_496
timestamp 1621261055
transform 1 0 48768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_509
timestamp 1621261055
transform 1 0 50016 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_512
timestamp 1621261055
transform 1 0 50304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_504
timestamp 1621261055
transform 1 0 49536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_521
timestamp 1621261055
transform 1 0 51168 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_517
timestamp 1621261055
transform 1 0 50784 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_520
timestamp 1621261055
transform 1 0 51072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_524
timestamp 1621261055
transform 1 0 51456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_528
timestamp 1621261055
transform 1 0 51840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1002
timestamp 1621261055
transform 1 0 51360 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_532
timestamp 1621261055
transform 1 0 52224 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_536
timestamp 1621261055
transform 1 0 52608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_540
timestamp 1621261055
transform 1 0 52992 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_544
timestamp 1621261055
transform 1 0 53376 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_554
timestamp 1621261055
transform 1 0 54336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_548
timestamp 1621261055
transform 1 0 53760 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_551
timestamp 1621261055
transform 1 0 54048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_548
timestamp 1621261055
transform 1 0 53760 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_190
timestamp 1621261055
transform -1 0 54048 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_992
timestamp 1621261055
transform 1 0 53952 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _181_
timestamp 1621261055
transform -1 0 54336 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_77_559
timestamp 1621261055
transform 1 0 54816 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_566
timestamp 1621261055
transform 1 0 55488 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_562
timestamp 1621261055
transform 1 0 55104 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_567
timestamp 1621261055
transform 1 0 55584 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_101
timestamp 1621261055
transform -1 0 55776 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _069_
timestamp 1621261055
transform -1 0 56064 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_576
timestamp 1621261055
transform 1 0 56448 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_572
timestamp 1621261055
transform 1 0 56064 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_575
timestamp 1621261055
transform 1 0 56352 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1003
timestamp 1621261055
transform 1 0 56640 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_587
timestamp 1621261055
transform 1 0 57504 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_579
timestamp 1621261055
transform 1 0 56736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_587
timestamp 1621261055
transform 1 0 57504 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_583
timestamp 1621261055
transform 1 0 57120 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_78_593
timestamp 1621261055
transform 1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_77_593
timestamp 1621261055
transform 1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output435
timestamp 1621261055
transform 1 0 57696 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output398
timestamp 1621261055
transform 1 0 57696 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_155
timestamp 1621261055
transform -1 0 58848 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_157
timestamp 1621261055
transform -1 0 58848 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_158
timestamp 1621261055
transform 1 0 1152 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output406
timestamp 1621261055
transform 1 0 1536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output428
timestamp 1621261055
transform 1 0 4320 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_33
timestamp 1621261055
transform 1 0 1920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_10
timestamp 1621261055
transform 1 0 2112 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_18
timestamp 1621261055
transform 1 0 2880 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_26
timestamp 1621261055
transform 1 0 3648 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_30
timestamp 1621261055
transform 1 0 4032 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_32
timestamp 1621261055
transform 1 0 4224 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1004
timestamp 1621261055
transform 1 0 6432 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output438
timestamp 1621261055
transform 1 0 7488 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_68
timestamp 1621261055
transform 1 0 7296 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_37
timestamp 1621261055
transform 1 0 4704 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_45
timestamp 1621261055
transform 1 0 5472 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_53
timestamp 1621261055
transform 1 0 6240 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_56
timestamp 1621261055
transform 1 0 6528 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output439
timestamp 1621261055
transform 1 0 9120 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_70
timestamp 1621261055
transform 1 0 7872 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_78
timestamp 1621261055
transform 1 0 8640 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_82
timestamp 1621261055
transform 1 0 9024 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_87
timestamp 1621261055
transform 1 0 9504 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_95
timestamp 1621261055
transform 1 0 10272 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_107
timestamp 1621261055
transform 1 0 11424 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_103
timestamp 1621261055
transform 1 0 11040 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_111
timestamp 1621261055
transform 1 0 11808 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_109
timestamp 1621261055
transform 1 0 11616 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_129
timestamp 1621261055
transform 1 0 12000 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1005
timestamp 1621261055
transform 1 0 11712 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _093_
timestamp 1621261055
transform 1 0 12192 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_79_118
timestamp 1621261055
transform 1 0 12480 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_126
timestamp 1621261055
transform 1 0 13248 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_72
timestamp 1621261055
transform -1 0 13824 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output442
timestamp 1621261055
transform -1 0 14208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1006
timestamp 1621261055
transform 1 0 16992 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_136
timestamp 1621261055
transform 1 0 14208 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_144
timestamp 1621261055
transform 1 0 14976 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_152
timestamp 1621261055
transform 1 0 15744 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_160
timestamp 1621261055
transform 1 0 16512 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_164
timestamp 1621261055
transform 1 0 16896 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output409
timestamp 1621261055
transform 1 0 20160 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_166
timestamp 1621261055
transform 1 0 17088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_174
timestamp 1621261055
transform 1 0 17856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_182
timestamp 1621261055
transform 1 0 18624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_190
timestamp 1621261055
transform 1 0 19392 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1007
timestamp 1621261055
transform 1 0 22272 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output411
timestamp 1621261055
transform -1 0 23712 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_39
timestamp 1621261055
transform -1 0 23328 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_202
timestamp 1621261055
transform 1 0 20544 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_210
timestamp 1621261055
transform 1 0 21312 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_218
timestamp 1621261055
transform 1 0 22080 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_221
timestamp 1621261055
transform 1 0 22368 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output412
timestamp 1621261055
transform 1 0 24864 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_41
timestamp 1621261055
transform 1 0 24672 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_235
timestamp 1621261055
transform 1 0 23712 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_243
timestamp 1621261055
transform 1 0 24480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_251
timestamp 1621261055
transform 1 0 25248 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_259
timestamp 1621261055
transform 1 0 26016 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1008
timestamp 1621261055
transform 1 0 27552 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_267
timestamp 1621261055
transform 1 0 26784 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_276
timestamp 1621261055
transform 1 0 27648 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_284
timestamp 1621261055
transform 1 0 28416 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_292
timestamp 1621261055
transform 1 0 29184 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1009
timestamp 1621261055
transform 1 0 32832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_300
timestamp 1621261055
transform 1 0 29952 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_308
timestamp 1621261055
transform 1 0 30720 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_316
timestamp 1621261055
transform 1 0 31488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_324
timestamp 1621261055
transform 1 0 32256 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_328
timestamp 1621261055
transform 1 0 32640 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_331
timestamp 1621261055
transform 1 0 32928 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_339
timestamp 1621261055
transform 1 0 33696 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_347
timestamp 1621261055
transform 1 0 34464 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_355
timestamp 1621261055
transform 1 0 35232 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_363
timestamp 1621261055
transform 1 0 36000 0 1 55278
box -38 -49 806 715
use HAX1  HAX1
timestamp 1623610208
transform 1 0 38784 0 1 55278
box 0 -48 3168 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1010
timestamp 1621261055
transform 1 0 38112 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_371
timestamp 1621261055
transform 1 0 36768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_379
timestamp 1621261055
transform 1 0 37536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_383
timestamp 1621261055
transform 1 0 37920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_386
timestamp 1621261055
transform 1 0 38208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_390
timestamp 1621261055
transform 1 0 38592 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output424
timestamp 1621261055
transform 1 0 42336 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_425
timestamp 1621261055
transform 1 0 41952 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1011
timestamp 1621261055
transform 1 0 43392 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output426
timestamp 1621261055
transform -1 0 45792 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_56
timestamp 1621261055
transform -1 0 45408 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_433
timestamp 1621261055
transform 1 0 42720 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_437
timestamp 1621261055
transform 1 0 43104 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_439
timestamp 1621261055
transform 1 0 43296 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_441
timestamp 1621261055
transform 1 0 43488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_449
timestamp 1621261055
transform 1 0 44256 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_457
timestamp 1621261055
transform 1 0 45024 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1012
timestamp 1621261055
transform 1 0 48672 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output427
timestamp 1621261055
transform -1 0 47328 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_58
timestamp 1621261055
transform -1 0 46944 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_59
timestamp 1621261055
transform -1 0 47520 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_465
timestamp 1621261055
transform 1 0 45792 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_473
timestamp 1621261055
transform 1 0 46560 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_483
timestamp 1621261055
transform 1 0 47520 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_491
timestamp 1621261055
transform 1 0 48288 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output431
timestamp 1621261055
transform 1 0 51744 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_496
timestamp 1621261055
transform 1 0 48768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_504
timestamp 1621261055
transform 1 0 49536 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_512
timestamp 1621261055
transform 1 0 50304 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_520
timestamp 1621261055
transform 1 0 51072 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_524
timestamp 1621261055
transform 1 0 51456 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_526
timestamp 1621261055
transform 1 0 51648 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1013
timestamp 1621261055
transform 1 0 53952 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_531
timestamp 1621261055
transform 1 0 52128 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_539
timestamp 1621261055
transform 1 0 52896 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_547
timestamp 1621261055
transform 1 0 53664 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_549
timestamp 1621261055
transform 1 0 53856 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_551
timestamp 1621261055
transform 1 0 54048 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_559
timestamp 1621261055
transform 1 0 54816 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_32
timestamp 1621261055
transform -1 0 55776 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _035_
timestamp 1621261055
transform -1 0 56064 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_79_572
timestamp 1621261055
transform 1 0 56064 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_580
timestamp 1621261055
transform 1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output434
timestamp 1621261055
transform 1 0 56448 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_584
timestamp 1621261055
transform 1 0 57216 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_26
timestamp 1621261055
transform -1 0 57504 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output397
timestamp 1621261055
transform -1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_593
timestamp 1621261055
transform 1 0 58080 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_27
timestamp 1621261055
transform -1 0 58080 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_159
timestamp 1621261055
transform -1 0 58848 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_8
timestamp 1621261055
transform 1 0 1920 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output368
timestamp 1621261055
transform 1 0 1536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_160
timestamp 1621261055
transform 1 0 1152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_16
timestamp 1621261055
transform 1 0 2688 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output417
timestamp 1621261055
transform 1 0 2784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_25
timestamp 1621261055
transform 1 0 3552 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_21
timestamp 1621261055
transform 1 0 3168 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_29
timestamp 1621261055
transform 1 0 3936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_27
timestamp 1621261055
transform 1 0 3744 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_17
timestamp 1621261055
transform 1 0 4128 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output390
timestamp 1621261055
transform 1 0 4320 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1014
timestamp 1621261055
transform 1 0 3840 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_41
timestamp 1621261055
transform 1 0 5088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_37
timestamp 1621261055
transform 1 0 4704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_48
timestamp 1621261055
transform 1 0 5760 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_43
timestamp 1621261055
transform 1 0 5280 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output399
timestamp 1621261055
transform 1 0 5376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_56
timestamp 1621261055
transform 1 0 6528 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output437
timestamp 1621261055
transform 1 0 6144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_65
timestamp 1621261055
transform 1 0 7392 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_80_60
timestamp 1621261055
transform 1 0 6912 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output400
timestamp 1621261055
transform 1 0 7008 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1015
timestamp 1621261055
transform 1 0 9120 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output401
timestamp 1621261055
transform 1 0 8352 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output402
timestamp 1621261055
transform 1 0 10176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_29
timestamp 1621261055
transform 1 0 9984 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_73
timestamp 1621261055
transform 1 0 8160 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_79
timestamp 1621261055
transform 1 0 8736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_84
timestamp 1621261055
transform 1 0 9216 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_98
timestamp 1621261055
transform 1 0 10560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output440
timestamp 1621261055
transform 1 0 10944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_106
timestamp 1621261055
transform 1 0 11328 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_31
timestamp 1621261055
transform 1 0 11520 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output403
timestamp 1621261055
transform 1 0 11712 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_114
timestamp 1621261055
transform 1 0 12096 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_70
timestamp 1621261055
transform 1 0 12288 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output441
timestamp 1621261055
transform 1 0 12480 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_122
timestamp 1621261055
transform 1 0 12864 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_126
timestamp 1621261055
transform 1 0 13248 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output404
timestamp 1621261055
transform 1 0 13344 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_131
timestamp 1621261055
transform 1 0 13728 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_139
timestamp 1621261055
transform 1 0 14496 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_137
timestamp 1621261055
transform 1 0 14304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_135
timestamp 1621261055
transform 1 0 14112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1016
timestamp 1621261055
transform 1 0 14400 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_147
timestamp 1621261055
transform 1 0 15264 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output405
timestamp 1621261055
transform 1 0 14880 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_155
timestamp 1621261055
transform 1 0 16032 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output443
timestamp 1621261055
transform 1 0 15648 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_35
timestamp 1621261055
transform 1 0 16800 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output407
timestamp 1621261055
transform 1 0 16992 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1017
timestamp 1621261055
transform 1 0 19680 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output371
timestamp 1621261055
transform 1 0 20160 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output408
timestamp 1621261055
transform 1 0 18528 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_169
timestamp 1621261055
transform 1 0 17376 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_177
timestamp 1621261055
transform 1 0 18144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_185
timestamp 1621261055
transform 1 0 18912 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_194
timestamp 1621261055
transform 1 0 19776 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_206
timestamp 1621261055
transform 1 0 20928 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_202
timestamp 1621261055
transform 1 0 20544 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_213
timestamp 1621261055
transform 1 0 21600 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_208
timestamp 1621261055
transform 1 0 21120 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_37
timestamp 1621261055
transform -1 0 21984 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output372
timestamp 1621261055
transform 1 0 21216 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_221
timestamp 1621261055
transform 1 0 22368 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output410
timestamp 1621261055
transform -1 0 22368 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_229
timestamp 1621261055
transform 1 0 23136 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output373
timestamp 1621261055
transform 1 0 22752 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1018
timestamp 1621261055
transform 1 0 24960 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output374
timestamp 1621261055
transform 1 0 24192 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output375
timestamp 1621261055
transform 1 0 25920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_237
timestamp 1621261055
transform 1 0 23904 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_239
timestamp 1621261055
transform 1 0 24096 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_244
timestamp 1621261055
transform 1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_249
timestamp 1621261055
transform 1 0 25056 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_80_257
timestamp 1621261055
transform 1 0 25824 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_262
timestamp 1621261055
transform 1 0 26304 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output413
timestamp 1621261055
transform 1 0 26688 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_270
timestamp 1621261055
transform 1 0 27072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_274
timestamp 1621261055
transform 1 0 27456 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output376
timestamp 1621261055
transform 1 0 27552 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_279
timestamp 1621261055
transform 1 0 27936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_43
timestamp 1621261055
transform -1 0 28320 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output414
timestamp 1621261055
transform -1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_287
timestamp 1621261055
transform 1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_291
timestamp 1621261055
transform 1 0 29088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_45
timestamp 1621261055
transform -1 0 29472 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output415
timestamp 1621261055
transform -1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1019
timestamp 1621261055
transform 1 0 30240 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output378
timestamp 1621261055
transform 1 0 30720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output380
timestamp 1621261055
transform 1 0 32256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output416
timestamp 1621261055
transform 1 0 31488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_299
timestamp 1621261055
transform 1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_304
timestamp 1621261055
transform 1 0 30336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_312
timestamp 1621261055
transform 1 0 31104 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_320
timestamp 1621261055
transform 1 0 31872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_328
timestamp 1621261055
transform 1 0 32640 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output418
timestamp 1621261055
transform 1 0 33024 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_336
timestamp 1621261055
transform 1 0 33408 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_7
timestamp 1621261055
transform 1 0 33600 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_344
timestamp 1621261055
transform 1 0 34176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output381
timestamp 1621261055
transform 1 0 33792 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_47
timestamp 1621261055
transform -1 0 34560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output419
timestamp 1621261055
transform -1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_354
timestamp 1621261055
transform 1 0 35136 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_48
timestamp 1621261055
transform -1 0 35136 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1020
timestamp 1621261055
transform 1 0 35520 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_359
timestamp 1621261055
transform 1 0 35616 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output382
timestamp 1621261055
transform 1 0 36000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_367
timestamp 1621261055
transform 1 0 36384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_50
timestamp 1621261055
transform -1 0 36768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output420
timestamp 1621261055
transform -1 0 37152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_375
timestamp 1621261055
transform 1 0 37152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_52
timestamp 1621261055
transform 1 0 37344 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output421
timestamp 1621261055
transform 1 0 37536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_387
timestamp 1621261055
transform 1 0 38304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_383
timestamp 1621261055
transform 1 0 37920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_9
timestamp 1621261055
transform -1 0 38592 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_394
timestamp 1621261055
transform 1 0 38976 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output384
timestamp 1621261055
transform -1 0 38976 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_404
timestamp 1621261055
transform 1 0 39936 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_402
timestamp 1621261055
transform 1 0 39744 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output385
timestamp 1621261055
transform 1 0 40032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_409
timestamp 1621261055
transform 1 0 40416 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_414
timestamp 1621261055
transform 1 0 40896 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1021
timestamp 1621261055
transform 1 0 40800 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_80_420
timestamp 1621261055
transform 1 0 41472 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_418
timestamp 1621261055
transform 1 0 41280 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_11
timestamp 1621261055
transform -1 0 41760 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output386
timestamp 1621261055
transform -1 0 42144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_427
timestamp 1621261055
transform 1 0 42144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_435
timestamp 1621261055
transform 1 0 42912 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_13
timestamp 1621261055
transform -1 0 43296 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output423
timestamp 1621261055
transform 1 0 42528 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_443
timestamp 1621261055
transform 1 0 43680 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_54
timestamp 1621261055
transform -1 0 44064 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output387
timestamp 1621261055
transform -1 0 43680 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_453
timestamp 1621261055
transform 1 0 44640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_451
timestamp 1621261055
transform 1 0 44448 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_15
timestamp 1621261055
transform 1 0 44736 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output425
timestamp 1621261055
transform -1 0 44448 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_460
timestamp 1621261055
transform 1 0 45312 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output388
timestamp 1621261055
transform 1 0 44928 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1022
timestamp 1621261055
transform 1 0 46080 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output389
timestamp 1621261055
transform 1 0 46560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output391
timestamp 1621261055
transform -1 0 48384 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_19
timestamp 1621261055
transform -1 0 48000 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_20
timestamp 1621261055
transform -1 0 48576 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_61
timestamp 1621261055
transform -1 0 48768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_469
timestamp 1621261055
transform 1 0 46176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_477
timestamp 1621261055
transform 1 0 46944 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_80_485
timestamp 1621261055
transform 1 0 47712 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output429
timestamp 1621261055
transform -1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_504
timestamp 1621261055
transform 1 0 49536 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_500
timestamp 1621261055
transform 1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_509
timestamp 1621261055
transform 1 0 50016 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output392
timestamp 1621261055
transform 1 0 49632 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_63
timestamp 1621261055
transform -1 0 50400 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output430
timestamp 1621261055
transform -1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_517
timestamp 1621261055
transform 1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_521
timestamp 1621261055
transform 1 0 51168 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1023
timestamp 1621261055
transform 1 0 51360 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_524
timestamp 1621261055
transform 1 0 51456 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_22
timestamp 1621261055
transform -1 0 51840 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output393
timestamp 1621261055
transform -1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_532
timestamp 1621261055
transform 1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_536
timestamp 1621261055
transform 1 0 52608 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_542
timestamp 1621261055
transform 1 0 53184 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output394
timestamp 1621261055
transform 1 0 52800 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_64
timestamp 1621261055
transform -1 0 53568 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output432
timestamp 1621261055
transform -1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_550
timestamp 1621261055
transform 1 0 53952 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_24
timestamp 1621261055
transform 1 0 54144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output395
timestamp 1621261055
transform 1 0 54336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_558
timestamp 1621261055
transform 1 0 54720 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_65
timestamp 1621261055
transform -1 0 55104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1024
timestamp 1621261055
transform 1 0 56640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input31
timestamp 1621261055
transform 1 0 57696 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output396
timestamp 1621261055
transform 1 0 55872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output433
timestamp 1621261055
transform -1 0 55488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_566
timestamp 1621261055
transform 1 0 55488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_574
timestamp 1621261055
transform 1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_579
timestamp 1621261055
transform 1 0 56736 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_587
timestamp 1621261055
transform 1 0 57504 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_593
timestamp 1621261055
transform 1 0 58080 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_161
timestamp 1621261055
transform -1 0 58848 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_162
timestamp 1621261055
transform 1 0 1152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1025
timestamp 1621261055
transform 1 0 3840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input1
timestamp 1621261055
transform 1 0 1536 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input12
timestamp 1621261055
transform 1 0 2304 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input23
timestamp 1621261055
transform 1 0 3072 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_8
timestamp 1621261055
transform 1 0 1920 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_16
timestamp 1621261055
transform 1 0 2688 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_24
timestamp 1621261055
transform 1 0 3456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_29
timestamp 1621261055
transform 1 0 3936 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_37
timestamp 1621261055
transform 1 0 4704 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input32
timestamp 1621261055
transform 1 0 4896 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_43
timestamp 1621261055
transform 1 0 5280 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_5
timestamp 1621261055
transform 1 0 5472 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output379
timestamp 1621261055
transform 1 0 5664 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_51
timestamp 1621261055
transform 1 0 6048 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_57
timestamp 1621261055
transform 1 0 6624 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_55
timestamp 1621261055
transform 1 0 6432 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1026
timestamp 1621261055
transform 1 0 6528 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_1  input33
timestamp 1621261055
transform 1 0 7008 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_65
timestamp 1621261055
transform 1 0 7392 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1027
timestamp 1621261055
transform 1 0 9216 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input34
timestamp 1621261055
transform 1 0 8064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input35
timestamp 1621261055
transform 1 0 9696 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_69
timestamp 1621261055
transform 1 0 7776 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_71
timestamp 1621261055
transform 1 0 7968 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_76
timestamp 1621261055
transform 1 0 8448 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_85
timestamp 1621261055
transform 1 0 9312 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_93
timestamp 1621261055
transform 1 0 10080 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_103
timestamp 1621261055
transform 1 0 11040 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_101
timestamp 1621261055
transform 1 0 10848 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input36
timestamp 1621261055
transform 1 0 11136 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_113
timestamp 1621261055
transform 1 0 12000 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_108
timestamp 1621261055
transform 1 0 11520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1028
timestamp 1621261055
transform 1 0 11904 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_125
timestamp 1621261055
transform 1 0 13152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input37
timestamp 1621261055
transform 1 0 12768 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_129
timestamp 1621261055
transform 1 0 13536 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_1
timestamp 1621261055
transform 1 0 13632 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output369
timestamp 1621261055
transform 1 0 13824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1029
timestamp 1621261055
transform 1 0 14592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  input2
timestamp 1621261055
transform 1 0 15936 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input38
timestamp 1621261055
transform 1 0 15072 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_136
timestamp 1621261055
transform 1 0 14208 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_141
timestamp 1621261055
transform 1 0 14688 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_149
timestamp 1621261055
transform 1 0 15456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_153
timestamp 1621261055
transform 1 0 15840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_158
timestamp 1621261055
transform 1 0 16320 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_169
timestamp 1621261055
transform 1 0 17376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_166
timestamp 1621261055
transform 1 0 17088 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  input3
timestamp 1621261055
transform 1 0 17760 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1030
timestamp 1621261055
transform 1 0 17280 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_177
timestamp 1621261055
transform 1 0 18144 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_191
timestamp 1621261055
transform 1 0 19488 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_185
timestamp 1621261055
transform 1 0 18912 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  input4
timestamp 1621261055
transform 1 0 19104 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_197
timestamp 1621261055
transform 1 0 20064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_195
timestamp 1621261055
transform 1 0 19872 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1031
timestamp 1621261055
transform 1 0 19968 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1032
timestamp 1621261055
transform 1 0 22656 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input5
timestamp 1621261055
transform 1 0 20640 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input6
timestamp 1621261055
transform 1 0 23136 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output370
timestamp 1621261055
transform 1 0 21504 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_3
timestamp 1621261055
transform 1 0 21312 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_201
timestamp 1621261055
transform 1 0 20448 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_208
timestamp 1621261055
transform 1 0 21120 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_216
timestamp 1621261055
transform 1 0 21888 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_225
timestamp 1621261055
transform 1 0 22752 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1033
timestamp 1621261055
transform 1 0 25344 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input7
timestamp 1621261055
transform 1 0 23904 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input8
timestamp 1621261055
transform 1 0 25824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_233
timestamp 1621261055
transform 1 0 23520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_241
timestamp 1621261055
transform 1 0 24288 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_249
timestamp 1621261055
transform 1 0 25056 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_251
timestamp 1621261055
transform 1 0 25248 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_253
timestamp 1621261055
transform 1 0 25440 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_261
timestamp 1621261055
transform 1 0 26208 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1034
timestamp 1621261055
transform 1 0 28032 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input9
timestamp 1621261055
transform 1 0 26976 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input10
timestamp 1621261055
transform 1 0 28608 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_273
timestamp 1621261055
transform 1 0 27360 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_277
timestamp 1621261055
transform 1 0 27744 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_279
timestamp 1621261055
transform 1 0 27936 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_281
timestamp 1621261055
transform 1 0 28128 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_285
timestamp 1621261055
transform 1 0 28512 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_290
timestamp 1621261055
transform 1 0 28992 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_304
timestamp 1621261055
transform 1 0 30336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_298
timestamp 1621261055
transform 1 0 29760 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input11
timestamp 1621261055
transform 1 0 29952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_309
timestamp 1621261055
transform 1 0 30816 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1035
timestamp 1621261055
transform 1 0 30720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_322
timestamp 1621261055
transform 1 0 32064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_317
timestamp 1621261055
transform 1 0 31584 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input13
timestamp 1621261055
transform 1 0 31680 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_330
timestamp 1621261055
transform 1 0 32832 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output377
timestamp 1621261055
transform 1 0 32448 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1036
timestamp 1621261055
transform 1 0 33408 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input14
timestamp 1621261055
transform 1 0 33888 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input15
timestamp 1621261055
transform 1 0 34848 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_334
timestamp 1621261055
transform 1 0 33216 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_337
timestamp 1621261055
transform 1 0 33504 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_346
timestamp 1621261055
transform 1 0 34368 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_350
timestamp 1621261055
transform 1 0 34752 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_355
timestamp 1621261055
transform 1 0 35232 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_363
timestamp 1621261055
transform 1 0 36000 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_365
timestamp 1621261055
transform 1 0 36192 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input16
timestamp 1621261055
transform 1 0 36576 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1037
timestamp 1621261055
transform 1 0 36096 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_373
timestamp 1621261055
transform 1 0 36960 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_388
timestamp 1621261055
transform 1 0 38400 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_383
timestamp 1621261055
transform 1 0 37920 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_381
timestamp 1621261055
transform 1 0 37728 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input17
timestamp 1621261055
transform 1 0 38016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_393
timestamp 1621261055
transform 1 0 38880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1038
timestamp 1621261055
transform 1 0 38784 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1039
timestamp 1621261055
transform 1 0 41472 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input18 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 39648 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input19
timestamp 1621261055
transform 1 0 41952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output383
timestamp 1621261055
transform 1 0 40608 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_407
timestamp 1621261055
transform 1 0 40224 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_415
timestamp 1621261055
transform 1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_419
timestamp 1621261055
transform 1 0 41376 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_421
timestamp 1621261055
transform 1 0 41568 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_429
timestamp 1621261055
transform 1 0 42336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1040
timestamp 1621261055
transform 1 0 44160 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input20
timestamp 1621261055
transform 1 0 42816 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input21
timestamp 1621261055
transform 1 0 44640 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_433
timestamp 1621261055
transform 1 0 42720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_439
timestamp 1621261055
transform 1 0 43296 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_447
timestamp 1621261055
transform 1 0 44064 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_449
timestamp 1621261055
transform 1 0 44256 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_457
timestamp 1621261055
transform 1 0 45024 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1041
timestamp 1621261055
transform 1 0 46848 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input22
timestamp 1621261055
transform 1 0 45888 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input24
timestamp 1621261055
transform 1 0 47520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input25
timestamp 1621261055
transform 1 0 48672 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_1  FILLER_81_465
timestamp 1621261055
transform 1 0 45792 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_472
timestamp 1621261055
transform 1 0 46464 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_477
timestamp 1621261055
transform 1 0 46944 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_481
timestamp 1621261055
transform 1 0 47328 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_487
timestamp 1621261055
transform 1 0 47904 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1042
timestamp 1621261055
transform 1 0 49536 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input26
timestamp 1621261055
transform 1 0 50688 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_500
timestamp 1621261055
transform 1 0 49152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_505
timestamp 1621261055
transform 1 0 49632 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_513
timestamp 1621261055
transform 1 0 50400 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_515
timestamp 1621261055
transform 1 0 50592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_521
timestamp 1621261055
transform 1 0 51168 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_533
timestamp 1621261055
transform 1 0 52320 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_531
timestamp 1621261055
transform 1 0 52128 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_529
timestamp 1621261055
transform 1 0 51936 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1043
timestamp 1621261055
transform 1 0 52224 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input27
timestamp 1621261055
transform 1 0 52704 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_547
timestamp 1621261055
transform 1 0 53664 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_543
timestamp 1621261055
transform 1 0 53280 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_553
timestamp 1621261055
transform 1 0 54240 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input28
timestamp 1621261055
transform 1 0 53856 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_561
timestamp 1621261055
transform 1 0 55008 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_559
timestamp 1621261055
transform 1 0 54816 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_557
timestamp 1621261055
transform 1 0 54624 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1044
timestamp 1621261055
transform 1 0 54912 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1045
timestamp 1621261055
transform 1 0 57600 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_1  input29
timestamp 1621261055
transform 1 0 55392 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  input30
timestamp 1621261055
transform 1 0 56832 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_569
timestamp 1621261055
transform 1 0 55776 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_577
timestamp 1621261055
transform 1 0 56544 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_579
timestamp 1621261055
transform 1 0 56736 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_584
timestamp 1621261055
transform 1 0 57216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_589
timestamp 1621261055
transform 1 0 57696 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_163
timestamp 1621261055
transform -1 0 58848 0 1 56610
box -38 -49 422 715
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 114 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 115 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 116 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 117 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 118 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 119 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 120 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 121 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 122 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 123 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 124 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 125 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 126 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 127 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 128 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 129 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 130 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 131 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 132 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 133 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 134 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 135 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 136 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 137 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 138 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 139 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 140 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 141 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 142 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 143 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 144 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 145 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 146 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 147 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 148 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 149 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 150 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 151 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 152 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 153 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 154 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 155 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 156 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 157 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 158 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 159 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 160 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 161 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 162 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 163 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 164 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 165 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 166 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 167 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 168 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 169 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 170 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 171 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 172 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 173 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 174 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 175 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 176 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 177 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 178 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 179 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 180 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 181 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 182 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 183 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 184 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 185 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 186 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 187 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 188 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 189 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 190 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 191 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 192 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 193 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 194 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 195 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 196 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 197 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 198 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 199 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 200 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 201 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 202 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 203 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 204 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 205 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 206 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 207 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 208 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 209 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 210 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 211 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 212 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 213 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 214 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 215 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 216 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 217 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 218 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 219 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 220 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 221 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 222 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 223 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 224 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 225 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 226 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 227 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 228 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 229 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 230 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 231 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 232 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 233 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 234 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 235 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 236 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 237 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 238 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 239 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 240 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 241 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 242 nsew signal tristate
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 243 nsew signal tristate
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 244 nsew signal tristate
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 245 nsew signal tristate
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 246 nsew signal tristate
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 247 nsew signal tristate
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 248 nsew signal tristate
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 249 nsew signal tristate
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 250 nsew signal tristate
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 251 nsew signal tristate
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 252 nsew signal tristate
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 253 nsew signal tristate
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 254 nsew signal tristate
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 255 nsew signal tristate
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 256 nsew signal tristate
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 257 nsew signal tristate
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 258 nsew signal tristate
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 259 nsew signal tristate
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 260 nsew signal tristate
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 261 nsew signal tristate
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 262 nsew signal tristate
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 263 nsew signal tristate
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 264 nsew signal tristate
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 265 nsew signal tristate
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 266 nsew signal tristate
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 267 nsew signal tristate
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 268 nsew signal tristate
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 269 nsew signal tristate
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 270 nsew signal tristate
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 271 nsew signal tristate
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 272 nsew signal tristate
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 273 nsew signal tristate
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 274 nsew signal tristate
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 275 nsew signal tristate
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 276 nsew signal tristate
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 277 nsew signal tristate
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 278 nsew signal tristate
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 279 nsew signal tristate
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 280 nsew signal tristate
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 281 nsew signal tristate
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 282 nsew signal tristate
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 283 nsew signal tristate
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 284 nsew signal tristate
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 285 nsew signal tristate
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 286 nsew signal tristate
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 287 nsew signal tristate
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 288 nsew signal tristate
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 289 nsew signal tristate
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 290 nsew signal tristate
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 291 nsew signal tristate
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 292 nsew signal tristate
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 293 nsew signal tristate
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 294 nsew signal tristate
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 295 nsew signal tristate
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 296 nsew signal tristate
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 297 nsew signal tristate
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 298 nsew signal tristate
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 299 nsew signal tristate
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 300 nsew signal tristate
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 301 nsew signal tristate
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 302 nsew signal tristate
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 303 nsew signal tristate
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 304 nsew signal tristate
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 305 nsew signal tristate
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 306 nsew signal tristate
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 307 nsew signal tristate
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 308 nsew signal tristate
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 309 nsew signal tristate
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 310 nsew signal tristate
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 311 nsew signal tristate
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 312 nsew signal tristate
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 313 nsew signal tristate
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 314 nsew signal tristate
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 315 nsew signal tristate
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 316 nsew signal tristate
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 317 nsew signal tristate
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 318 nsew signal tristate
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 319 nsew signal tristate
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 320 nsew signal tristate
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 321 nsew signal tristate
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 322 nsew signal tristate
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 323 nsew signal tristate
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 324 nsew signal tristate
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 325 nsew signal tristate
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 326 nsew signal tristate
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 327 nsew signal tristate
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 328 nsew signal tristate
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 329 nsew signal tristate
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 330 nsew signal tristate
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 331 nsew signal tristate
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 332 nsew signal tristate
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 333 nsew signal tristate
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 334 nsew signal tristate
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 335 nsew signal tristate
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 336 nsew signal tristate
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 337 nsew signal tristate
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 338 nsew signal tristate
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 339 nsew signal tristate
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 340 nsew signal tristate
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 341 nsew signal tristate
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 342 nsew signal tristate
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 343 nsew signal tristate
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 344 nsew signal tristate
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 345 nsew signal tristate
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 346 nsew signal tristate
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 347 nsew signal tristate
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 348 nsew signal tristate
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 349 nsew signal tristate
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 350 nsew signal tristate
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 351 nsew signal tristate
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 352 nsew signal tristate
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 353 nsew signal tristate
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 354 nsew signal tristate
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 355 nsew signal tristate
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 356 nsew signal tristate
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 357 nsew signal tristate
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 358 nsew signal tristate
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 359 nsew signal tristate
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 360 nsew signal tristate
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 361 nsew signal tristate
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 362 nsew signal tristate
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 363 nsew signal tristate
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 364 nsew signal tristate
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 365 nsew signal tristate
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 366 nsew signal tristate
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 367 nsew signal tristate
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 368 nsew signal tristate
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 369 nsew signal tristate
rlabel metal2 s 13172 0 13228 800 6 la_oen[0]
port 370 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oen[100]
port 371 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oen[101]
port 372 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oen[102]
port 373 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oen[103]
port 374 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oen[104]
port 375 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oen[105]
port 376 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oen[106]
port 377 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oen[107]
port 378 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oen[108]
port 379 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oen[109]
port 380 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oen[10]
port 381 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oen[110]
port 382 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oen[111]
port 383 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oen[112]
port 384 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oen[113]
port 385 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oen[114]
port 386 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oen[115]
port 387 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oen[116]
port 388 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oen[117]
port 389 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oen[118]
port 390 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oen[119]
port 391 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oen[120]
port 393 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oen[121]
port 394 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oen[122]
port 395 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oen[123]
port 396 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oen[124]
port 397 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oen[125]
port 398 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oen[126]
port 399 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oen[127]
port 400 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oen[12]
port 401 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oen[13]
port 402 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oen[14]
port 403 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oen[15]
port 404 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oen[16]
port 405 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oen[18]
port 407 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oen[19]
port 408 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oen[1]
port 409 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oen[20]
port 410 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oen[21]
port 411 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oen[22]
port 412 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oen[24]
port 414 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oen[25]
port 415 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oen[26]
port 416 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oen[27]
port 417 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oen[28]
port 418 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oen[2]
port 420 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oen[30]
port 421 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oen[31]
port 422 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oen[32]
port 423 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oen[33]
port 424 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oen[34]
port 425 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oen[36]
port 427 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oen[37]
port 428 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oen[38]
port 429 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oen[39]
port 430 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oen[3]
port 431 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oen[40]
port 432 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oen[42]
port 434 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oen[43]
port 435 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oen[44]
port 436 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oen[45]
port 437 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oen[46]
port 438 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oen[48]
port 440 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oen[49]
port 441 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oen[4]
port 442 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oen[50]
port 443 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oen[51]
port 444 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oen[52]
port 445 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oen[54]
port 447 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oen[55]
port 448 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oen[56]
port 449 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oen[57]
port 450 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oen[58]
port 451 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oen[60]
port 454 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oen[61]
port 455 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oen[62]
port 456 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oen[63]
port 457 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oen[64]
port 458 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oen[66]
port 460 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oen[67]
port 461 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oen[68]
port 462 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oen[69]
port 463 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oen[6]
port 464 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oen[70]
port 465 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oen[72]
port 467 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oen[73]
port 468 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oen[74]
port 469 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oen[75]
port 470 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oen[76]
port 471 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oen[78]
port 473 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oen[79]
port 474 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oen[7]
port 475 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oen[80]
port 476 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oen[81]
port 477 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oen[82]
port 478 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oen[84]
port 480 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oen[85]
port 481 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oen[86]
port 482 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oen[87]
port 483 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oen[88]
port 484 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oen[89]
port 485 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oen[8]
port 486 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oen[90]
port 487 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oen[91]
port 488 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oen[92]
port 489 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oen[93]
port 490 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oen[94]
port 491 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oen[95]
port 492 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oen[96]
port 493 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oen[97]
port 494 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oen[98]
port 495 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oen[99]
port 496 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oen[9]
port 497 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 498 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 499 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 500 nsew signal tristate
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 501 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 502 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 503 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 504 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 505 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 506 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 507 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 508 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 509 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 510 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 511 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 512 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 513 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 514 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 515 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 516 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 517 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 518 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 519 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 520 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 521 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 522 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 523 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 524 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 525 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 526 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 527 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 528 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 529 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 530 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 531 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 532 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 533 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 534 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 535 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 536 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 537 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 538 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 539 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 540 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 541 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 542 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 543 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 544 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 545 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 546 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 547 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 548 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 549 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 550 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 551 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 552 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 553 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 554 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 555 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 556 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 557 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 558 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 559 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 560 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 561 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 562 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 563 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 564 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 565 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 566 nsew signal tristate
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 567 nsew signal tristate
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 568 nsew signal tristate
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 569 nsew signal tristate
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 570 nsew signal tristate
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 571 nsew signal tristate
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 572 nsew signal tristate
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 573 nsew signal tristate
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 574 nsew signal tristate
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 575 nsew signal tristate
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 576 nsew signal tristate
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 577 nsew signal tristate
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 578 nsew signal tristate
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 579 nsew signal tristate
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 580 nsew signal tristate
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 581 nsew signal tristate
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 582 nsew signal tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew signal tristate
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 584 nsew signal tristate
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 585 nsew signal tristate
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 586 nsew signal tristate
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 587 nsew signal tristate
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 588 nsew signal tristate
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 589 nsew signal tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew signal tristate
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 591 nsew signal tristate
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 592 nsew signal tristate
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 593 nsew signal tristate
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 594 nsew signal tristate
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 595 nsew signal tristate
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 596 nsew signal tristate
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 597 nsew signal tristate
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 598 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 599 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 600 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 601 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 602 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 603 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 604 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 606 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 607 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 608 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 609 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 610 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 611 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 612 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 613 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 614 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 615 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 616 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 618 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 619 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
