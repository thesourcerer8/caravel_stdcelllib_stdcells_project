magic
tech sky130A
magscale 1 2
timestamp 1636962392
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2016 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
rect 1713 48 1743 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
rect 1713 450 1743 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 355 134 413 146
rect 355 132 367 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 1027 134 1085 146
rect 1027 132 1039 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 48 849 132
rect 879 100 1039 132
rect 1073 132 1085 134
rect 1507 134 1565 146
rect 1507 132 1519 134
rect 1073 100 1137 132
rect 879 48 1137 100
rect 1167 48 1425 132
rect 1455 100 1519 132
rect 1553 132 1565 134
rect 1795 134 1853 146
rect 1795 132 1807 134
rect 1553 100 1713 132
rect 1455 48 1713 100
rect 1743 100 1807 132
rect 1841 132 1853 134
rect 1841 100 1901 132
rect 1743 48 1901 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 127 485
rect 161 451 273 485
rect 115 450 273 451
rect 303 593 561 618
rect 303 559 367 593
rect 401 559 561 593
rect 303 450 561 559
rect 591 450 849 618
rect 879 566 1137 618
rect 879 532 943 566
rect 977 532 1137 566
rect 879 485 1137 532
rect 879 451 1039 485
rect 1073 451 1137 485
rect 879 450 1137 451
rect 1167 450 1425 618
rect 1455 593 1713 618
rect 1455 559 1519 593
rect 1553 559 1713 593
rect 1455 450 1713 559
rect 1743 485 1901 618
rect 1743 451 1807 485
rect 1841 451 1901 485
rect 1743 450 1901 451
rect 115 439 173 450
rect 1027 439 1085 450
rect 1795 439 1853 450
<< ndiffc >>
rect 127 100 161 134
rect 367 100 401 134
rect 1039 100 1073 134
rect 1519 100 1553 134
rect 1807 100 1841 134
<< pdiffc >>
rect 127 451 161 485
rect 367 559 401 593
rect 943 532 977 566
rect 1039 451 1073 485
rect 1519 559 1553 593
rect 1807 451 1841 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
rect 1713 22 1743 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 2016 683
rect 31 643 1985 649
rect 31 618 1469 643
rect 1603 618 1985 643
rect 351 593 417 618
rect 351 559 367 593
rect 401 559 417 593
rect 1503 593 1569 609
rect 351 543 417 559
rect 927 566 993 582
rect 927 532 943 566
rect 977 532 993 566
rect 1503 559 1519 593
rect 1553 559 1569 593
rect 1503 543 1569 559
rect 927 516 993 532
rect 111 485 177 501
rect 111 451 127 485
rect 161 451 177 485
rect 1027 485 1089 501
rect 1027 482 1039 485
rect 111 435 177 451
rect 1023 451 1039 482
rect 1073 451 1089 485
rect 1791 485 1857 501
rect 1791 452 1807 485
rect 1023 435 1089 451
rect 1795 451 1807 452
rect 1841 451 1857 485
rect 1795 435 1857 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 977 402
rect 831 352 897 368
rect 559 231 593 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 355 134 417 150
rect 355 131 367 134
rect 111 84 177 100
rect 351 100 367 131
rect 401 100 417 134
rect 943 134 977 368
rect 1039 150 1073 435
rect 1123 402 1185 418
rect 1123 401 1135 402
rect 1119 368 1135 401
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1119 215 1185 231
rect 1119 184 1135 215
rect 1123 181 1135 184
rect 1169 181 1185 215
rect 1123 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 184 1761 215
rect 1745 181 1757 184
rect 1695 165 1757 181
rect 1023 134 1089 150
rect 1023 100 1039 134
rect 1073 100 1089 134
rect 1507 134 1569 150
rect 1507 131 1519 134
rect 351 84 417 100
rect 1023 84 1089 100
rect 1503 100 1519 131
rect 1553 100 1569 134
rect 1503 84 1569 100
rect 1791 134 1857 150
rect 1791 100 1807 134
rect 1841 100 1857 134
rect 1791 84 1857 100
rect 367 48 401 84
rect 1519 48 1553 84
rect 31 17 1985 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 2016 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 367 559 401 593
rect 943 532 977 566
rect 1519 559 1553 593
rect 127 451 161 485
rect 1807 451 1841 485
rect 271 368 305 402
rect 559 368 593 402
rect 271 181 305 215
rect 847 181 881 215
rect 127 100 161 134
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 943 100 977 134
rect 1807 100 1841 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 2016 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 2016 683
rect 0 618 2016 649
rect 355 593 413 618
rect 355 559 367 593
rect 401 559 413 593
rect 1507 593 1565 618
rect 355 547 413 559
rect 931 566 989 578
rect 931 532 943 566
rect 977 532 989 566
rect 1507 559 1519 593
rect 1553 559 1565 593
rect 1507 547 1565 559
rect 931 520 989 532
rect 115 485 173 497
rect 115 451 127 485
rect 161 451 173 485
rect 1795 485 1853 497
rect 115 439 173 451
rect 562 454 1742 482
rect 130 146 158 439
rect 562 414 590 454
rect 1714 414 1742 454
rect 1795 451 1807 485
rect 1841 451 1853 485
rect 1795 439 1853 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 1123 402 1181 414
rect 1123 399 1135 402
rect 547 356 605 368
rect 850 371 1135 399
rect 274 227 302 356
rect 850 227 878 371
rect 1123 368 1135 371
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 1411 402 1469 414
rect 1411 368 1423 402
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1699 402 1757 414
rect 1699 368 1711 402
rect 1745 368 1757 402
rect 1699 356 1757 368
rect 1426 227 1454 356
rect 1714 227 1742 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 212 317 215
rect 835 215 893 227
rect 835 212 847 215
rect 305 184 847 212
rect 305 181 317 184
rect 259 169 317 181
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 1411 215 1469 227
rect 1411 181 1423 215
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 1699 215 1757 227
rect 1699 181 1711 215
rect 1745 181 1757 215
rect 1699 169 1757 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 131 173 134
rect 931 134 989 146
rect 931 131 943 134
rect 161 103 943 131
rect 161 100 173 103
rect 115 88 173 100
rect 931 100 943 103
rect 977 131 989 134
rect 1138 131 1166 169
rect 977 103 1166 131
rect 1426 131 1454 169
rect 1810 146 1838 439
rect 1795 134 1853 146
rect 1795 131 1807 134
rect 1426 103 1807 131
rect 977 100 989 103
rect 931 88 989 100
rect 1795 100 1807 103
rect 1841 100 1853 134
rect 1795 88 1853 100
rect 0 17 2016 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 2016 17
rect 0 -48 2016 -17
<< labels >>
rlabel metal1 0 618 2016 714 0 VPWR
port 3 se
rlabel metal1 0 618 2016 714 0 VPWR
port 3 se
rlabel metal1 0 -48 2016 48 0 VGND
port 2 se
rlabel metal1 0 -48 2016 48 0 VGND
port 2 se
rlabel metal1 931 520 989 578 0 Y
port 4 se
rlabel metal1 259 169 317 184 0 A
port 0 se
rlabel metal1 835 169 893 184 0 A
port 0 se
rlabel metal1 259 184 893 212 0 A
port 0 se
rlabel metal1 259 212 317 227 0 A
port 0 se
rlabel metal1 835 212 893 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 850 227 878 371 0 A
port 0 se
rlabel metal1 1123 356 1181 371 0 A
port 0 se
rlabel metal1 850 371 1181 399 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel metal1 1123 399 1181 414 0 A
port 0 se
rlabel metal1 1699 169 1757 227 0 B
port 1 se
rlabel metal1 1714 227 1742 356 0 B
port 1 se
rlabel metal1 547 356 605 414 0 B
port 1 se
rlabel metal1 1699 356 1757 414 0 B
port 1 se
rlabel metal1 562 414 590 454 0 B
port 1 se
rlabel metal1 1714 414 1742 454 0 B
port 1 se
rlabel metal1 562 454 1742 482 0 B
port 1 se
rlabel locali 0 -17 2016 17 4 VGND
port 2 se ground default abutment
rlabel locali 31 17 1985 48 4 VGND
port 2 se ground default abutment
rlabel locali 0 649 2016 683 4 VPWR
port 3 se power default abutment
rlabel metal1 31 618 1985 649 4 VGND
port 2 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2016 666
<< end >>
