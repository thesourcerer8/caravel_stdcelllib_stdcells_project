MACRO SUTHERLAND1989
 CLASS CORE ;
 FOREIGN SUTHERLAND1989 0 0 ;
 SIZE 11.52 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
    END
  END GND

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 7.77500000 0.84500000 8.06500000 0.92000000 ;
        RECT 9.93500000 0.84500000 10.22500000 0.92000000 ;
        RECT 7.77500000 0.92000000 10.22500000 1.06000000 ;
        RECT 7.77500000 1.06000000 8.06500000 1.13500000 ;
        RECT 9.93500000 1.06000000 10.22500000 1.13500000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 5.61500000 0.84500000 5.90500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 5.69000000 1.13500000 5.83000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 1.85500000 ;
        RECT 5.61500000 1.78000000 5.90500000 1.85500000 ;
        RECT 1.29500000 1.85500000 5.90500000 1.99500000 ;
        RECT 1.29500000 1.99500000 1.58500000 2.07000000 ;
        RECT 5.61500000 1.99500000 5.90500000 2.07000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 2.73500000 0.84500000 3.02500000 0.92000000 ;
        RECT 4.17500000 0.84500000 4.46500000 0.92000000 ;
        RECT 2.73500000 0.92000000 4.46500000 1.06000000 ;
        RECT 2.73500000 1.06000000 3.02500000 1.13500000 ;
        RECT 4.17500000 1.06000000 4.46500000 1.13500000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 9.99500000 0.90500000 10.16500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 9.99500000 1.84000000 10.16500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 5.19500000 2.25500000 5.36500000 2.42500000 ;
     RECT 7.83500000 2.25500000 8.00500000 2.42500000 ;
     RECT 9.27500000 2.25500000 9.44500000 2.42500000 ;
     RECT 10.47500000 2.25500000 10.64500000 2.42500000 ;
     RECT 3.27500000 2.79500000 3.44500000 2.96500000 ;
     RECT 6.15500000 2.79500000 6.32500000 2.96500000 ;

    LAYER ndiffc ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;
     RECT 5.19500000 0.50000000 5.36500000 0.67000000 ;
     RECT 6.15500000 0.50000000 6.32500000 0.67000000 ;
     RECT 7.83500000 0.50000000 8.00500000 0.67000000 ;
     RECT 9.27500000 0.50000000 9.44500000 0.67000000 ;
     RECT 10.47500000 0.50000000 10.64500000 0.67000000 ;

    LAYER li1 ;
     RECT 0.55500000 0.42000000 0.88500000 0.75000000 ;
     RECT 3.19500000 0.42000000 3.52500000 0.75000000 ;
     RECT 5.11500000 0.42000000 5.44500000 0.75000000 ;
     RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
     RECT 6.15500000 0.24000000 6.32500000 0.42000000 ;
     RECT 6.07500000 0.42000000 6.40500000 0.75000000 ;
     RECT 9.19500000 0.42000000 9.52500000 0.75000000 ;
     RECT 10.39500000 0.42000000 10.72500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 5.59500000 0.82500000 5.92500000 1.15500000 ;
     RECT 7.03500000 0.82500000 7.36500000 1.15500000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 2.79500000 1.15500000 2.96500000 1.76000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 4.15500000 0.82500000 4.48500000 1.15500000 ;
     RECT 4.23500000 1.15500000 4.40500000 1.76000000 ;
     RECT 4.15500000 1.76000000 4.48500000 2.09000000 ;
     RECT 5.59500000 1.76000000 5.92500000 2.09000000 ;
     RECT 7.03500000 1.76000000 7.36500000 2.09000000 ;
     RECT 9.91500000 0.82500000 10.24500000 1.15500000 ;
     RECT 9.99500000 1.15500000 10.16500000 1.76000000 ;
     RECT 9.91500000 1.76000000 10.24500000 2.09000000 ;
     RECT 0.55500000 2.17500000 0.88500000 2.50500000 ;
     RECT 5.11500000 2.17500000 5.44500000 2.50500000 ;
     RECT 7.75500000 0.42000000 8.08500000 0.75000000 ;
     RECT 7.83500000 0.75000000 8.00500000 2.17500000 ;
     RECT 7.75500000 2.17500000 8.08500000 2.50500000 ;
     RECT 9.19500000 2.17500000 9.52500000 2.50500000 ;
     RECT 10.39500000 2.17500000 10.72500000 2.50500000 ;
     RECT 3.19500000 2.71500000 3.52500000 3.04500000 ;
     RECT 6.07500000 2.71500000 6.40500000 3.04500000 ;
     RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;

    LAYER viali ;
     RECT 3.27500000 -0.08500000 3.44500000 0.08500000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;
     RECT 5.19500000 0.50000000 5.36500000 0.67000000 ;
     RECT 9.27500000 0.50000000 9.44500000 0.67000000 ;
     RECT 10.47500000 0.50000000 10.64500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 5.67500000 0.90500000 5.84500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 7.83500000 0.90500000 8.00500000 1.07500000 ;
     RECT 9.99500000 0.90500000 10.16500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 5.67500000 1.84000000 5.84500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 5.19500000 2.25500000 5.36500000 2.42500000 ;
     RECT 9.27500000 2.25500000 9.44500000 2.42500000 ;
     RECT 10.47500000 2.25500000 10.64500000 2.42500000 ;
     RECT 3.27500000 2.79500000 3.44500000 2.96500000 ;
     RECT 6.15500000 2.79500000 6.32500000 2.96500000 ;
     RECT 6.15500000 3.24500000 6.32500000 3.41500000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
     RECT 3.29000000 0.24000000 3.43000000 0.44000000 ;
     RECT 3.21500000 0.44000000 3.50500000 0.73000000 ;
     RECT 5.13500000 0.44000000 5.42500000 0.51500000 ;
     RECT 9.21500000 0.44000000 9.50500000 0.51500000 ;
     RECT 5.13500000 0.51500000 9.50500000 0.65500000 ;
     RECT 5.13500000 0.65500000 5.42500000 0.73000000 ;
     RECT 9.21500000 0.65500000 9.50500000 0.73000000 ;
     RECT 2.73500000 0.84500000 3.02500000 0.92000000 ;
     RECT 4.17500000 0.84500000 4.46500000 0.92000000 ;
     RECT 2.73500000 0.92000000 4.46500000 1.06000000 ;
     RECT 2.73500000 1.06000000 3.02500000 1.13500000 ;
     RECT 4.17500000 1.06000000 4.46500000 1.13500000 ;
     RECT 7.77500000 0.84500000 8.06500000 0.92000000 ;
     RECT 9.93500000 0.84500000 10.22500000 0.92000000 ;
     RECT 7.77500000 0.92000000 10.22500000 1.06000000 ;
     RECT 7.77500000 1.06000000 8.06500000 1.13500000 ;
     RECT 9.93500000 1.06000000 10.22500000 1.13500000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 5.61500000 0.84500000 5.90500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 5.69000000 1.13500000 5.83000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 1.85500000 ;
     RECT 5.61500000 1.78000000 5.90500000 1.85500000 ;
     RECT 1.29500000 1.85500000 5.90500000 1.99500000 ;
     RECT 1.29500000 1.99500000 1.58500000 2.07000000 ;
     RECT 5.61500000 1.99500000 5.90500000 2.07000000 ;
     RECT 0.57500000 0.44000000 0.86500000 0.73000000 ;
     RECT 0.65000000 0.73000000 0.79000000 2.19500000 ;
     RECT 0.57500000 2.19500000 0.86500000 2.48500000 ;
     RECT 5.13500000 2.19500000 5.42500000 2.27000000 ;
     RECT 9.21500000 2.19500000 9.50500000 2.27000000 ;
     RECT 5.13500000 2.27000000 9.50500000 2.41000000 ;
     RECT 5.13500000 2.41000000 5.42500000 2.48500000 ;
     RECT 9.21500000 2.41000000 9.50500000 2.48500000 ;
     RECT 10.41500000 0.44000000 10.70500000 0.73000000 ;
     RECT 7.05500000 0.84500000 7.34500000 1.13500000 ;
     RECT 7.13000000 1.13500000 7.27000000 1.78000000 ;
     RECT 7.05500000 1.78000000 7.34500000 1.85500000 ;
     RECT 10.49000000 0.73000000 10.63000000 1.85500000 ;
     RECT 7.05500000 1.85500000 10.63000000 1.99500000 ;
     RECT 7.05500000 1.99500000 7.34500000 2.07000000 ;
     RECT 10.49000000 1.99500000 10.63000000 2.19500000 ;
     RECT 10.41500000 2.19500000 10.70500000 2.48500000 ;
     RECT 3.21500000 2.73500000 3.50500000 3.09000000 ;
     RECT 6.09500000 2.73500000 6.38500000 3.09000000 ;
     RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;

 END
END SUTHERLAND1989
