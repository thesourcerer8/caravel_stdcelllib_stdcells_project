magic
tech sky130A
timestamp 1621277354
<< end >>
