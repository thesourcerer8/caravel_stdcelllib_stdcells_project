magic
tech sky130A
magscale 1 2
<<<<<<< HEAD
timestamp 1624954273
=======
timestamp 1631894554
>>>>>>> c5da9e9885e361d05dee2aa6303a69fc26423c8e
<< obsli1 >>
rect 1152 2647 58848 57293
<< obsm1 >>
<<<<<<< HEAD
rect 16 1417 59888 57325
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< obsm2 >>
rect 22 59144 156 59200
rect 324 59144 636 59200
rect 804 59144 1116 59200
rect 1284 59144 1692 59200
rect 1860 59144 2172 59200
rect 2340 59144 2748 59200
rect 2916 59144 3228 59200
rect 3396 59144 3804 59200
rect 3972 59144 4284 59200
rect 4452 59144 4860 59200
rect 5028 59144 5340 59200
rect 5508 59144 5916 59200
rect 6084 59144 6396 59200
rect 6564 59144 6972 59200
rect 7140 59144 7452 59200
rect 7620 59144 8028 59200
rect 8196 59144 8508 59200
rect 8676 59144 9084 59200
rect 9252 59144 9564 59200
rect 9732 59144 10140 59200
rect 10308 59144 10620 59200
rect 10788 59144 11196 59200
rect 11364 59144 11676 59200
rect 11844 59144 12252 59200
rect 12420 59144 12732 59200
rect 12900 59144 13308 59200
rect 13476 59144 13788 59200
rect 13956 59144 14364 59200
rect 14532 59144 14844 59200
rect 15012 59144 15324 59200
rect 15492 59144 15900 59200
rect 16068 59144 16380 59200
rect 16548 59144 16956 59200
rect 17124 59144 17436 59200
rect 17604 59144 18012 59200
rect 18180 59144 18492 59200
rect 18660 59144 19068 59200
rect 19236 59144 19548 59200
rect 19716 59144 20124 59200
rect 20292 59144 20604 59200
rect 20772 59144 21180 59200
rect 21348 59144 21660 59200
rect 21828 59144 22236 59200
rect 22404 59144 22716 59200
rect 22884 59144 23292 59200
rect 23460 59144 23772 59200
rect 23940 59144 24348 59200
rect 24516 59144 24828 59200
rect 24996 59144 25404 59200
rect 25572 59144 25884 59200
rect 26052 59144 26460 59200
rect 26628 59144 26940 59200
rect 27108 59144 27516 59200
rect 27684 59144 27996 59200
rect 28164 59144 28572 59200
rect 28740 59144 29052 59200
rect 29220 59144 29628 59200
rect 29796 59144 30108 59200
rect 30276 59144 30588 59200
rect 30756 59144 31164 59200
rect 31332 59144 31644 59200
rect 31812 59144 32220 59200
rect 32388 59144 32700 59200
rect 32868 59144 33276 59200
rect 33444 59144 33756 59200
rect 33924 59144 34332 59200
rect 34500 59144 34812 59200
rect 34980 59144 35388 59200
rect 35556 59144 35868 59200
rect 36036 59144 36444 59200
rect 36612 59144 36924 59200
rect 37092 59144 37500 59200
rect 37668 59144 37980 59200
rect 38148 59144 38556 59200
rect 38724 59144 39036 59200
rect 39204 59144 39612 59200
rect 39780 59144 40092 59200
rect 40260 59144 40668 59200
rect 40836 59144 41148 59200
rect 41316 59144 41724 59200
rect 41892 59144 42204 59200
rect 42372 59144 42780 59200
rect 42948 59144 43260 59200
rect 43428 59144 43836 59200
rect 44004 59144 44316 59200
rect 44484 59144 44892 59200
rect 45060 59144 45372 59200
rect 45540 59144 45852 59200
rect 46020 59144 46428 59200
rect 46596 59144 46908 59200
rect 47076 59144 47484 59200
rect 47652 59144 47964 59200
rect 48132 59144 48540 59200
rect 48708 59144 49020 59200
rect 49188 59144 49596 59200
rect 49764 59144 50076 59200
rect 50244 59144 50652 59200
rect 50820 59144 51132 59200
rect 51300 59144 51708 59200
rect 51876 59144 52188 59200
rect 52356 59144 52764 59200
rect 52932 59144 53244 59200
rect 53412 59144 53820 59200
rect 53988 59144 54300 59200
rect 54468 59144 54876 59200
rect 55044 59144 55356 59200
rect 55524 59144 55932 59200
rect 56100 59144 56412 59200
rect 56580 59144 56988 59200
rect 57156 59144 57468 59200
rect 57636 59144 58044 59200
rect 58212 59144 58524 59200
rect 58692 59144 59100 59200
rect 59268 59144 59580 59200
rect 59748 59144 59882 59200
rect 22 856 59882 59144
rect 420 800 444 856
rect 900 800 924 856
rect 1284 800 1308 856
rect 1764 800 1788 856
rect 2244 800 2268 856
rect 2628 800 2652 856
rect 3108 800 3132 856
rect 3588 800 3612 856
rect 3972 800 3996 856
rect 4452 800 4476 856
rect 4836 800 4860 856
rect 5316 800 5340 856
rect 5796 800 5820 856
rect 6180 800 6204 856
rect 6660 800 6684 856
rect 7140 800 7164 856
rect 7524 800 7548 856
rect 8004 800 8028 856
rect 8388 800 8412 856
rect 8868 800 8892 856
rect 9348 800 9372 856
rect 9732 800 9756 856
rect 10212 800 10236 856
rect 10692 800 10716 856
rect 11076 800 11100 856
rect 11556 800 11580 856
rect 11940 800 11964 856
rect 12420 800 12444 856
rect 12900 800 12924 856
rect 13284 800 13308 856
rect 13764 800 13788 856
rect 14244 800 14268 856
rect 14628 800 14652 856
rect 15108 800 15132 856
rect 15588 800 15612 856
rect 15972 800 15996 856
rect 16452 800 16476 856
rect 16836 800 16860 856
rect 17316 800 17340 856
rect 17796 800 17820 856
rect 18180 800 18204 856
rect 18660 800 18684 856
rect 19140 800 19164 856
rect 19524 800 19548 856
rect 20004 800 20028 856
rect 20388 800 20412 856
rect 20868 800 20892 856
rect 21348 800 21372 856
rect 21732 800 21756 856
rect 22212 800 22236 856
rect 22692 800 22716 856
rect 23076 800 23100 856
rect 23556 800 23580 856
rect 23940 800 23964 856
rect 24420 800 24444 856
rect 24900 800 24924 856
rect 25284 800 25308 856
rect 25764 800 25788 856
rect 26244 800 26268 856
rect 26628 800 26652 856
rect 27108 800 27132 856
rect 27588 800 27612 856
rect 27972 800 27996 856
rect 28452 800 28476 856
rect 28836 800 28860 856
rect 29316 800 29340 856
rect 29796 800 29820 856
rect 30180 800 30204 856
rect 30660 800 30684 856
rect 31140 800 31164 856
rect 31524 800 31548 856
rect 32004 800 32028 856
rect 32388 800 32412 856
rect 32868 800 32892 856
rect 33348 800 33372 856
rect 33732 800 33756 856
rect 34212 800 34236 856
rect 34692 800 34716 856
rect 35076 800 35100 856
rect 35556 800 35580 856
rect 35940 800 35964 856
rect 36420 800 36444 856
rect 36900 800 36924 856
rect 37284 800 37308 856
rect 37764 800 37788 856
rect 38244 800 38268 856
rect 38628 800 38652 856
rect 39108 800 39132 856
rect 39588 800 39612 856
rect 39972 800 39996 856
rect 40452 800 40476 856
rect 40836 800 40860 856
rect 41316 800 41340 856
rect 41796 800 41820 856
rect 42180 800 42204 856
rect 42660 800 42684 856
rect 43140 800 43164 856
rect 43524 800 43548 856
rect 44004 800 44028 856
rect 44388 800 44412 856
rect 44868 800 44892 856
rect 45348 800 45372 856
rect 45732 800 45756 856
rect 46212 800 46236 856
rect 46692 800 46716 856
rect 47076 800 47100 856
rect 47556 800 47580 856
rect 47940 800 47964 856
rect 48420 800 48444 856
rect 48900 800 48924 856
rect 49284 800 49308 856
rect 49764 800 49788 856
rect 50244 800 50268 856
rect 50628 800 50652 856
rect 51108 800 51132 856
rect 51588 800 51612 856
rect 51972 800 51996 856
rect 52452 800 52476 856
rect 52836 800 52860 856
rect 53316 800 53340 856
rect 53796 800 53820 856
rect 54180 800 54204 856
rect 54660 800 54684 856
rect 55140 800 55164 856
rect 55524 800 55548 856
rect 56004 800 56028 856
rect 56388 800 56412 856
rect 56868 800 56892 856
rect 57348 800 57372 856
rect 57732 800 57756 856
rect 58212 800 58236 856
rect 58692 800 58716 856
rect 59076 800 59100 856
rect 59556 800 59580 856
<< metal3 >>
rect 0 44858 800 44978
rect 59200 29910 60000 30030
rect 0 14962 800 15082
<< obsm3 >>
rect 800 45058 59200 57309
rect 880 44778 59200 45058
rect 800 30110 59200 44778
rect 800 29830 59120 30110
rect 800 15162 59200 29830
rect 880 14882 59200 15162
rect 800 2409 59200 14882
<< metal4 >>
rect 4256 2616 4576 57324
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 2616 19936 57324
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 2616 35296 57324
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 2616 50656 57324
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
=======
rect 106 1232 179846 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10230 119200 10286 120000
rect 11794 119200 11850 120000
rect 13358 119200 13414 120000
rect 14922 119200 14978 120000
rect 16486 119200 16542 120000
rect 18050 119200 18106 120000
rect 19706 119200 19762 120000
rect 21270 119200 21326 120000
rect 22834 119200 22890 120000
rect 24398 119200 24454 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 29182 119200 29238 120000
rect 30746 119200 30802 120000
rect 32310 119200 32366 120000
rect 33874 119200 33930 120000
rect 35438 119200 35494 120000
rect 37002 119200 37058 120000
rect 38658 119200 38714 120000
rect 40222 119200 40278 120000
rect 41786 119200 41842 120000
rect 43350 119200 43406 120000
rect 44914 119200 44970 120000
rect 46478 119200 46534 120000
rect 48134 119200 48190 120000
rect 49698 119200 49754 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54390 119200 54446 120000
rect 55954 119200 56010 120000
rect 57610 119200 57666 120000
rect 59174 119200 59230 120000
rect 60738 119200 60794 120000
rect 62302 119200 62358 120000
rect 63866 119200 63922 120000
rect 65430 119200 65486 120000
rect 67086 119200 67142 120000
rect 68650 119200 68706 120000
rect 70214 119200 70270 120000
rect 71778 119200 71834 120000
rect 73342 119200 73398 120000
rect 74906 119200 74962 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79690 119200 79746 120000
rect 81254 119200 81310 120000
rect 82818 119200 82874 120000
rect 84382 119200 84438 120000
rect 86038 119200 86094 120000
rect 87602 119200 87658 120000
rect 89166 119200 89222 120000
rect 90730 119200 90786 120000
rect 92294 119200 92350 120000
rect 93858 119200 93914 120000
rect 95514 119200 95570 120000
rect 97078 119200 97134 120000
rect 98642 119200 98698 120000
rect 100206 119200 100262 120000
rect 101770 119200 101826 120000
rect 103334 119200 103390 120000
rect 104990 119200 105046 120000
rect 106554 119200 106610 120000
rect 108118 119200 108174 120000
rect 109682 119200 109738 120000
rect 111246 119200 111302 120000
rect 112810 119200 112866 120000
rect 114466 119200 114522 120000
rect 116030 119200 116086 120000
rect 117594 119200 117650 120000
rect 119158 119200 119214 120000
rect 120722 119200 120778 120000
rect 122286 119200 122342 120000
rect 123942 119200 123998 120000
rect 125506 119200 125562 120000
rect 127070 119200 127126 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131762 119200 131818 120000
rect 133418 119200 133474 120000
rect 134982 119200 135038 120000
rect 136546 119200 136602 120000
rect 138110 119200 138166 120000
rect 139674 119200 139730 120000
rect 141238 119200 141294 120000
rect 142894 119200 142950 120000
rect 144458 119200 144514 120000
rect 146022 119200 146078 120000
rect 147586 119200 147642 120000
rect 149150 119200 149206 120000
rect 150714 119200 150770 120000
rect 152370 119200 152426 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 157062 119200 157118 120000
rect 158626 119200 158682 120000
rect 160190 119200 160246 120000
rect 161846 119200 161902 120000
rect 163410 119200 163466 120000
rect 164974 119200 165030 120000
rect 166538 119200 166594 120000
rect 168102 119200 168158 120000
rect 169666 119200 169722 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39854 0 39910 800
rect 40222 0 40278 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97170 0 97226 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100114 0 100170 800
rect 100482 0 100538 800
rect 100850 0 100906 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102690 0 102746 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141422 0 141478 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 145010 0 145066 800
rect 145378 0 145434 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146850 0 146906 800
rect 147218 0 147274 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149794 0 149850 800
rect 150162 0 150218 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151266 0 151322 800
rect 151634 0 151690 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160742 0 160798 800
rect 161110 0 161166 800
rect 161478 0 161534 800
rect 161846 0 161902 800
rect 162214 0 162270 800
rect 162582 0 162638 800
rect 162950 0 163006 800
rect 163318 0 163374 800
rect 163686 0 163742 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164790 0 164846 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165894 0 165950 800
rect 166262 0 166318 800
rect 166630 0 166686 800
rect 166998 0 167054 800
rect 167366 0 167422 800
rect 167734 0 167790 800
rect 168102 0 168158 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 112 119144 698 119218
rect 866 119144 2262 119218
rect 2430 119144 3826 119218
rect 3994 119144 5390 119218
rect 5558 119144 6954 119218
rect 7122 119144 8518 119218
rect 8686 119144 10174 119218
rect 10342 119144 11738 119218
rect 11906 119144 13302 119218
rect 13470 119144 14866 119218
rect 15034 119144 16430 119218
rect 16598 119144 17994 119218
rect 18162 119144 19650 119218
rect 19818 119144 21214 119218
rect 21382 119144 22778 119218
rect 22946 119144 24342 119218
rect 24510 119144 25906 119218
rect 26074 119144 27470 119218
rect 27638 119144 29126 119218
rect 29294 119144 30690 119218
rect 30858 119144 32254 119218
rect 32422 119144 33818 119218
rect 33986 119144 35382 119218
rect 35550 119144 36946 119218
rect 37114 119144 38602 119218
rect 38770 119144 40166 119218
rect 40334 119144 41730 119218
rect 41898 119144 43294 119218
rect 43462 119144 44858 119218
rect 45026 119144 46422 119218
rect 46590 119144 48078 119218
rect 48246 119144 49642 119218
rect 49810 119144 51206 119218
rect 51374 119144 52770 119218
rect 52938 119144 54334 119218
rect 54502 119144 55898 119218
rect 56066 119144 57554 119218
rect 57722 119144 59118 119218
rect 59286 119144 60682 119218
rect 60850 119144 62246 119218
rect 62414 119144 63810 119218
rect 63978 119144 65374 119218
rect 65542 119144 67030 119218
rect 67198 119144 68594 119218
rect 68762 119144 70158 119218
rect 70326 119144 71722 119218
rect 71890 119144 73286 119218
rect 73454 119144 74850 119218
rect 75018 119144 76506 119218
rect 76674 119144 78070 119218
rect 78238 119144 79634 119218
rect 79802 119144 81198 119218
rect 81366 119144 82762 119218
rect 82930 119144 84326 119218
rect 84494 119144 85982 119218
rect 86150 119144 87546 119218
rect 87714 119144 89110 119218
rect 89278 119144 90674 119218
rect 90842 119144 92238 119218
rect 92406 119144 93802 119218
rect 93970 119144 95458 119218
rect 95626 119144 97022 119218
rect 97190 119144 98586 119218
rect 98754 119144 100150 119218
rect 100318 119144 101714 119218
rect 101882 119144 103278 119218
rect 103446 119144 104934 119218
rect 105102 119144 106498 119218
rect 106666 119144 108062 119218
rect 108230 119144 109626 119218
rect 109794 119144 111190 119218
rect 111358 119144 112754 119218
rect 112922 119144 114410 119218
rect 114578 119144 115974 119218
rect 116142 119144 117538 119218
rect 117706 119144 119102 119218
rect 119270 119144 120666 119218
rect 120834 119144 122230 119218
rect 122398 119144 123886 119218
rect 124054 119144 125450 119218
rect 125618 119144 127014 119218
rect 127182 119144 128578 119218
rect 128746 119144 130142 119218
rect 130310 119144 131706 119218
rect 131874 119144 133362 119218
rect 133530 119144 134926 119218
rect 135094 119144 136490 119218
rect 136658 119144 138054 119218
rect 138222 119144 139618 119218
rect 139786 119144 141182 119218
rect 141350 119144 142838 119218
rect 143006 119144 144402 119218
rect 144570 119144 145966 119218
rect 146134 119144 147530 119218
rect 147698 119144 149094 119218
rect 149262 119144 150658 119218
rect 150826 119144 152314 119218
rect 152482 119144 153878 119218
rect 154046 119144 155442 119218
rect 155610 119144 157006 119218
rect 157174 119144 158570 119218
rect 158738 119144 160134 119218
rect 160302 119144 161790 119218
rect 161958 119144 163354 119218
rect 163522 119144 164918 119218
rect 165086 119144 166482 119218
rect 166650 119144 168046 119218
rect 168214 119144 169610 119218
rect 169778 119144 171266 119218
rect 171434 119144 172830 119218
rect 172998 119144 174394 119218
rect 174562 119144 175958 119218
rect 176126 119144 177522 119218
rect 177690 119144 179086 119218
rect 179254 119144 179840 119218
rect 112 856 179840 119144
rect 222 734 330 856
rect 498 734 698 856
rect 866 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7322 856
rect 7490 734 7690 856
rect 7858 734 8058 856
rect 8226 734 8426 856
rect 8594 734 8794 856
rect 8962 734 9162 856
rect 9330 734 9530 856
rect 9698 734 9898 856
rect 10066 734 10266 856
rect 10434 734 10634 856
rect 10802 734 11002 856
rect 11170 734 11370 856
rect 11538 734 11738 856
rect 11906 734 12014 856
rect 12182 734 12382 856
rect 12550 734 12750 856
rect 12918 734 13118 856
rect 13286 734 13486 856
rect 13654 734 13854 856
rect 14022 734 14222 856
rect 14390 734 14590 856
rect 14758 734 14958 856
rect 15126 734 15326 856
rect 15494 734 15694 856
rect 15862 734 16062 856
rect 16230 734 16430 856
rect 16598 734 16798 856
rect 16966 734 17166 856
rect 17334 734 17534 856
rect 17702 734 17902 856
rect 18070 734 18270 856
rect 18438 734 18638 856
rect 18806 734 19006 856
rect 19174 734 19374 856
rect 19542 734 19742 856
rect 19910 734 20110 856
rect 20278 734 20478 856
rect 20646 734 20846 856
rect 21014 734 21214 856
rect 21382 734 21582 856
rect 21750 734 21950 856
rect 22118 734 22318 856
rect 22486 734 22686 856
rect 22854 734 23054 856
rect 23222 734 23422 856
rect 23590 734 23790 856
rect 23958 734 24066 856
rect 24234 734 24434 856
rect 24602 734 24802 856
rect 24970 734 25170 856
rect 25338 734 25538 856
rect 25706 734 25906 856
rect 26074 734 26274 856
rect 26442 734 26642 856
rect 26810 734 27010 856
rect 27178 734 27378 856
rect 27546 734 27746 856
rect 27914 734 28114 856
rect 28282 734 28482 856
rect 28650 734 28850 856
rect 29018 734 29218 856
rect 29386 734 29586 856
rect 29754 734 29954 856
rect 30122 734 30322 856
rect 30490 734 30690 856
rect 30858 734 31058 856
rect 31226 734 31426 856
rect 31594 734 31794 856
rect 31962 734 32162 856
rect 32330 734 32530 856
rect 32698 734 32898 856
rect 33066 734 33266 856
rect 33434 734 33634 856
rect 33802 734 34002 856
rect 34170 734 34370 856
rect 34538 734 34738 856
rect 34906 734 35106 856
rect 35274 734 35474 856
rect 35642 734 35842 856
rect 36010 734 36118 856
rect 36286 734 36486 856
rect 36654 734 36854 856
rect 37022 734 37222 856
rect 37390 734 37590 856
rect 37758 734 37958 856
rect 38126 734 38326 856
rect 38494 734 38694 856
rect 38862 734 39062 856
rect 39230 734 39430 856
rect 39598 734 39798 856
rect 39966 734 40166 856
rect 40334 734 40534 856
rect 40702 734 40902 856
rect 41070 734 41270 856
rect 41438 734 41638 856
rect 41806 734 42006 856
rect 42174 734 42374 856
rect 42542 734 42742 856
rect 42910 734 43110 856
rect 43278 734 43478 856
rect 43646 734 43846 856
rect 44014 734 44214 856
rect 44382 734 44582 856
rect 44750 734 44950 856
rect 45118 734 45318 856
rect 45486 734 45686 856
rect 45854 734 46054 856
rect 46222 734 46422 856
rect 46590 734 46790 856
rect 46958 734 47158 856
rect 47326 734 47526 856
rect 47694 734 47894 856
rect 48062 734 48170 856
rect 48338 734 48538 856
rect 48706 734 48906 856
rect 49074 734 49274 856
rect 49442 734 49642 856
rect 49810 734 50010 856
rect 50178 734 50378 856
rect 50546 734 50746 856
rect 50914 734 51114 856
rect 51282 734 51482 856
rect 51650 734 51850 856
rect 52018 734 52218 856
rect 52386 734 52586 856
rect 52754 734 52954 856
rect 53122 734 53322 856
rect 53490 734 53690 856
rect 53858 734 54058 856
rect 54226 734 54426 856
rect 54594 734 54794 856
rect 54962 734 55162 856
rect 55330 734 55530 856
rect 55698 734 55898 856
rect 56066 734 56266 856
rect 56434 734 56634 856
rect 56802 734 57002 856
rect 57170 734 57370 856
rect 57538 734 57738 856
rect 57906 734 58106 856
rect 58274 734 58474 856
rect 58642 734 58842 856
rect 59010 734 59210 856
rect 59378 734 59578 856
rect 59746 734 59946 856
rect 60114 734 60222 856
rect 60390 734 60590 856
rect 60758 734 60958 856
rect 61126 734 61326 856
rect 61494 734 61694 856
rect 61862 734 62062 856
rect 62230 734 62430 856
rect 62598 734 62798 856
rect 62966 734 63166 856
rect 63334 734 63534 856
rect 63702 734 63902 856
rect 64070 734 64270 856
rect 64438 734 64638 856
rect 64806 734 65006 856
rect 65174 734 65374 856
rect 65542 734 65742 856
rect 65910 734 66110 856
rect 66278 734 66478 856
rect 66646 734 66846 856
rect 67014 734 67214 856
rect 67382 734 67582 856
rect 67750 734 67950 856
rect 68118 734 68318 856
rect 68486 734 68686 856
rect 68854 734 69054 856
rect 69222 734 69422 856
rect 69590 734 69790 856
rect 69958 734 70158 856
rect 70326 734 70526 856
rect 70694 734 70894 856
rect 71062 734 71262 856
rect 71430 734 71630 856
rect 71798 734 71998 856
rect 72166 734 72274 856
rect 72442 734 72642 856
rect 72810 734 73010 856
rect 73178 734 73378 856
rect 73546 734 73746 856
rect 73914 734 74114 856
rect 74282 734 74482 856
rect 74650 734 74850 856
rect 75018 734 75218 856
rect 75386 734 75586 856
rect 75754 734 75954 856
rect 76122 734 76322 856
rect 76490 734 76690 856
rect 76858 734 77058 856
rect 77226 734 77426 856
rect 77594 734 77794 856
rect 77962 734 78162 856
rect 78330 734 78530 856
rect 78698 734 78898 856
rect 79066 734 79266 856
rect 79434 734 79634 856
rect 79802 734 80002 856
rect 80170 734 80370 856
rect 80538 734 80738 856
rect 80906 734 81106 856
rect 81274 734 81474 856
rect 81642 734 81842 856
rect 82010 734 82210 856
rect 82378 734 82578 856
rect 82746 734 82946 856
rect 83114 734 83314 856
rect 83482 734 83682 856
rect 83850 734 84050 856
rect 84218 734 84326 856
rect 84494 734 84694 856
rect 84862 734 85062 856
rect 85230 734 85430 856
rect 85598 734 85798 856
rect 85966 734 86166 856
rect 86334 734 86534 856
rect 86702 734 86902 856
rect 87070 734 87270 856
rect 87438 734 87638 856
rect 87806 734 88006 856
rect 88174 734 88374 856
rect 88542 734 88742 856
rect 88910 734 89110 856
rect 89278 734 89478 856
rect 89646 734 89846 856
rect 90014 734 90214 856
rect 90382 734 90582 856
rect 90750 734 90950 856
rect 91118 734 91318 856
rect 91486 734 91686 856
rect 91854 734 92054 856
rect 92222 734 92422 856
rect 92590 734 92790 856
rect 92958 734 93158 856
rect 93326 734 93526 856
rect 93694 734 93894 856
rect 94062 734 94262 856
rect 94430 734 94630 856
rect 94798 734 94998 856
rect 95166 734 95366 856
rect 95534 734 95734 856
rect 95902 734 96010 856
rect 96178 734 96378 856
rect 96546 734 96746 856
rect 96914 734 97114 856
rect 97282 734 97482 856
rect 97650 734 97850 856
rect 98018 734 98218 856
rect 98386 734 98586 856
rect 98754 734 98954 856
rect 99122 734 99322 856
rect 99490 734 99690 856
rect 99858 734 100058 856
rect 100226 734 100426 856
rect 100594 734 100794 856
rect 100962 734 101162 856
rect 101330 734 101530 856
rect 101698 734 101898 856
rect 102066 734 102266 856
rect 102434 734 102634 856
rect 102802 734 103002 856
rect 103170 734 103370 856
rect 103538 734 103738 856
rect 103906 734 104106 856
rect 104274 734 104474 856
rect 104642 734 104842 856
rect 105010 734 105210 856
rect 105378 734 105578 856
rect 105746 734 105946 856
rect 106114 734 106314 856
rect 106482 734 106682 856
rect 106850 734 107050 856
rect 107218 734 107418 856
rect 107586 734 107786 856
rect 107954 734 108062 856
rect 108230 734 108430 856
rect 108598 734 108798 856
rect 108966 734 109166 856
rect 109334 734 109534 856
rect 109702 734 109902 856
rect 110070 734 110270 856
rect 110438 734 110638 856
rect 110806 734 111006 856
rect 111174 734 111374 856
rect 111542 734 111742 856
rect 111910 734 112110 856
rect 112278 734 112478 856
rect 112646 734 112846 856
rect 113014 734 113214 856
rect 113382 734 113582 856
rect 113750 734 113950 856
rect 114118 734 114318 856
rect 114486 734 114686 856
rect 114854 734 115054 856
rect 115222 734 115422 856
rect 115590 734 115790 856
rect 115958 734 116158 856
rect 116326 734 116526 856
rect 116694 734 116894 856
rect 117062 734 117262 856
rect 117430 734 117630 856
rect 117798 734 117998 856
rect 118166 734 118366 856
rect 118534 734 118734 856
rect 118902 734 119102 856
rect 119270 734 119470 856
rect 119638 734 119838 856
rect 120006 734 120114 856
rect 120282 734 120482 856
rect 120650 734 120850 856
rect 121018 734 121218 856
rect 121386 734 121586 856
rect 121754 734 121954 856
rect 122122 734 122322 856
rect 122490 734 122690 856
rect 122858 734 123058 856
rect 123226 734 123426 856
rect 123594 734 123794 856
rect 123962 734 124162 856
rect 124330 734 124530 856
rect 124698 734 124898 856
rect 125066 734 125266 856
rect 125434 734 125634 856
rect 125802 734 126002 856
rect 126170 734 126370 856
rect 126538 734 126738 856
rect 126906 734 127106 856
rect 127274 734 127474 856
rect 127642 734 127842 856
rect 128010 734 128210 856
rect 128378 734 128578 856
rect 128746 734 128946 856
rect 129114 734 129314 856
rect 129482 734 129682 856
rect 129850 734 130050 856
rect 130218 734 130418 856
rect 130586 734 130786 856
rect 130954 734 131154 856
rect 131322 734 131522 856
rect 131690 734 131890 856
rect 132058 734 132166 856
rect 132334 734 132534 856
rect 132702 734 132902 856
rect 133070 734 133270 856
rect 133438 734 133638 856
rect 133806 734 134006 856
rect 134174 734 134374 856
rect 134542 734 134742 856
rect 134910 734 135110 856
rect 135278 734 135478 856
rect 135646 734 135846 856
rect 136014 734 136214 856
rect 136382 734 136582 856
rect 136750 734 136950 856
rect 137118 734 137318 856
rect 137486 734 137686 856
rect 137854 734 138054 856
rect 138222 734 138422 856
rect 138590 734 138790 856
rect 138958 734 139158 856
rect 139326 734 139526 856
rect 139694 734 139894 856
rect 140062 734 140262 856
rect 140430 734 140630 856
rect 140798 734 140998 856
rect 141166 734 141366 856
rect 141534 734 141734 856
rect 141902 734 142102 856
rect 142270 734 142470 856
rect 142638 734 142838 856
rect 143006 734 143206 856
rect 143374 734 143574 856
rect 143742 734 143942 856
rect 144110 734 144218 856
rect 144386 734 144586 856
rect 144754 734 144954 856
rect 145122 734 145322 856
rect 145490 734 145690 856
rect 145858 734 146058 856
rect 146226 734 146426 856
rect 146594 734 146794 856
rect 146962 734 147162 856
rect 147330 734 147530 856
rect 147698 734 147898 856
rect 148066 734 148266 856
rect 148434 734 148634 856
rect 148802 734 149002 856
rect 149170 734 149370 856
rect 149538 734 149738 856
rect 149906 734 150106 856
rect 150274 734 150474 856
rect 150642 734 150842 856
rect 151010 734 151210 856
rect 151378 734 151578 856
rect 151746 734 151946 856
rect 152114 734 152314 856
rect 152482 734 152682 856
rect 152850 734 153050 856
rect 153218 734 153418 856
rect 153586 734 153786 856
rect 153954 734 154154 856
rect 154322 734 154522 856
rect 154690 734 154890 856
rect 155058 734 155258 856
rect 155426 734 155626 856
rect 155794 734 155994 856
rect 156162 734 156270 856
rect 156438 734 156638 856
rect 156806 734 157006 856
rect 157174 734 157374 856
rect 157542 734 157742 856
rect 157910 734 158110 856
rect 158278 734 158478 856
rect 158646 734 158846 856
rect 159014 734 159214 856
rect 159382 734 159582 856
rect 159750 734 159950 856
rect 160118 734 160318 856
rect 160486 734 160686 856
rect 160854 734 161054 856
rect 161222 734 161422 856
rect 161590 734 161790 856
rect 161958 734 162158 856
rect 162326 734 162526 856
rect 162694 734 162894 856
rect 163062 734 163262 856
rect 163430 734 163630 856
rect 163798 734 163998 856
rect 164166 734 164366 856
rect 164534 734 164734 856
rect 164902 734 165102 856
rect 165270 734 165470 856
rect 165638 734 165838 856
rect 166006 734 166206 856
rect 166374 734 166574 856
rect 166742 734 166942 856
rect 167110 734 167310 856
rect 167478 734 167678 856
rect 167846 734 168046 856
rect 168214 734 168322 856
rect 168490 734 168690 856
rect 168858 734 169058 856
rect 169226 734 169426 856
rect 169594 734 169794 856
rect 169962 734 170162 856
rect 170330 734 170530 856
rect 170698 734 170898 856
rect 171066 734 171266 856
rect 171434 734 171634 856
rect 171802 734 172002 856
rect 172170 734 172370 856
rect 172538 734 172738 856
rect 172906 734 173106 856
rect 173274 734 173474 856
rect 173642 734 173842 856
rect 174010 734 174210 856
rect 174378 734 174578 856
rect 174746 734 174946 856
rect 175114 734 175314 856
rect 175482 734 175682 856
rect 175850 734 176050 856
rect 176218 734 176418 856
rect 176586 734 176786 856
rect 176954 734 177154 856
rect 177322 734 177522 856
rect 177690 734 177890 856
rect 178058 734 178258 856
rect 178426 734 178626 856
rect 178794 734 178994 856
rect 179162 734 179362 856
rect 179530 734 179730 856
<< obsm3 >>
rect 1669 1803 173488 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
<< obsm4 >>
rect 34928 1803 173488 117552
>>>>>>> c5da9e9885e361d05dee2aa6303a69fc26423c8e
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 114 nsew signal output
<<<<<<< HEAD
rlabel metal3 s 0 14962 800 15082 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 59200 29910 60000 30030 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 44858 800 44978 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 13172 0 13228 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 610 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 611 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 612 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 613 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 614 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 615 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 616 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 617 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 618 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 619 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 620 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 621 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 622 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 623 nsew ground bidirectional
=======
rlabel metal2 s 179050 0 179106 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 158534 0 158590 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 160742 0 160798 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 161846 0 161902 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 164054 0 164110 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 165158 0 165214 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 126794 0 126850 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 609 nsew signal input
>>>>>>> c5da9e9885e361d05dee2aa6303a69fc26423c8e
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
<<<<<<< HEAD
string GDS_END 2182180
string GDS_START 251226
=======
string GDS_END 8095954
string GDS_START 360410
>>>>>>> c5da9e9885e361d05dee2aa6303a69fc26423c8e
<< end >>

