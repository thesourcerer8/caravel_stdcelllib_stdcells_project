magic
tech sky130A
timestamp 1624067522
<< nwell >>
rect 0 179 576 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
<< ndiff >>
rect 226 67 255 73
rect 226 66 232 67
rect 58 49 137 66
rect 58 32 64 49
rect 81 32 137 49
rect 58 24 137 32
rect 152 50 232 66
rect 249 66 255 67
rect 466 67 495 73
rect 466 66 472 67
rect 249 50 281 66
rect 152 24 281 50
rect 296 49 425 66
rect 296 32 328 49
rect 345 32 425 49
rect 296 24 425 32
rect 440 50 472 66
rect 489 66 495 67
rect 489 50 519 66
rect 440 24 519 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 88 243
rect 105 226 137 243
rect 58 225 137 226
rect 152 225 281 309
rect 296 301 425 309
rect 296 284 328 301
rect 345 284 425 301
rect 296 225 425 284
rect 440 243 519 309
rect 440 226 472 243
rect 489 226 519 243
rect 440 225 519 226
rect 82 220 111 225
rect 466 220 495 225
<< ndiffc >>
rect 64 32 81 49
rect 232 50 249 67
rect 328 32 345 49
rect 472 50 489 67
<< pdiffc >>
rect 88 226 105 243
rect 328 284 345 301
rect 472 226 489 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
<< locali >>
rect 320 301 353 309
rect 320 284 328 301
rect 345 284 353 301
rect 320 276 353 284
rect 80 243 113 251
rect 80 226 88 243
rect 105 226 113 243
rect 464 243 497 251
rect 464 226 472 243
rect 489 226 497 243
rect 80 218 111 226
rect 466 218 497 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 136 116 153 131
rect 280 116 297 176
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 272 108 305 116
rect 272 92 280 108
rect 128 83 161 91
rect 274 91 280 92
rect 297 91 305 108
rect 274 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 224 67 257 75
rect 56 49 89 57
rect 56 32 64 49
rect 81 32 89 49
rect 224 50 232 67
rect 249 50 257 67
rect 466 67 497 75
rect 466 66 472 67
rect 224 42 257 50
rect 320 49 353 57
rect 56 24 89 32
rect 320 32 328 49
rect 345 32 353 49
rect 464 50 472 66
rect 489 50 497 67
rect 464 42 497 50
rect 320 24 353 32
<< viali >>
rect 328 284 345 301
rect 88 226 105 243
rect 472 226 489 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 131 153 148
rect 424 91 441 108
rect 64 32 81 49
rect 232 50 249 67
rect 328 32 345 49
rect 472 50 489 67
<< metal1 >>
rect 0 309 576 357
rect 322 301 351 309
rect 322 284 328 301
rect 345 284 351 301
rect 322 278 351 284
rect 82 243 111 249
rect 82 226 88 243
rect 105 226 111 243
rect 82 220 111 226
rect 466 243 495 249
rect 466 226 472 243
rect 489 226 495 243
rect 466 220 495 226
rect 89 106 103 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 137 154 151 178
rect 130 148 159 154
rect 130 131 136 148
rect 153 131 159 148
rect 130 125 159 131
rect 425 114 439 178
rect 418 108 447 114
rect 418 106 424 108
rect 89 92 424 106
rect 233 73 247 92
rect 418 91 424 92
rect 441 91 447 108
rect 418 85 447 91
rect 473 73 487 220
rect 226 67 255 73
rect 58 49 87 55
rect 58 32 64 49
rect 81 32 87 49
rect 226 50 232 67
rect 249 50 255 67
rect 466 67 495 73
rect 226 44 255 50
rect 322 49 351 55
rect 58 24 87 32
rect 322 32 328 49
rect 345 32 351 49
rect 466 50 472 67
rect 489 50 495 67
rect 466 44 495 50
rect 322 24 351 32
rect 0 -24 576 24
<< labels >>
rlabel metal1 0 309 576 357 0 VDD
port 1 se
rlabel metal1 0 -24 576 24 0 GND
port 2 se
rlabel metal1 466 44 495 73 0 Y
port 3 se
rlabel metal1 473 73 487 220 0 Y
port 4 se
rlabel metal1 466 220 495 249 0 Y
port 5 se
rlabel metal1 130 125 159 154 0 A
port 6 se
rlabel metal1 137 154 151 178 0 A
port 7 se
rlabel metal1 130 178 159 207 0 A
port 8 se
rlabel metal1 274 178 303 207 0 B
port 9 se
<< properties >>
string FIXED_BBOX 0 0 576 333
<< end >>
