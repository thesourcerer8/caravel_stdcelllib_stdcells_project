VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LOFTY
  CLASS CORE ;
  FOREIGN LOFTY ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.600 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 21.600 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 21.600 0.240 ;
    END
  END gnd
  PIN Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.020 2.290 2.550 2.580 ;
        RECT 2.090 0.690 2.230 2.290 ;
        RECT 2.020 0.400 2.310 0.690 ;
    END
  END Q
  PIN ASEL_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.750 5.910 2.040 ;
        RECT 5.690 1.090 5.830 1.750 ;
        RECT 5.620 0.800 5.910 1.090 ;
    END
  END ASEL_P
  PIN USEXOR_N
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 15.700 0.750 15.990 0.820 ;
        RECT 20.020 0.750 20.310 0.820 ;
        RECT 15.700 0.610 20.310 0.750 ;
        RECT 15.700 0.530 15.990 0.610 ;
        RECT 20.020 0.530 20.310 0.610 ;
    END
  END USEXOR_N
  PIN USEMUX_N
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.890 2.230 1.750 2.370 ;
        RECT 0.890 0.690 1.030 2.230 ;
        RECT 1.540 2.170 1.750 2.230 ;
        RECT 1.540 2.040 1.830 2.170 ;
        RECT 1.300 1.880 1.830 2.040 ;
        RECT 1.300 1.750 1.590 1.880 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
        RECT 0.820 0.400 1.110 0.690 ;
    END
  END USEMUX_N
  PIN USEXOR_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 17.140 1.750 17.430 2.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.500 1.750 8.790 2.040 ;
    END
  END USEXOR_P
  PIN ASEL_N
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.060 1.340 7.350 1.630 ;
        RECT 7.130 1.090 7.270 1.340 ;
        RECT 7.060 0.800 7.350 1.090 ;
    END
  END ASEL_N
  PIN BSEL_N
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 18.580 1.340 18.870 2.040 ;
    END
  END BSEL_N
  PIN BSEL_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 14.260 1.340 14.550 1.630 ;
    END
  END BSEL_P
  PIN MUXSEL_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.540 2.500 7.830 2.580 ;
        RECT 7.540 2.360 9.190 2.500 ;
        RECT 7.540 2.290 7.830 2.360 ;
        RECT 9.050 2.230 9.190 2.360 ;
        RECT 10.420 2.230 10.710 2.310 ;
        RECT 11.620 2.230 11.910 2.310 ;
        RECT 9.050 2.090 10.710 2.230 ;
        RECT 10.420 2.040 10.710 2.090 ;
        RECT 10.970 2.090 11.910 2.230 ;
        RECT 10.970 2.040 11.110 2.090 ;
        RECT 10.420 2.020 11.110 2.040 ;
        RECT 11.620 2.040 11.910 2.090 ;
        RECT 11.620 2.020 12.150 2.040 ;
        RECT 10.660 1.820 11.110 2.020 ;
        RECT 10.660 1.750 10.950 1.820 ;
        RECT 11.860 1.750 12.150 2.020 ;
    END
  END MUXSEL_P
  PIN USEMUX_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.570 2.230 3.430 2.370 ;
        RECT 2.570 2.170 2.790 2.230 ;
        RECT 2.500 2.040 2.790 2.170 ;
        RECT 2.500 1.880 3.030 2.040 ;
        RECT 2.740 1.750 3.030 1.880 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 3.290 1.500 3.430 2.230 ;
        RECT 3.220 1.210 3.510 1.500 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END USEMUX_P
END LOFTY
END LIBRARY

