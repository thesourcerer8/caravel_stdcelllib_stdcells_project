magic
tech sky130A
timestamp 1624190759
<< nwell >>
rect 0 179 1008 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
rect 857 24 872 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
rect 857 225 872 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 514 67 543 73
rect 514 66 520 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 51 281 66
rect 152 34 184 51
rect 201 34 281 51
rect 152 24 281 34
rect 296 24 425 66
rect 440 50 520 66
rect 537 66 543 67
rect 898 67 927 73
rect 898 66 904 67
rect 537 50 569 66
rect 440 24 569 50
rect 584 24 713 66
rect 728 51 857 66
rect 728 34 760 51
rect 777 34 857 51
rect 728 24 857 34
rect 872 50 904 66
rect 921 66 927 67
rect 921 50 951 66
rect 872 24 951 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 225 425 309
rect 440 243 569 309
rect 440 226 520 243
rect 537 226 569 243
rect 440 225 569 226
rect 584 225 713 309
rect 728 299 857 309
rect 728 282 760 299
rect 777 282 857 299
rect 728 225 857 282
rect 872 243 951 309
rect 872 226 904 243
rect 921 226 951 243
rect 872 225 951 226
rect 58 220 87 225
rect 514 220 543 225
rect 898 220 927 225
<< ndiffc >>
rect 64 50 81 67
rect 184 34 201 51
rect 520 50 537 67
rect 760 34 777 51
rect 904 50 921 67
<< pdiffc >>
rect 64 226 81 243
rect 184 282 201 299
rect 520 226 537 243
rect 760 282 777 299
rect 904 226 921 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 713 309 728 322
rect 857 309 872 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 713 209 728 225
rect 857 209 872 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 848 201 881 209
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 713 66 728 83
rect 857 66 872 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
rect 857 11 872 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 856 184 873 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
rect 856 91 873 108
<< locali >>
rect 760 307 777 325
rect 176 299 209 307
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 752 299 785 307
rect 752 282 760 299
rect 777 282 785 299
rect 752 274 785 282
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 512 243 545 251
rect 512 226 520 243
rect 537 226 545 243
rect 896 243 929 251
rect 896 226 904 243
rect 921 226 929 243
rect 512 218 543 226
rect 898 218 929 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 416 201 449 209
rect 272 184 280 201
rect 297 184 305 201
rect 345 184 424 201
rect 441 184 449 201
rect 272 176 305 184
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 848 201 881 209
rect 848 184 856 201
rect 873 184 881 201
rect 848 176 881 184
rect 280 116 297 176
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 560 108 593 116
rect 560 92 568 108
rect 416 83 449 91
rect 562 91 568 92
rect 585 91 593 108
rect 562 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 848 108 881 116
rect 848 91 856 108
rect 873 91 881 108
rect 848 83 881 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 512 67 545 75
rect 56 42 89 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 512 50 520 67
rect 537 50 545 67
rect 898 67 929 75
rect 898 66 904 67
rect 512 42 545 50
rect 752 51 785 59
rect 176 26 209 34
rect 752 34 760 51
rect 777 34 785 51
rect 896 50 904 66
rect 921 50 929 67
rect 896 42 929 50
rect 752 26 785 34
rect 184 9 201 26
rect 760 9 777 26
<< viali >>
rect 760 325 777 342
rect 184 282 201 299
rect 64 226 81 243
rect 520 226 537 243
rect 904 226 921 243
rect 136 184 153 201
rect 280 184 297 201
rect 328 184 345 201
rect 568 184 585 201
rect 712 184 729 201
rect 856 184 873 201
rect 136 91 153 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
rect 856 91 873 108
rect 64 50 81 67
rect 520 50 537 67
rect 904 50 921 67
rect 184 -9 201 9
rect 760 -9 777 9
<< metal1 >>
rect 0 342 1008 357
rect 0 325 760 342
rect 777 325 1008 342
rect 0 309 1008 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 281 268 871 282
rect 58 243 87 249
rect 58 226 64 243
rect 81 241 87 243
rect 81 227 199 241
rect 81 226 87 227
rect 58 220 87 226
rect 65 73 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 137 114 151 178
rect 185 160 199 227
rect 281 207 295 268
rect 514 243 543 249
rect 514 226 520 243
rect 537 241 543 243
rect 537 227 631 241
rect 537 226 543 227
rect 514 220 543 226
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 322 201 351 207
rect 322 184 328 201
rect 345 184 351 201
rect 562 201 591 207
rect 562 200 568 201
rect 322 178 351 184
rect 425 186 568 200
rect 329 160 343 178
rect 185 146 343 160
rect 425 114 439 186
rect 562 184 568 186
rect 585 184 591 201
rect 562 178 591 184
rect 130 108 159 114
rect 130 91 136 108
rect 153 106 159 108
rect 418 108 447 114
rect 418 106 424 108
rect 153 92 424 106
rect 153 91 159 92
rect 130 85 159 91
rect 418 91 424 92
rect 441 91 447 108
rect 562 108 591 114
rect 562 106 568 108
rect 418 85 447 91
rect 473 92 568 106
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 473 66 487 92
rect 562 91 568 92
rect 585 91 591 108
rect 562 85 591 91
rect 81 52 487 66
rect 514 67 543 73
rect 81 50 87 52
rect 58 44 87 50
rect 514 50 520 67
rect 537 66 543 67
rect 617 66 631 227
rect 857 207 871 268
rect 898 243 927 249
rect 898 226 904 243
rect 921 226 927 243
rect 898 220 927 226
rect 706 201 735 207
rect 706 184 712 201
rect 729 184 735 201
rect 706 178 735 184
rect 850 201 879 207
rect 850 184 856 201
rect 873 184 879 201
rect 850 178 879 184
rect 713 114 727 178
rect 857 114 871 178
rect 706 108 735 114
rect 706 91 712 108
rect 729 91 735 108
rect 706 85 735 91
rect 850 108 879 114
rect 850 91 856 108
rect 873 91 879 108
rect 850 85 879 91
rect 537 52 631 66
rect 713 66 727 85
rect 905 73 919 220
rect 898 67 927 73
rect 898 66 904 67
rect 713 52 904 66
rect 537 50 543 52
rect 514 44 543 50
rect 898 50 904 52
rect 921 50 927 67
rect 898 44 927 50
rect 0 9 1008 24
rect 0 -9 184 9
rect 201 -9 760 9
rect 777 -9 1008 9
rect 0 -24 1008 -9
<< labels >>
rlabel metal1 0 309 1008 357 0 VDD
port 1 se
rlabel metal1 0 -24 1008 24 0 GND
port 2 se
rlabel metal1 514 44 543 52 0 Y
port 3 se
rlabel metal1 514 52 631 66 0 Y
port 4 se
rlabel metal1 514 66 543 73 0 Y
port 5 se
rlabel metal1 514 220 543 227 0 Y
port 6 se
rlabel metal1 617 66 631 227 0 Y
port 7 se
rlabel metal1 514 227 631 241 0 Y
port 8 se
rlabel metal1 514 241 543 249 0 Y
port 9 se
rlabel metal1 130 85 159 92 0 A
port 10 se
rlabel metal1 418 85 447 92 0 A
port 11 se
rlabel metal1 130 92 447 106 0 A
port 12 se
rlabel metal1 130 106 159 114 0 A
port 13 se
rlabel metal1 418 106 447 114 0 A
port 14 se
rlabel metal1 137 114 151 178 0 A
port 15 se
rlabel metal1 425 114 439 186 0 A
port 16 se
rlabel metal1 562 178 591 186 0 A
port 17 se
rlabel metal1 425 186 591 200 0 A
port 18 se
rlabel metal1 130 178 159 207 0 A
port 19 se
rlabel metal1 562 200 591 207 0 A
port 20 se
rlabel metal1 850 85 879 114 0 B
port 21 se
rlabel metal1 857 114 871 178 0 B
port 22 se
rlabel metal1 274 178 303 207 0 B
port 23 se
rlabel metal1 850 178 879 207 0 B
port 24 se
rlabel metal1 281 207 295 268 0 B
port 25 se
rlabel metal1 857 207 871 268 0 B
port 26 se
rlabel metal1 281 268 871 282 0 B
port 27 se
<< properties >>
string FIXED_BBOX 0 0 1008 333
<< end >>
