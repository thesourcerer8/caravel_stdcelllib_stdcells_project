VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ASYNC2
  CLASS CORE ;
  FOREIGN ASYNC2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 2.735 0.845 3.025 1.135 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA 0.189000 ;
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 6.095 2.410 6.385 2.485 ;
        RECT 4.250 2.270 6.385 2.410 ;
        RECT 4.250 2.070 4.390 2.270 ;
        RECT 6.095 2.195 6.385 2.270 ;
        RECT 4.175 1.780 4.465 2.070 ;
        RECT 6.170 0.730 6.310 2.195 ;
        RECT 6.095 0.440 6.385 0.730 ;
    END
  END C
  PIN CN
    ANTENNAGATEAREA 0.189000 ;
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 3.215 2.195 3.505 2.485 ;
        RECT 3.290 1.060 3.430 2.195 ;
        RECT 5.615 1.780 5.905 2.070 ;
        RECT 5.690 1.135 5.830 1.780 ;
        RECT 5.615 1.060 5.905 1.135 ;
        RECT 3.290 0.920 5.905 1.060 ;
        RECT 3.290 0.730 3.430 0.920 ;
        RECT 5.615 0.845 5.905 0.920 ;
        RECT 3.215 0.440 3.505 0.730 ;
    END
  END CN
  PIN VGND
    ANTENNADIFFAREA 0.914200 ;
    PORT
      LAYER met1 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 0.650 0.240 0.790 0.440 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
        RECT 0.575 2.735 0.865 3.090 ;
        RECT 4.655 2.735 4.945 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 0.663600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 7.200 3.415 ;
        RECT 0.155 3.215 7.045 3.245 ;
        RECT 0.155 3.090 4.465 3.215 ;
        RECT 5.135 3.090 7.045 3.215 ;
        RECT 0.555 2.715 0.885 3.090 ;
      LAYER mcon ;
        RECT 4.715 3.245 4.885 3.415 ;
        RECT 0.635 2.795 0.805 2.965 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 7.200 3.330 ;
      LAYER li1 ;
        RECT 4.635 2.715 4.965 3.045 ;
        RECT 3.195 2.260 3.525 2.505 ;
        RECT 6.075 2.260 6.405 2.505 ;
        RECT 3.215 2.175 3.525 2.260 ;
        RECT 6.095 2.175 6.405 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 4.235 1.155 4.405 1.760 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 2.715 0.825 3.025 0.920 ;
        RECT 4.155 0.825 4.485 1.155 ;
        RECT 5.595 0.920 5.925 1.155 ;
        RECT 5.595 0.825 5.905 0.920 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 3.195 0.420 3.525 0.750 ;
        RECT 4.655 0.655 4.965 0.750 ;
        RECT 4.635 0.420 4.965 0.655 ;
        RECT 6.075 0.420 6.405 0.750 ;
        RECT 4.715 0.240 4.885 0.420 ;
        RECT 0.155 0.085 7.045 0.240 ;
        RECT 0.000 -0.085 7.200 0.085 ;
      LAYER mcon ;
        RECT 4.715 2.795 4.885 2.965 ;
        RECT 3.275 2.255 3.445 2.425 ;
        RECT 6.155 2.255 6.325 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 5.675 1.840 5.845 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 6.155 0.500 6.325 0.670 ;
        RECT 4.715 -0.085 4.885 0.085 ;
  END
END ASYNC2
END LIBRARY

