magic
tech sky130A
magscale 1 2
timestamp 1624893035
<< locali >>
rect 23935 52742 23969 52856
rect 22399 40828 22433 40942
rect 8479 26512 8801 26546
rect 8479 26472 8513 26512
rect 8383 26438 8513 26472
rect 8767 26472 8801 26512
rect 8383 26398 8417 26438
rect 30079 23438 30113 23552
rect 8191 22476 8225 22516
rect 8095 22442 8225 22476
rect 8095 22106 8129 22442
rect 7903 18480 7937 18520
rect 8191 18480 8225 18520
rect 7903 18446 8225 18480
rect 7039 8342 7073 8530
rect 7999 5530 8033 5644
rect 21631 5530 21665 5644
rect 26623 5530 26657 5644
rect 37951 5530 37985 5644
rect 7711 5160 7745 5200
rect 7903 5200 8225 5234
rect 7903 5160 7937 5200
rect 7711 5126 7937 5160
rect 8191 5160 8225 5200
rect 8479 5160 8513 5200
rect 8191 5126 8513 5160
rect 21151 2866 21185 3054
<< viali >>
rect 9919 57000 9953 57034
rect 14047 57000 14081 57034
rect 32575 57000 32609 57034
rect 1951 56926 1985 56960
rect 2815 56926 2849 56960
rect 5311 56926 5345 56960
rect 5791 56926 5825 56960
rect 7423 56926 7457 56960
rect 8095 56926 8129 56960
rect 11455 56926 11489 56960
rect 13183 56926 13217 56960
rect 15103 56926 15137 56960
rect 16351 56926 16385 56960
rect 18175 56926 18209 56960
rect 19519 56926 19553 56960
rect 21055 56926 21089 56960
rect 22015 56926 22049 56960
rect 24223 56926 24257 56960
rect 25951 56926 25985 56960
rect 27391 56926 27425 56960
rect 28639 56926 28673 56960
rect 30271 56926 30305 56960
rect 31711 56926 31745 56960
rect 34303 56926 34337 56960
rect 34879 56926 34913 56960
rect 38047 56926 38081 56960
rect 41983 56926 42017 56960
rect 44671 56926 44705 56960
rect 47551 56926 47585 56960
rect 53887 56926 53921 56960
rect 1759 56852 1793 56886
rect 2623 56852 2657 56886
rect 5119 56852 5153 56886
rect 7231 56852 7265 56886
rect 11263 56852 11297 56886
rect 12991 56852 13025 56886
rect 13951 56852 13985 56886
rect 16159 56852 16193 56886
rect 17983 56852 18017 56886
rect 19327 56852 19361 56886
rect 20863 56852 20897 56886
rect 24031 56852 24065 56886
rect 27199 56852 27233 56886
rect 30079 56852 30113 56886
rect 32671 56852 32705 56886
rect 34111 56852 34145 56886
rect 36991 56852 37025 56886
rect 40063 56852 40097 56886
rect 40543 56852 40577 56886
rect 40735 56852 40769 56886
rect 43231 56852 43265 56886
rect 46303 56852 46337 56886
rect 48991 56852 49025 56886
rect 51103 56852 51137 56886
rect 53119 56852 53153 56886
rect 55807 56852 55841 56886
rect 57055 56852 57089 56886
rect 9823 56704 9857 56738
rect 13663 56704 13697 56738
rect 36703 56704 36737 56738
rect 39775 56704 39809 56738
rect 40831 56704 40865 56738
rect 42943 56704 42977 56738
rect 46015 56704 46049 56738
rect 48703 56704 48737 56738
rect 50815 56704 50849 56738
rect 52831 56704 52865 56738
rect 55519 56704 55553 56738
rect 56767 56704 56801 56738
rect 1663 56482 1697 56516
rect 2431 56482 2465 56516
rect 3199 56482 3233 56516
rect 4447 56482 4481 56516
rect 5503 56482 5537 56516
rect 6271 56482 6305 56516
rect 7135 56482 7169 56516
rect 8575 56482 8609 56516
rect 10303 56482 10337 56516
rect 11071 56482 11105 56516
rect 11839 56482 11873 56516
rect 12607 56482 12641 56516
rect 13567 56482 13601 56516
rect 15007 56482 15041 56516
rect 17119 56482 17153 56516
rect 18175 56482 18209 56516
rect 18943 56482 18977 56516
rect 20287 56482 20321 56516
rect 21343 56482 21377 56516
rect 22111 56482 22145 56516
rect 22879 56482 22913 56516
rect 24319 56482 24353 56516
rect 26047 56482 26081 56516
rect 26911 56482 26945 56516
rect 27775 56482 27809 56516
rect 28543 56482 28577 56516
rect 29695 56482 29729 56516
rect 30847 56482 30881 56516
rect 31615 56482 31649 56516
rect 32383 56482 32417 56516
rect 33919 56482 33953 56516
rect 34783 56482 34817 56516
rect 36991 56482 37025 56516
rect 37663 56482 37697 56516
rect 38815 56482 38849 56516
rect 40159 56482 40193 56516
rect 41887 56482 41921 56516
rect 42751 56482 42785 56516
rect 43519 56482 43553 56516
rect 44287 56482 44321 56516
rect 45151 56482 45185 56516
rect 46687 56482 46721 56516
rect 48127 56482 48161 56516
rect 49759 56482 49793 56516
rect 50527 56482 50561 56516
rect 53023 56482 53057 56516
rect 53791 56482 53825 56516
rect 54463 56482 54497 56516
rect 55327 56482 55361 56516
rect 56095 56482 56129 56516
rect 4543 56334 4577 56368
rect 15487 56334 15521 56368
rect 15775 56334 15809 56368
rect 19039 56334 19073 56368
rect 1759 56260 1793 56294
rect 24415 56260 24449 56294
rect 52639 56260 52673 56294
rect 52927 56260 52961 56294
rect 55711 56260 55745 56294
rect 55999 56260 56033 56294
rect 57823 56260 57857 56294
rect 2527 56186 2561 56220
rect 3007 56186 3041 56220
rect 3295 56186 3329 56220
rect 5599 56186 5633 56220
rect 5983 56186 6017 56220
rect 6367 56186 6401 56220
rect 7231 56186 7265 56220
rect 8191 56186 8225 56220
rect 8479 56186 8513 56220
rect 10111 56186 10145 56220
rect 10399 56186 10433 56220
rect 11167 56186 11201 56220
rect 11935 56186 11969 56220
rect 12703 56186 12737 56220
rect 13279 56186 13313 56220
rect 13471 56186 13505 56220
rect 15103 56186 15137 56220
rect 15871 56186 15905 56220
rect 17215 56186 17249 56220
rect 18271 56186 18305 56220
rect 20383 56186 20417 56220
rect 21151 56186 21185 56220
rect 21439 56186 21473 56220
rect 21919 56186 21953 56220
rect 22207 56186 22241 56220
rect 22975 56186 23009 56220
rect 26143 56186 26177 56220
rect 26623 56186 26657 56220
rect 26815 56186 26849 56220
rect 27487 56186 27521 56220
rect 27679 56186 27713 56220
rect 28159 56186 28193 56220
rect 28447 56186 28481 56220
rect 29311 56186 29345 56220
rect 29599 56186 29633 56220
rect 30943 56186 30977 56220
rect 31423 56186 31457 56220
rect 31711 56186 31745 56220
rect 32479 56186 32513 56220
rect 32863 56186 32897 56220
rect 33151 56186 33185 56220
rect 33247 56186 33281 56220
rect 33727 56186 33761 56220
rect 34015 56186 34049 56220
rect 34399 56186 34433 56220
rect 34687 56186 34721 56220
rect 35839 56186 35873 56220
rect 36127 56186 36161 56220
rect 36223 56186 36257 56220
rect 36703 56186 36737 56220
rect 36895 56186 36929 56220
rect 37471 56186 37505 56220
rect 37759 56186 37793 56220
rect 38527 56186 38561 56220
rect 38719 56186 38753 56220
rect 39871 56186 39905 56220
rect 40255 56186 40289 56220
rect 41983 56186 42017 56220
rect 42463 56186 42497 56220
rect 42655 56186 42689 56220
rect 43231 56186 43265 56220
rect 43423 56186 43457 56220
rect 43999 56186 44033 56220
rect 44191 56186 44225 56220
rect 44863 56186 44897 56220
rect 45055 56186 45089 56220
rect 46783 56186 46817 56220
rect 48223 56186 48257 56220
rect 48703 56186 48737 56220
rect 48895 56186 48929 56220
rect 48991 56186 49025 56220
rect 49855 56186 49889 56220
rect 50623 56186 50657 56220
rect 51679 56186 51713 56220
rect 51967 56186 52001 56220
rect 52063 56186 52097 56220
rect 53503 56186 53537 56220
rect 53695 56186 53729 56220
rect 54559 56186 54593 56220
rect 55039 56186 55073 56220
rect 55231 56186 55265 56220
rect 55519 56186 55553 56220
rect 9727 55742 9761 55776
rect 9919 55742 9953 55776
rect 1663 55668 1697 55702
rect 4447 55668 4481 55702
rect 7615 55668 7649 55702
rect 9343 55668 9377 55702
rect 13951 55668 13985 55702
rect 20287 55668 20321 55702
rect 23551 55668 23585 55702
rect 25087 55668 25121 55702
rect 39295 55668 39329 55702
rect 40927 55668 40961 55702
rect 45631 55668 45665 55702
rect 47167 55668 47201 55702
rect 48031 55668 48065 55702
rect 51967 55668 52001 55702
rect 56671 55668 56705 55702
rect 57727 55668 57761 55702
rect 14047 55594 14081 55628
rect 1759 55520 1793 55554
rect 1951 55520 1985 55554
rect 4255 55520 4289 55554
rect 4543 55520 4577 55554
rect 7423 55520 7457 55554
rect 7711 55520 7745 55554
rect 9247 55520 9281 55554
rect 12511 55520 12545 55554
rect 12799 55520 12833 55554
rect 15295 55520 15329 55554
rect 15583 55520 15617 55554
rect 20383 55520 20417 55554
rect 23455 55520 23489 55554
rect 24991 55520 25025 55554
rect 25663 55520 25697 55554
rect 29119 55520 29153 55554
rect 39199 55520 39233 55554
rect 40831 55520 40865 55554
rect 41119 55520 41153 55554
rect 42559 55520 42593 55554
rect 45535 55520 45569 55554
rect 47071 55520 47105 55554
rect 47359 55520 47393 55554
rect 51871 55520 51905 55554
rect 55807 55520 55841 55554
rect 56575 55520 56609 55554
rect 57631 55520 57665 55554
rect 14719 55446 14753 55480
rect 8959 55372 8993 55406
rect 23167 55372 23201 55406
rect 24799 55372 24833 55406
rect 25567 55372 25601 55406
rect 38911 55372 38945 55406
rect 40543 55372 40577 55406
rect 42175 55372 42209 55406
rect 45247 55372 45281 55406
rect 46783 55372 46817 55406
rect 51583 55372 51617 55406
rect 55615 55372 55649 55406
rect 56287 55372 56321 55406
rect 57343 55372 57377 55406
rect 57823 55150 57857 55184
rect 12031 55002 12065 55036
rect 57631 54854 57665 54888
rect 57919 54854 57953 54888
rect 25855 54706 25889 54740
rect 26143 54706 26177 54740
rect 44671 54706 44705 54740
rect 44863 54706 44897 54740
rect 55807 54706 55841 54740
rect 55999 54706 56033 54740
rect 57919 54336 57953 54370
rect 14143 54188 14177 54222
rect 49087 54188 49121 54222
rect 49375 54188 49409 54222
rect 57631 54188 57665 54222
rect 57823 54188 57857 54222
rect 13855 54114 13889 54148
rect 57919 53818 57953 53852
rect 57823 53522 57857 53556
rect 26815 53374 26849 53408
rect 27007 53374 27041 53408
rect 57631 53374 57665 53408
rect 23935 52856 23969 52890
rect 24223 52856 24257 52890
rect 40831 52856 40865 52890
rect 41119 52856 41153 52890
rect 21343 52782 21377 52816
rect 23935 52708 23969 52742
rect 24031 52708 24065 52742
rect 37087 52190 37121 52224
rect 42847 52042 42881 52076
rect 43039 52042 43073 52076
rect 1663 51524 1697 51558
rect 1951 51524 1985 51558
rect 5695 51524 5729 51558
rect 5983 51524 6017 51558
rect 20095 51524 20129 51558
rect 19807 51450 19841 51484
rect 25375 50710 25409 50744
rect 25663 50710 25697 50744
rect 31519 50710 31553 50744
rect 31711 50710 31745 50744
rect 29791 50266 29825 50300
rect 30079 50266 30113 50300
rect 49183 50192 49217 50226
rect 57727 50192 57761 50226
rect 57823 50192 57857 50226
rect 49087 50044 49121 50078
rect 38143 49378 38177 49412
rect 38431 49378 38465 49412
rect 50335 49378 50369 49412
rect 50623 49378 50657 49412
rect 52063 49378 52097 49412
rect 40543 49156 40577 49190
rect 19135 48860 19169 48894
rect 19423 48860 19457 48894
rect 47839 48860 47873 48894
rect 47743 48712 47777 48746
rect 54943 48046 54977 48080
rect 55135 48046 55169 48080
rect 31423 47824 31457 47858
rect 27967 47602 28001 47636
rect 28255 47602 28289 47636
rect 54367 47528 54401 47562
rect 54463 47528 54497 47562
rect 6655 47158 6689 47192
rect 2719 46714 2753 46748
rect 3007 46714 3041 46748
rect 13087 46714 13121 46748
rect 13279 46714 13313 46748
rect 10879 46492 10913 46526
rect 24799 46270 24833 46304
rect 43711 46270 43745 46304
rect 43903 46270 43937 46304
rect 27967 46196 28001 46230
rect 28255 46196 28289 46230
rect 31423 46048 31457 46082
rect 6271 45382 6305 45416
rect 6559 45382 6593 45416
rect 41119 45382 41153 45416
rect 41311 45382 41345 45416
rect 44095 44864 44129 44898
rect 47551 44864 47585 44898
rect 47647 44864 47681 44898
rect 43903 44716 43937 44750
rect 12031 44124 12065 44158
rect 17119 44050 17153 44084
rect 17311 44050 17345 44084
rect 21631 43532 21665 43566
rect 21439 43384 21473 43418
rect 2143 42718 2177 42752
rect 2335 42718 2369 42752
rect 33247 42200 33281 42234
rect 33535 42200 33569 42234
rect 46495 42200 46529 42234
rect 30943 42126 30977 42160
rect 40159 42126 40193 42160
rect 46303 42052 46337 42086
rect 25375 41386 25409 41420
rect 25663 41386 25697 41420
rect 48319 41386 48353 41420
rect 15391 40942 15425 40976
rect 15679 40942 15713 40976
rect 22399 40942 22433 40976
rect 1759 40868 1793 40902
rect 17407 40868 17441 40902
rect 17695 40868 17729 40902
rect 22399 40794 22433 40828
rect 1951 40720 1985 40754
rect 2815 40350 2849 40384
rect 32959 40054 32993 40088
rect 33151 40054 33185 40088
rect 49183 39536 49217 39570
rect 48991 39388 49025 39422
rect 58015 38796 58049 38830
rect 12319 38722 12353 38756
rect 12607 38722 12641 38756
rect 24127 38722 24161 38756
rect 52351 38722 52385 38756
rect 52543 38722 52577 38756
rect 10879 38204 10913 38238
rect 12799 38204 12833 38238
rect 13087 38204 13121 38238
rect 10687 38056 10721 38090
rect 10015 37538 10049 37572
rect 10303 37390 10337 37424
rect 11455 37390 11489 37424
rect 29503 37390 29537 37424
rect 29599 37390 29633 37424
rect 5023 37168 5057 37202
rect 33823 36872 33857 36906
rect 34111 36872 34145 36906
rect 2431 36502 2465 36536
rect 7327 36132 7361 36166
rect 16447 36058 16481 36092
rect 16831 36058 16865 36092
rect 13279 35540 13313 35574
rect 39103 35540 39137 35574
rect 43903 35540 43937 35574
rect 13087 35392 13121 35426
rect 43711 35392 43745 35426
rect 33151 35022 33185 35056
rect 51679 34874 51713 34908
rect 51871 34874 51905 34908
rect 6079 34800 6113 34834
rect 22783 34800 22817 34834
rect 22975 34800 23009 34834
rect 52351 34800 52385 34834
rect 52543 34800 52577 34834
rect 21055 34726 21089 34760
rect 21343 34726 21377 34760
rect 28543 34726 28577 34760
rect 28735 34726 28769 34760
rect 22975 34208 23009 34242
rect 55807 34208 55841 34242
rect 28159 33542 28193 33576
rect 28351 33542 28385 33576
rect 57631 33468 57665 33502
rect 17119 33394 17153 33428
rect 17311 33394 17345 33428
rect 18751 33394 18785 33428
rect 43135 33394 43169 33428
rect 44767 33172 44801 33206
rect 2527 33024 2561 33058
rect 46783 32950 46817 32984
rect 46975 32950 47009 32984
rect 40063 32876 40097 32910
rect 39871 32728 39905 32762
rect 8479 32136 8513 32170
rect 32191 32062 32225 32096
rect 43039 32062 43073 32096
rect 21343 31692 21377 31726
rect 34687 31692 34721 31726
rect 29023 31618 29057 31652
rect 54751 31026 54785 31060
rect 7999 30730 8033 30764
rect 8287 30730 8321 30764
rect 16159 30286 16193 30320
rect 5791 29620 5825 29654
rect 6079 29620 6113 29654
rect 18367 29398 18401 29432
rect 47359 28806 47393 28840
rect 47551 28732 47585 28766
rect 31039 28214 31073 28248
rect 31231 28214 31265 28248
rect 9919 28066 9953 28100
rect 21343 28066 21377 28100
rect 57343 28066 57377 28100
rect 14431 27844 14465 27878
rect 14623 27844 14657 27878
rect 5311 27548 5345 27582
rect 57727 27548 57761 27582
rect 38623 27178 38657 27212
rect 38815 27030 38849 27064
rect 42271 26808 42305 26842
rect 15103 26734 15137 26768
rect 36223 26734 36257 26768
rect 1951 26512 1985 26546
rect 8767 26438 8801 26472
rect 8383 26364 8417 26398
rect 57727 26216 57761 26250
rect 57823 26216 57857 26250
rect 25375 25550 25409 25584
rect 25663 25550 25697 25584
rect 33535 25476 33569 25510
rect 26815 24884 26849 24918
rect 33535 24884 33569 24918
rect 51295 24884 51329 24918
rect 10495 24070 10529 24104
rect 36607 24070 36641 24104
rect 41503 24070 41537 24104
rect 19903 23626 19937 23660
rect 20191 23626 20225 23660
rect 29983 23552 30017 23586
rect 30079 23552 30113 23586
rect 41791 23552 41825 23586
rect 44671 23552 44705 23586
rect 46975 23552 47009 23586
rect 30079 23404 30113 23438
rect 10207 22738 10241 22772
rect 37567 22738 37601 22772
rect 8191 22516 8225 22550
rect 7615 22072 7649 22106
rect 8095 22072 8129 22106
rect 7999 21628 8033 21662
rect 8287 21628 8321 21662
rect 32863 21406 32897 21440
rect 7615 20740 7649 20774
rect 24031 20148 24065 20182
rect 24319 20148 24353 20182
rect 16159 20074 16193 20108
rect 27583 20074 27617 20108
rect 7615 19852 7649 19886
rect 6847 19556 6881 19590
rect 7135 19556 7169 19590
rect 34783 19556 34817 19590
rect 48703 18890 48737 18924
rect 48895 18890 48929 18924
rect 21247 18742 21281 18776
rect 52063 18742 52097 18776
rect 7615 18520 7649 18554
rect 7903 18520 7937 18554
rect 8191 18520 8225 18554
rect 1759 18224 1793 18258
rect 24511 18224 24545 18258
rect 40735 18224 40769 18258
rect 51199 18224 51233 18258
rect 26143 18076 26177 18110
rect 26431 18076 26465 18110
rect 51007 18076 51041 18110
rect 30655 17632 30689 17666
rect 30943 17632 30977 17666
rect 1951 17410 1985 17444
rect 56767 16966 56801 17000
rect 5983 16892 6017 16926
rect 7135 16892 7169 16926
rect 46879 16892 46913 16926
rect 55999 16892 56033 16926
rect 7615 16744 7649 16778
rect 27103 16078 27137 16112
rect 46879 15560 46913 15594
rect 47071 15560 47105 15594
rect 7615 15412 7649 15446
rect 12319 15190 12353 15224
rect 12607 15190 12641 15224
rect 24031 15190 24065 15224
rect 24223 15042 24257 15076
rect 57727 15042 57761 15076
rect 58015 15042 58049 15076
rect 23743 14820 23777 14854
rect 3583 14524 3617 14558
rect 3871 14524 3905 14558
rect 12703 14450 12737 14484
rect 17503 14376 17537 14410
rect 17791 14376 17825 14410
rect 4447 14080 4481 14114
rect 4735 14080 4769 14114
rect 7615 14080 7649 14114
rect 47647 13710 47681 13744
rect 15103 13414 15137 13448
rect 47359 13414 47393 13448
rect 7615 13192 7649 13226
rect 26719 13118 26753 13152
rect 48991 13044 49025 13078
rect 49183 13044 49217 13078
rect 58015 12970 58049 13004
rect 57727 12378 57761 12412
rect 31327 12230 31361 12264
rect 57631 12230 57665 12264
rect 31039 12156 31073 12190
rect 5023 12082 5057 12116
rect 15199 12082 15233 12116
rect 18751 12082 18785 12116
rect 29599 12082 29633 12116
rect 1759 11860 1793 11894
rect 1855 11860 1889 11894
rect 5215 11860 5249 11894
rect 7615 11860 7649 11894
rect 56479 11712 56513 11746
rect 9247 11638 9281 11672
rect 9535 11638 9569 11672
rect 56959 11638 56993 11672
rect 57247 11638 57281 11672
rect 37663 11564 37697 11598
rect 54655 11564 54689 11598
rect 56575 11564 56609 11598
rect 57343 11416 57377 11450
rect 55807 11046 55841 11080
rect 55999 11046 56033 11080
rect 56287 11046 56321 11080
rect 56959 10972 56993 11006
rect 57247 10972 57281 11006
rect 56095 10898 56129 10932
rect 57343 10898 57377 10932
rect 12127 10750 12161 10784
rect 7615 10528 7649 10562
rect 56383 10528 56417 10562
rect 56863 10528 56897 10562
rect 57055 10454 57089 10488
rect 55039 10380 55073 10414
rect 55135 10380 55169 10414
rect 56671 10380 56705 10414
rect 57343 10380 57377 10414
rect 29215 10306 29249 10340
rect 28447 10232 28481 10266
rect 41503 10232 41537 10266
rect 55807 10232 55841 10266
rect 56575 10232 56609 10266
rect 55519 10158 55553 10192
rect 55903 10084 55937 10118
rect 57439 10084 57473 10118
rect 55903 9862 55937 9896
rect 55999 9714 56033 9748
rect 55231 9640 55265 9674
rect 57631 9640 57665 9674
rect 54367 9566 54401 9600
rect 54463 9566 54497 9600
rect 55135 9566 55169 9600
rect 25855 9418 25889 9452
rect 32383 9418 32417 9452
rect 53023 9196 53057 9230
rect 55135 9196 55169 9230
rect 55615 9196 55649 9230
rect 5311 9122 5345 9156
rect 5599 9122 5633 9156
rect 53311 9048 53345 9082
rect 53407 9048 53441 9082
rect 55423 9048 55457 9082
rect 55327 8974 55361 9008
rect 56575 8974 56609 9008
rect 57247 8974 57281 9008
rect 25663 8900 25697 8934
rect 54559 8900 54593 8934
rect 54271 8826 54305 8860
rect 7615 8752 7649 8786
rect 54655 8752 54689 8786
rect 1951 8530 1985 8564
rect 7039 8530 7073 8564
rect 9535 8530 9569 8564
rect 13567 8530 13601 8564
rect 48607 8530 48641 8564
rect 52447 8530 52481 8564
rect 1759 8382 1793 8416
rect 2527 8382 2561 8416
rect 7615 8382 7649 8416
rect 7903 8382 7937 8416
rect 9823 8382 9857 8416
rect 11071 8382 11105 8416
rect 11359 8382 11393 8416
rect 13663 8382 13697 8416
rect 16255 8382 16289 8416
rect 17023 8382 17057 8416
rect 38431 8382 38465 8416
rect 38623 8382 38657 8416
rect 47935 8382 47969 8416
rect 48127 8382 48161 8416
rect 48895 8382 48929 8416
rect 49759 8382 49793 8416
rect 52543 8382 52577 8416
rect 53023 8382 53057 8416
rect 53215 8382 53249 8416
rect 54079 8382 54113 8416
rect 3295 8308 3329 8342
rect 7039 8308 7073 8342
rect 12127 8308 12161 8342
rect 12895 8308 12929 8342
rect 55231 8308 55265 8342
rect 55999 8308 56033 8342
rect 57151 8308 57185 8342
rect 1663 8234 1697 8268
rect 2431 8234 2465 8268
rect 3199 8234 3233 8268
rect 4447 8234 4481 8268
rect 4543 8234 4577 8268
rect 7807 8234 7841 8268
rect 9727 8234 9761 8268
rect 10495 8234 10529 8268
rect 10591 8234 10625 8268
rect 11263 8234 11297 8268
rect 12031 8234 12065 8268
rect 12799 8234 12833 8268
rect 16159 8234 16193 8268
rect 16927 8234 16961 8268
rect 48223 8234 48257 8268
rect 48991 8234 49025 8268
rect 49663 8234 49697 8268
rect 53311 8234 53345 8268
rect 53983 8234 54017 8268
rect 10207 8160 10241 8194
rect 25663 8160 25697 8194
rect 4255 8086 4289 8120
rect 5503 8086 5537 8120
rect 18367 8086 18401 8120
rect 29599 8086 29633 8120
rect 45151 8086 45185 8120
rect 36511 7864 36545 7898
rect 40831 7864 40865 7898
rect 42271 7864 42305 7898
rect 45247 7864 45281 7898
rect 46111 7864 46145 7898
rect 47551 7864 47585 7898
rect 48991 7864 49025 7898
rect 53023 7864 53057 7898
rect 2239 7790 2273 7824
rect 7615 7790 7649 7824
rect 2527 7716 2561 7750
rect 3295 7716 3329 7750
rect 10111 7716 10145 7750
rect 13087 7716 13121 7750
rect 13663 7716 13697 7750
rect 13951 7716 13985 7750
rect 20671 7716 20705 7750
rect 20959 7716 20993 7750
rect 23647 7716 23681 7750
rect 23935 7716 23969 7750
rect 25471 7716 25505 7750
rect 26239 7716 26273 7750
rect 27007 7716 27041 7750
rect 28063 7716 28097 7750
rect 28351 7716 28385 7750
rect 29407 7716 29441 7750
rect 30175 7716 30209 7750
rect 31231 7716 31265 7750
rect 34591 7716 34625 7750
rect 35359 7716 35393 7750
rect 36127 7716 36161 7750
rect 36799 7716 36833 7750
rect 40351 7716 40385 7750
rect 41023 7716 41057 7750
rect 41887 7716 41921 7750
rect 42559 7716 42593 7750
rect 44095 7716 44129 7750
rect 44575 7716 44609 7750
rect 44863 7716 44897 7750
rect 45631 7716 45665 7750
rect 46399 7716 46433 7750
rect 47167 7716 47201 7750
rect 47839 7716 47873 7750
rect 49375 7716 49409 7750
rect 51583 7716 51617 7750
rect 51775 7716 51809 7750
rect 52639 7716 52673 7750
rect 53407 7716 53441 7750
rect 1567 7642 1601 7676
rect 3775 7642 3809 7676
rect 4063 7642 4097 7676
rect 4831 7642 4865 7676
rect 9055 7642 9089 7676
rect 9439 7642 9473 7676
rect 10207 7642 10241 7676
rect 12415 7642 12449 7676
rect 14815 7642 14849 7676
rect 15103 7642 15137 7676
rect 15871 7642 15905 7676
rect 29887 7642 29921 7676
rect 30079 7642 30113 7676
rect 46303 7642 46337 7676
rect 49279 7642 49313 7676
rect 51103 7642 51137 7676
rect 53311 7642 53345 7676
rect 55135 7642 55169 7676
rect 55807 7642 55841 7676
rect 56575 7642 56609 7676
rect 57343 7642 57377 7676
rect 5599 7568 5633 7602
rect 10687 7568 10721 7602
rect 10975 7568 11009 7602
rect 13183 7568 13217 7602
rect 24703 7568 24737 7602
rect 33823 7568 33857 7602
rect 38815 7568 38849 7602
rect 39583 7568 39617 7602
rect 41119 7568 41153 7602
rect 45535 7568 45569 7602
rect 49759 7568 49793 7602
rect 50047 7568 50081 7602
rect 2431 7420 2465 7454
rect 3199 7420 3233 7454
rect 3967 7420 4001 7454
rect 4735 7420 4769 7454
rect 5503 7420 5537 7454
rect 9343 7420 9377 7454
rect 10879 7420 10913 7454
rect 12319 7420 12353 7454
rect 13855 7420 13889 7454
rect 15775 7420 15809 7454
rect 20863 7420 20897 7454
rect 23839 7420 23873 7454
rect 24607 7420 24641 7454
rect 25375 7420 25409 7454
rect 26143 7420 26177 7454
rect 26911 7420 26945 7454
rect 28255 7420 28289 7454
rect 29311 7420 29345 7454
rect 31135 7420 31169 7454
rect 33727 7420 33761 7454
rect 34495 7420 34529 7454
rect 35263 7420 35297 7454
rect 36031 7420 36065 7454
rect 36895 7420 36929 7454
rect 38719 7420 38753 7454
rect 39487 7420 39521 7454
rect 40255 7420 40289 7454
rect 41791 7420 41825 7454
rect 42655 7420 42689 7454
rect 43999 7420 44033 7454
rect 44767 7420 44801 7454
rect 47071 7420 47105 7454
rect 47935 7420 47969 7454
rect 50143 7420 50177 7454
rect 51007 7420 51041 7454
rect 51871 7420 51905 7454
rect 52543 7420 52577 7454
rect 10303 7124 10337 7158
rect 20767 7124 20801 7158
rect 23935 7124 23969 7158
rect 26815 7124 26849 7158
rect 29119 7124 29153 7158
rect 36607 7124 36641 7158
rect 37471 7124 37505 7158
rect 39679 7124 39713 7158
rect 41119 7124 41153 7158
rect 41887 7124 41921 7158
rect 43423 7124 43457 7158
rect 45055 7124 45089 7158
rect 48799 7124 48833 7158
rect 52447 7124 52481 7158
rect 4543 7050 4577 7084
rect 5791 7050 5825 7084
rect 6079 7050 6113 7084
rect 15871 7050 15905 7084
rect 17023 7050 17057 7084
rect 17311 7050 17345 7084
rect 17791 7050 17825 7084
rect 18079 7050 18113 7084
rect 18847 7050 18881 7084
rect 20095 7050 20129 7084
rect 20383 7050 20417 7084
rect 21055 7050 21089 7084
rect 21919 7050 21953 7084
rect 22399 7050 22433 7084
rect 22687 7050 22721 7084
rect 24223 7050 24257 7084
rect 25663 7050 25697 7084
rect 26431 7050 26465 7084
rect 27103 7050 27137 7084
rect 27679 7050 27713 7084
rect 27967 7050 28001 7084
rect 28735 7050 28769 7084
rect 29407 7050 29441 7084
rect 30943 7050 30977 7084
rect 31711 7050 31745 7084
rect 32191 7050 32225 7084
rect 32383 7050 32417 7084
rect 32959 7050 32993 7084
rect 33247 7050 33281 7084
rect 34783 7050 34817 7084
rect 36223 7050 36257 7084
rect 36895 7050 36929 7084
rect 37759 7050 37793 7084
rect 38527 7050 38561 7084
rect 39295 7050 39329 7084
rect 39967 7050 40001 7084
rect 41407 7050 41441 7084
rect 42175 7050 42209 7084
rect 42751 7050 42785 7084
rect 42943 7050 42977 7084
rect 43807 7050 43841 7084
rect 45247 7050 45281 7084
rect 46495 7050 46529 7084
rect 46687 7050 46721 7084
rect 47551 7050 47585 7084
rect 48319 7050 48353 7084
rect 48991 7050 49025 7084
rect 50047 7050 50081 7084
rect 50239 7050 50273 7084
rect 52063 7050 52097 7084
rect 52735 7050 52769 7084
rect 1663 6976 1697 7010
rect 2527 6976 2561 7010
rect 5023 6976 5057 7010
rect 5311 6976 5345 7010
rect 6463 6976 6497 7010
rect 6847 6976 6881 7010
rect 7615 6976 7649 7010
rect 8095 6976 8129 7010
rect 10591 6976 10625 7010
rect 11263 6976 11297 7010
rect 12703 6976 12737 7010
rect 15103 6976 15137 7010
rect 23455 6976 23489 7010
rect 34015 6976 34049 7010
rect 44287 6976 44321 7010
rect 44575 6976 44609 7010
rect 54079 6976 54113 7010
rect 54751 6976 54785 7010
rect 55519 6976 55553 7010
rect 57823 6976 57857 7010
rect 4447 6902 4481 6936
rect 5215 6902 5249 6936
rect 5983 6902 6017 6936
rect 6751 6902 6785 6936
rect 7519 6902 7553 6936
rect 8287 6902 8321 6936
rect 8383 6902 8417 6936
rect 9727 6902 9761 6936
rect 9823 6902 9857 6936
rect 10495 6902 10529 6936
rect 13567 6902 13601 6936
rect 13663 6902 13697 6936
rect 15007 6902 15041 6936
rect 15775 6902 15809 6936
rect 17215 6902 17249 6936
rect 17983 6902 18017 6936
rect 18751 6902 18785 6936
rect 20287 6902 20321 6936
rect 21151 6902 21185 6936
rect 21823 6902 21857 6936
rect 22591 6902 22625 6936
rect 23359 6902 23393 6936
rect 24127 6902 24161 6936
rect 25567 6902 25601 6936
rect 26335 6902 26369 6936
rect 27199 6902 27233 6936
rect 27871 6902 27905 6936
rect 28639 6902 28673 6936
rect 29503 6902 29537 6936
rect 30847 6902 30881 6936
rect 31615 6902 31649 6936
rect 32479 6902 32513 6936
rect 33151 6902 33185 6936
rect 33919 6902 33953 6936
rect 34687 6902 34721 6936
rect 36127 6902 36161 6936
rect 36991 6902 37025 6936
rect 37663 6902 37697 6936
rect 38431 6902 38465 6936
rect 39199 6902 39233 6936
rect 40063 6902 40097 6936
rect 41503 6902 41537 6936
rect 42271 6902 42305 6936
rect 43039 6902 43073 6936
rect 43711 6902 43745 6936
rect 44479 6902 44513 6936
rect 45343 6902 45377 6936
rect 46783 6902 46817 6936
rect 47455 6902 47489 6936
rect 48223 6902 48257 6936
rect 49087 6902 49121 6936
rect 50335 6902 50369 6936
rect 51967 6902 52001 6936
rect 52831 6902 52865 6936
rect 5407 6532 5441 6566
rect 15967 6532 16001 6566
rect 30271 6532 30305 6566
rect 31807 6532 31841 6566
rect 34783 6532 34817 6566
rect 36895 6532 36929 6566
rect 51295 6532 51329 6566
rect 7615 6458 7649 6492
rect 13663 6458 13697 6492
rect 39871 6458 39905 6492
rect 5695 6384 5729 6418
rect 7135 6384 7169 6418
rect 13855 6384 13889 6418
rect 13951 6384 13985 6418
rect 15487 6384 15521 6418
rect 16255 6384 16289 6418
rect 17407 6384 17441 6418
rect 17695 6384 17729 6418
rect 18463 6384 18497 6418
rect 18943 6384 18977 6418
rect 19135 6384 19169 6418
rect 19711 6384 19745 6418
rect 19999 6384 20033 6418
rect 20767 6384 20801 6418
rect 21535 6384 21569 6418
rect 23743 6384 23777 6418
rect 24223 6384 24257 6418
rect 24511 6384 24545 6418
rect 28255 6384 28289 6418
rect 29023 6384 29057 6418
rect 30559 6384 30593 6418
rect 32095 6384 32129 6418
rect 32191 6384 32225 6418
rect 33535 6384 33569 6418
rect 34015 6384 34049 6418
rect 34207 6384 34241 6418
rect 34975 6384 35009 6418
rect 37279 6384 37313 6418
rect 42559 6384 42593 6418
rect 42751 6384 42785 6418
rect 44863 6384 44897 6418
rect 50911 6384 50945 6418
rect 51583 6384 51617 6418
rect 52447 6384 52481 6418
rect 1567 6310 1601 6344
rect 2335 6310 2369 6344
rect 3199 6310 3233 6344
rect 3967 6310 4001 6344
rect 4735 6310 4769 6344
rect 9439 6310 9473 6344
rect 10207 6310 10241 6344
rect 10975 6310 11009 6344
rect 12223 6310 12257 6344
rect 12991 6310 13025 6344
rect 22975 6310 23009 6344
rect 25663 6310 25697 6344
rect 26815 6310 26849 6344
rect 29695 6310 29729 6344
rect 31231 6310 31265 6344
rect 36319 6310 36353 6344
rect 38911 6310 38945 6344
rect 40351 6310 40385 6344
rect 41887 6310 41921 6344
rect 45535 6310 45569 6344
rect 46975 6310 47009 6344
rect 47743 6310 47777 6344
rect 49183 6310 49217 6344
rect 49951 6310 49985 6344
rect 53311 6310 53345 6344
rect 54463 6310 54497 6344
rect 55231 6310 55265 6344
rect 55999 6310 56033 6344
rect 57055 6310 57089 6344
rect 57823 6310 57857 6344
rect 14719 6236 14753 6270
rect 41311 6236 41345 6270
rect 44095 6236 44129 6270
rect 5599 6088 5633 6122
rect 7039 6088 7073 6122
rect 14623 6088 14657 6122
rect 15391 6088 15425 6122
rect 16159 6088 16193 6122
rect 17599 6088 17633 6122
rect 18367 6088 18401 6122
rect 19231 6088 19265 6122
rect 19903 6088 19937 6122
rect 20671 6088 20705 6122
rect 21439 6088 21473 6122
rect 22879 6088 22913 6122
rect 23647 6088 23681 6122
rect 24415 6088 24449 6122
rect 28159 6088 28193 6122
rect 28927 6088 28961 6122
rect 30655 6088 30689 6122
rect 33439 6088 33473 6122
rect 34303 6088 34337 6122
rect 35071 6088 35105 6122
rect 37183 6088 37217 6122
rect 41215 6088 41249 6122
rect 42847 6088 42881 6122
rect 43999 6088 44033 6122
rect 44767 6088 44801 6122
rect 50815 6088 50849 6122
rect 51679 6088 51713 6122
rect 52351 6088 52385 6122
rect 55423 5718 55457 5752
rect 1567 5644 1601 5678
rect 2911 5644 2945 5678
rect 4447 5644 4481 5678
rect 5119 5644 5153 5678
rect 6847 5644 6881 5678
rect 7615 5644 7649 5678
rect 7999 5644 8033 5678
rect 8383 5644 8417 5678
rect 9631 5644 9665 5678
rect 10399 5644 10433 5678
rect 11167 5644 11201 5678
rect 12607 5644 12641 5678
rect 13375 5644 13409 5678
rect 15007 5644 15041 5678
rect 15871 5644 15905 5678
rect 16543 5644 16577 5678
rect 17311 5644 17345 5678
rect 18751 5644 18785 5678
rect 20191 5644 20225 5678
rect 20959 5644 20993 5678
rect 21631 5644 21665 5678
rect 21727 5644 21761 5678
rect 22495 5644 22529 5678
rect 23263 5644 23297 5678
rect 24031 5644 24065 5678
rect 25471 5644 25505 5678
rect 26239 5644 26273 5678
rect 26623 5644 26657 5678
rect 27007 5644 27041 5678
rect 27775 5644 27809 5678
rect 28543 5644 28577 5678
rect 29311 5644 29345 5678
rect 30751 5644 30785 5678
rect 31519 5644 31553 5678
rect 32287 5644 32321 5678
rect 33151 5644 33185 5678
rect 33823 5644 33857 5678
rect 34687 5644 34721 5678
rect 36031 5644 36065 5678
rect 36799 5644 36833 5678
rect 37567 5644 37601 5678
rect 37951 5644 37985 5678
rect 38335 5644 38369 5678
rect 39103 5644 39137 5678
rect 39871 5644 39905 5678
rect 41311 5644 41345 5678
rect 42079 5644 42113 5678
rect 42847 5644 42881 5678
rect 43615 5644 43649 5678
rect 44383 5644 44417 5678
rect 45151 5644 45185 5678
rect 46591 5644 46625 5678
rect 47359 5644 47393 5678
rect 48127 5644 48161 5678
rect 48991 5644 49025 5678
rect 49663 5644 49697 5678
rect 50527 5644 50561 5678
rect 52159 5644 52193 5678
rect 52927 5644 52961 5678
rect 53695 5644 53729 5678
rect 54463 5644 54497 5678
rect 55999 5644 56033 5678
rect 57439 5644 57473 5678
rect 5983 5570 6017 5604
rect 6079 5570 6113 5604
rect 5791 5496 5825 5530
rect 7999 5496 8033 5530
rect 21631 5496 21665 5530
rect 26623 5496 26657 5530
rect 37951 5496 37985 5530
rect 7519 5200 7553 5234
rect 7711 5200 7745 5234
rect 8479 5200 8513 5234
rect 1567 4978 1601 5012
rect 2335 4978 2369 5012
rect 3103 4978 3137 5012
rect 4159 4978 4193 5012
rect 5407 4978 5441 5012
rect 6943 4978 6977 5012
rect 9247 4978 9281 5012
rect 10015 4978 10049 5012
rect 10783 4978 10817 5012
rect 12223 4978 12257 5012
rect 12991 4978 13025 5012
rect 13951 4978 13985 5012
rect 14719 4978 14753 5012
rect 15487 4978 15521 5012
rect 16351 4978 16385 5012
rect 17503 4978 17537 5012
rect 18271 4978 18305 5012
rect 19039 4978 19073 5012
rect 19807 4978 19841 5012
rect 20575 4978 20609 5012
rect 21343 4978 21377 5012
rect 22783 4978 22817 5012
rect 23551 4978 23585 5012
rect 24319 4978 24353 5012
rect 25087 4978 25121 5012
rect 25855 4978 25889 5012
rect 26623 4978 26657 5012
rect 28063 4978 28097 5012
rect 28927 4978 28961 5012
rect 29599 4978 29633 5012
rect 30367 4978 30401 5012
rect 31135 4978 31169 5012
rect 31903 4978 31937 5012
rect 33343 4978 33377 5012
rect 34111 4978 34145 5012
rect 34879 4978 34913 5012
rect 35647 4978 35681 5012
rect 36415 4978 36449 5012
rect 37183 4978 37217 5012
rect 38623 4978 38657 5012
rect 39391 4978 39425 5012
rect 40159 4978 40193 5012
rect 40927 4978 40961 5012
rect 41695 4978 41729 5012
rect 42463 4978 42497 5012
rect 43903 4978 43937 5012
rect 44767 4978 44801 5012
rect 45439 4978 45473 5012
rect 46207 4978 46241 5012
rect 46975 4978 47009 5012
rect 47743 4978 47777 5012
rect 49375 4978 49409 5012
rect 50431 4978 50465 5012
rect 51103 4978 51137 5012
rect 51871 4978 51905 5012
rect 52639 4978 52673 5012
rect 54463 4978 54497 5012
rect 55615 4978 55649 5012
rect 56383 4978 56417 5012
rect 57055 4978 57089 5012
rect 15775 4534 15809 4568
rect 16543 4460 16577 4494
rect 1567 4312 1601 4346
rect 2335 4312 2369 4346
rect 3103 4312 3137 4346
rect 4351 4312 4385 4346
rect 5119 4312 5153 4346
rect 5887 4312 5921 4346
rect 6655 4312 6689 4346
rect 7423 4312 7457 4346
rect 8191 4312 8225 4346
rect 9631 4312 9665 4346
rect 10399 4312 10433 4346
rect 11167 4312 11201 4346
rect 11935 4312 11969 4346
rect 12703 4312 12737 4346
rect 13567 4312 13601 4346
rect 15487 4312 15521 4346
rect 16255 4312 16289 4346
rect 17023 4312 17057 4346
rect 17791 4312 17825 4346
rect 18559 4312 18593 4346
rect 20287 4312 20321 4346
rect 21055 4312 21089 4346
rect 21823 4312 21857 4346
rect 23263 4312 23297 4346
rect 24031 4312 24065 4346
rect 25471 4312 25505 4346
rect 26239 4312 26273 4346
rect 27007 4312 27041 4346
rect 28351 4312 28385 4346
rect 29119 4312 29153 4346
rect 30943 4312 30977 4346
rect 31711 4312 31745 4346
rect 32767 4312 32801 4346
rect 33919 4312 33953 4346
rect 34687 4312 34721 4346
rect 36031 4312 36065 4346
rect 36799 4312 36833 4346
rect 37567 4312 37601 4346
rect 39007 4312 39041 4346
rect 39775 4312 39809 4346
rect 41983 4312 42017 4346
rect 42751 4312 42785 4346
rect 43519 4312 43553 4346
rect 44959 4312 44993 4346
rect 46783 4312 46817 4346
rect 47551 4312 47585 4346
rect 48319 4312 48353 4346
rect 49087 4312 49121 4346
rect 49855 4312 49889 4346
rect 50623 4312 50657 4346
rect 51871 4312 51905 4346
rect 52639 4312 52673 4346
rect 53407 4312 53441 4346
rect 54175 4312 54209 4346
rect 55615 4312 55649 4346
rect 57151 4312 57185 4346
rect 44479 4238 44513 4272
rect 41503 4090 41537 4124
rect 12415 3868 12449 3902
rect 13951 3868 13985 3902
rect 15487 3868 15521 3902
rect 18559 3868 18593 3902
rect 1567 3646 1601 3680
rect 2335 3646 2369 3680
rect 3103 3646 3137 3680
rect 3871 3646 3905 3680
rect 4639 3646 4673 3680
rect 5599 3646 5633 3680
rect 6943 3646 6977 3680
rect 7711 3646 7745 3680
rect 8479 3646 8513 3680
rect 9247 3646 9281 3680
rect 10015 3646 10049 3680
rect 10783 3646 10817 3680
rect 12991 3646 13025 3680
rect 13663 3646 13697 3680
rect 14431 3646 14465 3680
rect 15199 3646 15233 3680
rect 15967 3646 16001 3680
rect 17503 3646 17537 3680
rect 18271 3646 18305 3680
rect 19039 3646 19073 3680
rect 19807 3646 19841 3680
rect 20575 3646 20609 3680
rect 21343 3646 21377 3680
rect 22783 3646 22817 3680
rect 23551 3646 23585 3680
rect 24319 3646 24353 3680
rect 25087 3646 25121 3680
rect 25855 3646 25889 3680
rect 26623 3646 26657 3680
rect 28063 3646 28097 3680
rect 28831 3646 28865 3680
rect 29695 3646 29729 3680
rect 30367 3646 30401 3680
rect 31135 3646 31169 3680
rect 31903 3646 31937 3680
rect 33343 3646 33377 3680
rect 34111 3646 34145 3680
rect 34879 3646 34913 3680
rect 35647 3646 35681 3680
rect 36415 3646 36449 3680
rect 37183 3646 37217 3680
rect 38623 3646 38657 3680
rect 39391 3646 39425 3680
rect 40159 3646 40193 3680
rect 40927 3646 40961 3680
rect 41695 3646 41729 3680
rect 42463 3646 42497 3680
rect 43903 3646 43937 3680
rect 44671 3646 44705 3680
rect 45439 3646 45473 3680
rect 46207 3646 46241 3680
rect 46975 3646 47009 3680
rect 47743 3646 47777 3680
rect 49183 3646 49217 3680
rect 50527 3646 50561 3680
rect 51199 3646 51233 3680
rect 51967 3646 52001 3680
rect 52735 3646 52769 3680
rect 54463 3646 54497 3680
rect 55231 3646 55265 3680
rect 55999 3646 56033 3680
rect 56767 3646 56801 3680
rect 57535 3646 57569 3680
rect 13279 3202 13313 3236
rect 14047 3202 14081 3236
rect 15391 3202 15425 3236
rect 16831 3202 16865 3236
rect 18079 3202 18113 3236
rect 18847 3202 18881 3236
rect 21151 3054 21185 3088
rect 24607 3054 24641 3088
rect 24895 3054 24929 3088
rect 1567 2980 1601 3014
rect 2335 2980 2369 3014
rect 3103 2980 3137 3014
rect 4927 2980 4961 3014
rect 5695 2980 5729 3014
rect 7039 2980 7073 3014
rect 7807 2980 7841 3014
rect 9727 2980 9761 3014
rect 10495 2980 10529 3014
rect 12991 2980 13025 3014
rect 13759 2980 13793 3014
rect 15103 2980 15137 3014
rect 16639 2980 16673 3014
rect 17791 2980 17825 3014
rect 18559 2980 18593 3014
rect 20479 2980 20513 3014
rect 8479 2906 8513 2940
rect 21247 2980 21281 3014
rect 23167 2980 23201 3014
rect 23935 2980 23969 3014
rect 25855 2980 25889 3014
rect 26623 2980 26657 3014
rect 28543 2980 28577 3014
rect 29311 2980 29345 3014
rect 31231 2980 31265 3014
rect 31999 2980 32033 3014
rect 33919 2980 33953 3014
rect 34687 2980 34721 3014
rect 36607 2980 36641 3014
rect 37375 2980 37409 3014
rect 39295 2980 39329 3014
rect 40063 2980 40097 3014
rect 41983 2980 42017 3014
rect 42751 2980 42785 3014
rect 44671 2980 44705 3014
rect 45439 2980 45473 3014
rect 47359 2980 47393 3014
rect 48127 2980 48161 3014
rect 50047 2980 50081 3014
rect 50815 2980 50849 3014
rect 52735 2980 52769 3014
rect 53503 2980 53537 3014
rect 55423 2980 55457 3014
rect 56191 2980 56225 3014
rect 27295 2906 27329 2940
rect 8767 2832 8801 2866
rect 11455 2832 11489 2866
rect 21151 2832 21185 2866
rect 27583 2832 27617 2866
rect 30271 2832 30305 2866
rect 38335 2832 38369 2866
rect 41023 2758 41057 2792
rect 46399 2758 46433 2792
rect 49087 2758 49121 2792
<< metal1 >>
rect 1152 57302 58848 57324
rect 1152 57250 4294 57302
rect 4346 57250 4358 57302
rect 4410 57250 4422 57302
rect 4474 57250 4486 57302
rect 4538 57250 35014 57302
rect 35066 57250 35078 57302
rect 35130 57250 35142 57302
rect 35194 57250 35206 57302
rect 35258 57250 58848 57302
rect 1152 57228 58848 57250
rect 1744 56991 1750 57043
rect 1802 57031 1808 57043
rect 1802 57003 2846 57031
rect 1802 56991 1808 57003
rect 208 56917 214 56969
rect 266 56957 272 56969
rect 2818 56966 2846 57003
rect 3280 56991 3286 57043
rect 3338 57031 3344 57043
rect 3338 57003 5822 57031
rect 3338 56991 3344 57003
rect 1939 56960 1997 56966
rect 1939 56957 1951 56960
rect 266 56929 1951 56957
rect 266 56917 272 56929
rect 1939 56926 1951 56929
rect 1985 56926 1997 56960
rect 1939 56920 1997 56926
rect 2803 56960 2861 56966
rect 2803 56926 2815 56960
rect 2849 56926 2861 56960
rect 2803 56920 2861 56926
rect 4912 56917 4918 56969
rect 4970 56957 4976 56969
rect 5794 56966 5822 57003
rect 9616 56991 9622 57043
rect 9674 57031 9680 57043
rect 9907 57034 9965 57040
rect 9907 57031 9919 57034
rect 9674 57003 9919 57031
rect 9674 56991 9680 57003
rect 9907 57000 9919 57003
rect 9953 57000 9965 57034
rect 9907 56994 9965 57000
rect 11248 56991 11254 57043
rect 11306 57031 11312 57043
rect 14035 57034 14093 57040
rect 11306 57003 11486 57031
rect 11306 56991 11312 57003
rect 5299 56960 5357 56966
rect 5299 56957 5311 56960
rect 4970 56929 5311 56957
rect 4970 56917 4976 56929
rect 5299 56926 5311 56929
rect 5345 56926 5357 56960
rect 5299 56920 5357 56926
rect 5779 56960 5837 56966
rect 5779 56926 5791 56960
rect 5825 56926 5837 56960
rect 5779 56920 5837 56926
rect 6448 56917 6454 56969
rect 6506 56957 6512 56969
rect 7411 56960 7469 56966
rect 7411 56957 7423 56960
rect 6506 56929 7423 56957
rect 6506 56917 6512 56929
rect 7411 56926 7423 56929
rect 7457 56926 7469 56960
rect 8080 56957 8086 56969
rect 8041 56929 8086 56957
rect 7411 56920 7469 56926
rect 8080 56917 8086 56929
rect 8138 56917 8144 56969
rect 11458 56966 11486 57003
rect 14035 57000 14047 57034
rect 14081 57031 14093 57034
rect 16432 57031 16438 57043
rect 14081 57003 16438 57031
rect 14081 57000 14093 57003
rect 14035 56994 14093 57000
rect 16432 56991 16438 57003
rect 16490 56991 16496 57043
rect 29104 56991 29110 57043
rect 29162 57031 29168 57043
rect 32563 57034 32621 57040
rect 32563 57031 32575 57034
rect 29162 57003 32575 57031
rect 29162 56991 29168 57003
rect 32563 57000 32575 57003
rect 32609 57000 32621 57034
rect 32563 56994 32621 57000
rect 11443 56960 11501 56966
rect 11443 56926 11455 56960
rect 11489 56926 11501 56960
rect 11443 56920 11501 56926
rect 12784 56917 12790 56969
rect 12842 56957 12848 56969
rect 13171 56960 13229 56966
rect 13171 56957 13183 56960
rect 12842 56929 13183 56957
rect 12842 56917 12848 56929
rect 13171 56926 13183 56929
rect 13217 56926 13229 56960
rect 13171 56920 13229 56926
rect 14416 56917 14422 56969
rect 14474 56957 14480 56969
rect 15091 56960 15149 56966
rect 15091 56957 15103 56960
rect 14474 56929 15103 56957
rect 14474 56917 14480 56929
rect 15091 56926 15103 56929
rect 15137 56926 15149 56960
rect 15091 56920 15149 56926
rect 15952 56917 15958 56969
rect 16010 56957 16016 56969
rect 16339 56960 16397 56966
rect 16339 56957 16351 56960
rect 16010 56929 16351 56957
rect 16010 56917 16016 56929
rect 16339 56926 16351 56929
rect 16385 56926 16397 56960
rect 16339 56920 16397 56926
rect 17488 56917 17494 56969
rect 17546 56957 17552 56969
rect 18163 56960 18221 56966
rect 18163 56957 18175 56960
rect 17546 56929 18175 56957
rect 17546 56917 17552 56929
rect 18163 56926 18175 56929
rect 18209 56926 18221 56960
rect 18163 56920 18221 56926
rect 19120 56917 19126 56969
rect 19178 56957 19184 56969
rect 19507 56960 19565 56966
rect 19507 56957 19519 56960
rect 19178 56929 19519 56957
rect 19178 56917 19184 56929
rect 19507 56926 19519 56929
rect 19553 56926 19565 56960
rect 19507 56920 19565 56926
rect 20656 56917 20662 56969
rect 20714 56957 20720 56969
rect 21043 56960 21101 56966
rect 21043 56957 21055 56960
rect 20714 56929 21055 56957
rect 20714 56917 20720 56929
rect 21043 56926 21055 56929
rect 21089 56926 21101 56960
rect 21043 56920 21101 56926
rect 22003 56960 22061 56966
rect 22003 56926 22015 56960
rect 22049 56957 22061 56960
rect 22288 56957 22294 56969
rect 22049 56929 22294 56957
rect 22049 56926 22061 56929
rect 22003 56920 22061 56926
rect 22288 56917 22294 56929
rect 22346 56917 22352 56969
rect 23824 56917 23830 56969
rect 23882 56957 23888 56969
rect 24211 56960 24269 56966
rect 24211 56957 24223 56960
rect 23882 56929 24223 56957
rect 23882 56917 23888 56929
rect 24211 56926 24223 56929
rect 24257 56926 24269 56960
rect 24211 56920 24269 56926
rect 25456 56917 25462 56969
rect 25514 56957 25520 56969
rect 25939 56960 25997 56966
rect 25939 56957 25951 56960
rect 25514 56929 25951 56957
rect 25514 56917 25520 56929
rect 25939 56926 25951 56929
rect 25985 56926 25997 56960
rect 25939 56920 25997 56926
rect 26992 56917 26998 56969
rect 27050 56957 27056 56969
rect 27379 56960 27437 56966
rect 27379 56957 27391 56960
rect 27050 56929 27391 56957
rect 27050 56917 27056 56929
rect 27379 56926 27391 56929
rect 27425 56926 27437 56960
rect 28624 56957 28630 56969
rect 28585 56929 28630 56957
rect 27379 56920 27437 56926
rect 28624 56917 28630 56929
rect 28682 56917 28688 56969
rect 30256 56957 30262 56969
rect 30217 56929 30262 56957
rect 30256 56917 30262 56929
rect 30314 56917 30320 56969
rect 31696 56957 31702 56969
rect 31657 56929 31702 56957
rect 31696 56917 31702 56929
rect 31754 56917 31760 56969
rect 33328 56917 33334 56969
rect 33386 56957 33392 56969
rect 34291 56960 34349 56966
rect 34291 56957 34303 56960
rect 33386 56929 34303 56957
rect 33386 56917 33392 56929
rect 34291 56926 34303 56929
rect 34337 56926 34349 56960
rect 34864 56957 34870 56969
rect 34825 56929 34870 56957
rect 34291 56920 34349 56926
rect 34864 56917 34870 56929
rect 34922 56917 34928 56969
rect 38032 56957 38038 56969
rect 37993 56929 38038 56957
rect 38032 56917 38038 56929
rect 38090 56917 38096 56969
rect 41200 56917 41206 56969
rect 41258 56957 41264 56969
rect 41971 56960 42029 56966
rect 41971 56957 41983 56960
rect 41258 56929 41983 56957
rect 41258 56917 41264 56929
rect 41971 56926 41983 56929
rect 42017 56926 42029 56960
rect 41971 56920 42029 56926
rect 44368 56917 44374 56969
rect 44426 56957 44432 56969
rect 44659 56960 44717 56966
rect 44659 56957 44671 56960
rect 44426 56929 44671 56957
rect 44426 56917 44432 56929
rect 44659 56926 44671 56929
rect 44705 56926 44717 56960
rect 47536 56957 47542 56969
rect 47497 56929 47542 56957
rect 44659 56920 44717 56926
rect 47536 56917 47542 56929
rect 47594 56917 47600 56969
rect 53872 56957 53878 56969
rect 53833 56929 53878 56957
rect 53872 56917 53878 56929
rect 53930 56917 53936 56969
rect 1747 56886 1805 56892
rect 1747 56852 1759 56886
rect 1793 56852 1805 56886
rect 1747 56846 1805 56852
rect 2611 56886 2669 56892
rect 2611 56852 2623 56886
rect 2657 56883 2669 56886
rect 3664 56883 3670 56895
rect 2657 56855 3670 56883
rect 2657 56852 2669 56855
rect 2611 56846 2669 56852
rect 1762 56809 1790 56846
rect 3664 56843 3670 56855
rect 3722 56843 3728 56895
rect 5104 56883 5110 56895
rect 5065 56855 5110 56883
rect 5104 56843 5110 56855
rect 5162 56843 5168 56895
rect 7219 56886 7277 56892
rect 7219 56852 7231 56886
rect 7265 56883 7277 56886
rect 8272 56883 8278 56895
rect 7265 56855 8278 56883
rect 7265 56852 7277 56855
rect 7219 56846 7277 56852
rect 8272 56843 8278 56855
rect 8330 56843 8336 56895
rect 11248 56883 11254 56895
rect 11209 56855 11254 56883
rect 11248 56843 11254 56855
rect 11306 56843 11312 56895
rect 12976 56883 12982 56895
rect 12937 56855 12982 56883
rect 12976 56843 12982 56855
rect 13034 56843 13040 56895
rect 13648 56843 13654 56895
rect 13706 56883 13712 56895
rect 13939 56886 13997 56892
rect 13939 56883 13951 56886
rect 13706 56855 13951 56883
rect 13706 56843 13712 56855
rect 13939 56852 13951 56855
rect 13985 56852 13997 56886
rect 16144 56883 16150 56895
rect 16105 56855 16150 56883
rect 13939 56846 13997 56852
rect 16144 56843 16150 56855
rect 16202 56843 16208 56895
rect 17968 56883 17974 56895
rect 17929 56855 17974 56883
rect 17968 56843 17974 56855
rect 18026 56843 18032 56895
rect 19312 56883 19318 56895
rect 19273 56855 19318 56883
rect 19312 56843 19318 56855
rect 19370 56843 19376 56895
rect 20851 56886 20909 56892
rect 20851 56852 20863 56886
rect 20897 56852 20909 56886
rect 24016 56883 24022 56895
rect 23977 56855 24022 56883
rect 20851 56846 20909 56852
rect 3568 56809 3574 56821
rect 1762 56781 3574 56809
rect 3568 56769 3574 56781
rect 3626 56769 3632 56821
rect 10768 56769 10774 56821
rect 10826 56809 10832 56821
rect 20866 56809 20894 56846
rect 24016 56843 24022 56855
rect 24074 56843 24080 56895
rect 27184 56883 27190 56895
rect 27145 56855 27190 56883
rect 27184 56843 27190 56855
rect 27242 56843 27248 56895
rect 29968 56843 29974 56895
rect 30026 56883 30032 56895
rect 30067 56886 30125 56892
rect 30067 56883 30079 56886
rect 30026 56855 30079 56883
rect 30026 56843 30032 56855
rect 30067 56852 30079 56855
rect 30113 56852 30125 56886
rect 30067 56846 30125 56852
rect 32659 56886 32717 56892
rect 32659 56852 32671 56886
rect 32705 56852 32717 56886
rect 34096 56883 34102 56895
rect 34057 56855 34102 56883
rect 32659 56846 32717 56852
rect 10826 56781 20894 56809
rect 32674 56809 32702 56846
rect 34096 56843 34102 56855
rect 34154 56843 34160 56895
rect 36496 56843 36502 56895
rect 36554 56883 36560 56895
rect 36979 56886 37037 56892
rect 36979 56883 36991 56886
rect 36554 56855 36991 56883
rect 36554 56843 36560 56855
rect 36979 56852 36991 56855
rect 37025 56852 37037 56886
rect 36979 56846 37037 56852
rect 39664 56843 39670 56895
rect 39722 56883 39728 56895
rect 40051 56886 40109 56892
rect 40051 56883 40063 56886
rect 39722 56855 40063 56883
rect 39722 56843 39728 56855
rect 40051 56852 40063 56855
rect 40097 56852 40109 56886
rect 40051 56846 40109 56852
rect 40531 56886 40589 56892
rect 40531 56852 40543 56886
rect 40577 56883 40589 56886
rect 40624 56883 40630 56895
rect 40577 56855 40630 56883
rect 40577 56852 40589 56855
rect 40531 56846 40589 56852
rect 40624 56843 40630 56855
rect 40682 56883 40688 56895
rect 40723 56886 40781 56892
rect 40723 56883 40735 56886
rect 40682 56855 40735 56883
rect 40682 56843 40688 56855
rect 40723 56852 40735 56855
rect 40769 56852 40781 56886
rect 40723 56846 40781 56852
rect 42832 56843 42838 56895
rect 42890 56883 42896 56895
rect 43219 56886 43277 56892
rect 43219 56883 43231 56886
rect 42890 56855 43231 56883
rect 42890 56843 42896 56855
rect 43219 56852 43231 56855
rect 43265 56852 43277 56886
rect 43219 56846 43277 56852
rect 46096 56843 46102 56895
rect 46154 56883 46160 56895
rect 46291 56886 46349 56892
rect 46291 56883 46303 56886
rect 46154 56855 46303 56883
rect 46154 56843 46160 56855
rect 46291 56852 46303 56855
rect 46337 56852 46349 56886
rect 46291 56846 46349 56852
rect 48979 56886 49037 56892
rect 48979 56852 48991 56886
rect 49025 56883 49037 56886
rect 49072 56883 49078 56895
rect 49025 56855 49078 56883
rect 49025 56852 49037 56855
rect 48979 56846 49037 56852
rect 49072 56843 49078 56855
rect 49130 56843 49136 56895
rect 50704 56843 50710 56895
rect 50762 56883 50768 56895
rect 51091 56886 51149 56892
rect 51091 56883 51103 56886
rect 50762 56855 51103 56883
rect 50762 56843 50768 56855
rect 51091 56852 51103 56855
rect 51137 56852 51149 56886
rect 51091 56846 51149 56852
rect 52240 56843 52246 56895
rect 52298 56883 52304 56895
rect 53107 56886 53165 56892
rect 53107 56883 53119 56886
rect 52298 56855 53119 56883
rect 52298 56843 52304 56855
rect 53107 56852 53119 56855
rect 53153 56852 53165 56886
rect 53107 56846 53165 56852
rect 55408 56843 55414 56895
rect 55466 56883 55472 56895
rect 55795 56886 55853 56892
rect 55795 56883 55807 56886
rect 55466 56855 55807 56883
rect 55466 56843 55472 56855
rect 55795 56852 55807 56855
rect 55841 56852 55853 56886
rect 57040 56883 57046 56895
rect 57001 56855 57046 56883
rect 55795 56846 55853 56852
rect 57040 56843 57046 56855
rect 57098 56843 57104 56895
rect 40336 56809 40342 56821
rect 32674 56781 40342 56809
rect 10826 56769 10832 56781
rect 40336 56769 40342 56781
rect 40394 56769 40400 56821
rect 9808 56735 9814 56747
rect 9769 56707 9814 56735
rect 9808 56695 9814 56707
rect 9866 56695 9872 56747
rect 13648 56735 13654 56747
rect 13609 56707 13654 56735
rect 13648 56695 13654 56707
rect 13706 56695 13712 56747
rect 36688 56735 36694 56747
rect 36649 56707 36694 56735
rect 36688 56695 36694 56707
rect 36746 56695 36752 56747
rect 39760 56735 39766 56747
rect 39721 56707 39766 56735
rect 39760 56695 39766 56707
rect 39818 56695 39824 56747
rect 40816 56735 40822 56747
rect 40777 56707 40822 56735
rect 40816 56695 40822 56707
rect 40874 56695 40880 56747
rect 42928 56735 42934 56747
rect 42889 56707 42934 56735
rect 42928 56695 42934 56707
rect 42986 56695 42992 56747
rect 46003 56738 46061 56744
rect 46003 56704 46015 56738
rect 46049 56735 46061 56738
rect 46096 56735 46102 56747
rect 46049 56707 46102 56735
rect 46049 56704 46061 56707
rect 46003 56698 46061 56704
rect 46096 56695 46102 56707
rect 46154 56695 46160 56747
rect 48688 56735 48694 56747
rect 48649 56707 48694 56735
rect 48688 56695 48694 56707
rect 48746 56695 48752 56747
rect 50800 56735 50806 56747
rect 50761 56707 50806 56735
rect 50800 56695 50806 56707
rect 50858 56695 50864 56747
rect 52816 56735 52822 56747
rect 52777 56707 52822 56735
rect 52816 56695 52822 56707
rect 52874 56695 52880 56747
rect 55408 56695 55414 56747
rect 55466 56735 55472 56747
rect 55507 56738 55565 56744
rect 55507 56735 55519 56738
rect 55466 56707 55519 56735
rect 55466 56695 55472 56707
rect 55507 56704 55519 56707
rect 55553 56704 55565 56738
rect 56752 56735 56758 56747
rect 56713 56707 56758 56735
rect 55507 56698 55565 56704
rect 56752 56695 56758 56707
rect 56810 56695 56816 56747
rect 1152 56636 58848 56658
rect 1152 56584 19654 56636
rect 19706 56584 19718 56636
rect 19770 56584 19782 56636
rect 19834 56584 19846 56636
rect 19898 56584 50374 56636
rect 50426 56584 50438 56636
rect 50490 56584 50502 56636
rect 50554 56584 50566 56636
rect 50618 56584 58848 56636
rect 1152 56562 58848 56584
rect 688 56473 694 56525
rect 746 56513 752 56525
rect 1651 56516 1709 56522
rect 1651 56513 1663 56516
rect 746 56485 1663 56513
rect 746 56473 752 56485
rect 1651 56482 1663 56485
rect 1697 56482 1709 56516
rect 1651 56476 1709 56482
rect 2224 56473 2230 56525
rect 2282 56513 2288 56525
rect 2419 56516 2477 56522
rect 2419 56513 2431 56516
rect 2282 56485 2431 56513
rect 2282 56473 2288 56485
rect 2419 56482 2431 56485
rect 2465 56482 2477 56516
rect 2419 56476 2477 56482
rect 2800 56473 2806 56525
rect 2858 56513 2864 56525
rect 3187 56516 3245 56522
rect 3187 56513 3199 56516
rect 2858 56485 3199 56513
rect 2858 56473 2864 56485
rect 3187 56482 3199 56485
rect 3233 56482 3245 56516
rect 3187 56476 3245 56482
rect 3856 56473 3862 56525
rect 3914 56513 3920 56525
rect 4435 56516 4493 56522
rect 4435 56513 4447 56516
rect 3914 56485 4447 56513
rect 3914 56473 3920 56485
rect 4435 56482 4447 56485
rect 4481 56482 4493 56516
rect 4435 56476 4493 56482
rect 5392 56473 5398 56525
rect 5450 56513 5456 56525
rect 5491 56516 5549 56522
rect 5491 56513 5503 56516
rect 5450 56485 5503 56513
rect 5450 56473 5456 56485
rect 5491 56482 5503 56485
rect 5537 56482 5549 56516
rect 5491 56476 5549 56482
rect 5968 56473 5974 56525
rect 6026 56513 6032 56525
rect 6259 56516 6317 56522
rect 6259 56513 6271 56516
rect 6026 56485 6271 56513
rect 6026 56473 6032 56485
rect 6259 56482 6271 56485
rect 6305 56482 6317 56516
rect 6259 56476 6317 56482
rect 7024 56473 7030 56525
rect 7082 56513 7088 56525
rect 7123 56516 7181 56522
rect 7123 56513 7135 56516
rect 7082 56485 7135 56513
rect 7082 56473 7088 56485
rect 7123 56482 7135 56485
rect 7169 56482 7181 56516
rect 8560 56513 8566 56525
rect 8521 56485 8566 56513
rect 7123 56476 7181 56482
rect 8560 56473 8566 56485
rect 8618 56473 8624 56525
rect 10192 56473 10198 56525
rect 10250 56513 10256 56525
rect 10291 56516 10349 56522
rect 10291 56513 10303 56516
rect 10250 56485 10303 56513
rect 10250 56473 10256 56485
rect 10291 56482 10303 56485
rect 10337 56482 10349 56516
rect 10291 56476 10349 56482
rect 10672 56473 10678 56525
rect 10730 56513 10736 56525
rect 11059 56516 11117 56522
rect 11059 56513 11071 56516
rect 10730 56485 11071 56513
rect 10730 56473 10736 56485
rect 11059 56482 11071 56485
rect 11105 56482 11117 56516
rect 11059 56476 11117 56482
rect 11728 56473 11734 56525
rect 11786 56513 11792 56525
rect 11827 56516 11885 56522
rect 11827 56513 11839 56516
rect 11786 56485 11839 56513
rect 11786 56473 11792 56485
rect 11827 56482 11839 56485
rect 11873 56482 11885 56516
rect 11827 56476 11885 56482
rect 12304 56473 12310 56525
rect 12362 56513 12368 56525
rect 12595 56516 12653 56522
rect 12595 56513 12607 56516
rect 12362 56485 12607 56513
rect 12362 56473 12368 56485
rect 12595 56482 12607 56485
rect 12641 56482 12653 56516
rect 12595 56476 12653 56482
rect 13360 56473 13366 56525
rect 13418 56513 13424 56525
rect 13555 56516 13613 56522
rect 13555 56513 13567 56516
rect 13418 56485 13567 56513
rect 13418 56473 13424 56485
rect 13555 56482 13567 56485
rect 13601 56482 13613 56516
rect 13555 56476 13613 56482
rect 14896 56473 14902 56525
rect 14954 56513 14960 56525
rect 14995 56516 15053 56522
rect 14995 56513 15007 56516
rect 14954 56485 15007 56513
rect 14954 56473 14960 56485
rect 14995 56482 15007 56485
rect 15041 56482 15053 56516
rect 14995 56476 15053 56482
rect 17008 56473 17014 56525
rect 17066 56513 17072 56525
rect 17107 56516 17165 56522
rect 17107 56513 17119 56516
rect 17066 56485 17119 56513
rect 17066 56473 17072 56485
rect 17107 56482 17119 56485
rect 17153 56482 17165 56516
rect 17107 56476 17165 56482
rect 18064 56473 18070 56525
rect 18122 56513 18128 56525
rect 18163 56516 18221 56522
rect 18163 56513 18175 56516
rect 18122 56485 18175 56513
rect 18122 56473 18128 56485
rect 18163 56482 18175 56485
rect 18209 56482 18221 56516
rect 18163 56476 18221 56482
rect 18544 56473 18550 56525
rect 18602 56513 18608 56525
rect 18931 56516 18989 56522
rect 18931 56513 18943 56516
rect 18602 56485 18943 56513
rect 18602 56473 18608 56485
rect 18931 56482 18943 56485
rect 18977 56482 18989 56516
rect 18931 56476 18989 56482
rect 19984 56473 19990 56525
rect 20042 56513 20048 56525
rect 20275 56516 20333 56522
rect 20275 56513 20287 56516
rect 20042 56485 20287 56513
rect 20042 56473 20048 56485
rect 20275 56482 20287 56485
rect 20321 56482 20333 56516
rect 20275 56476 20333 56482
rect 21232 56473 21238 56525
rect 21290 56513 21296 56525
rect 21331 56516 21389 56522
rect 21331 56513 21343 56516
rect 21290 56485 21343 56513
rect 21290 56473 21296 56485
rect 21331 56482 21343 56485
rect 21377 56482 21389 56516
rect 21331 56476 21389 56482
rect 21712 56473 21718 56525
rect 21770 56513 21776 56525
rect 22099 56516 22157 56522
rect 22099 56513 22111 56516
rect 21770 56485 22111 56513
rect 21770 56473 21776 56485
rect 22099 56482 22111 56485
rect 22145 56482 22157 56516
rect 22099 56476 22157 56482
rect 22768 56473 22774 56525
rect 22826 56513 22832 56525
rect 22867 56516 22925 56522
rect 22867 56513 22879 56516
rect 22826 56485 22879 56513
rect 22826 56473 22832 56485
rect 22867 56482 22879 56485
rect 22913 56482 22925 56516
rect 22867 56476 22925 56482
rect 24307 56516 24365 56522
rect 24307 56482 24319 56516
rect 24353 56513 24365 56516
rect 24400 56513 24406 56525
rect 24353 56485 24406 56513
rect 24353 56482 24365 56485
rect 24307 56476 24365 56482
rect 24400 56473 24406 56485
rect 24458 56473 24464 56525
rect 25936 56473 25942 56525
rect 25994 56513 26000 56525
rect 26035 56516 26093 56522
rect 26035 56513 26047 56516
rect 25994 56485 26047 56513
rect 25994 56473 26000 56485
rect 26035 56482 26047 56485
rect 26081 56482 26093 56516
rect 26035 56476 26093 56482
rect 26512 56473 26518 56525
rect 26570 56513 26576 56525
rect 26899 56516 26957 56522
rect 26899 56513 26911 56516
rect 26570 56485 26911 56513
rect 26570 56473 26576 56485
rect 26899 56482 26911 56485
rect 26945 56482 26957 56516
rect 26899 56476 26957 56482
rect 27568 56473 27574 56525
rect 27626 56513 27632 56525
rect 27763 56516 27821 56522
rect 27763 56513 27775 56516
rect 27626 56485 27775 56513
rect 27626 56473 27632 56485
rect 27763 56482 27775 56485
rect 27809 56482 27821 56516
rect 27763 56476 27821 56482
rect 28048 56473 28054 56525
rect 28106 56513 28112 56525
rect 28531 56516 28589 56522
rect 28531 56513 28543 56516
rect 28106 56485 28543 56513
rect 28106 56473 28112 56485
rect 28531 56482 28543 56485
rect 28577 56482 28589 56516
rect 29680 56513 29686 56525
rect 29641 56485 29686 56513
rect 28531 56476 28589 56482
rect 29680 56473 29686 56485
rect 29738 56473 29744 56525
rect 30640 56473 30646 56525
rect 30698 56513 30704 56525
rect 30835 56516 30893 56522
rect 30835 56513 30847 56516
rect 30698 56485 30847 56513
rect 30698 56473 30704 56485
rect 30835 56482 30847 56485
rect 30881 56482 30893 56516
rect 30835 56476 30893 56482
rect 31216 56473 31222 56525
rect 31274 56513 31280 56525
rect 31603 56516 31661 56522
rect 31603 56513 31615 56516
rect 31274 56485 31615 56513
rect 31274 56473 31280 56485
rect 31603 56482 31615 56485
rect 31649 56482 31661 56516
rect 31603 56476 31661 56482
rect 32272 56473 32278 56525
rect 32330 56513 32336 56525
rect 32371 56516 32429 56522
rect 32371 56513 32383 56516
rect 32330 56485 32383 56513
rect 32330 56473 32336 56485
rect 32371 56482 32383 56485
rect 32417 56482 32429 56516
rect 32371 56476 32429 56482
rect 33808 56473 33814 56525
rect 33866 56513 33872 56525
rect 33907 56516 33965 56522
rect 33907 56513 33919 56516
rect 33866 56485 33919 56513
rect 33866 56473 33872 56485
rect 33907 56482 33919 56485
rect 33953 56482 33965 56516
rect 33907 56476 33965 56482
rect 34576 56473 34582 56525
rect 34634 56513 34640 56525
rect 34771 56516 34829 56522
rect 34771 56513 34783 56516
rect 34634 56485 34783 56513
rect 34634 56473 34640 56485
rect 34771 56482 34783 56485
rect 34817 56482 34829 56516
rect 34771 56476 34829 56482
rect 36016 56473 36022 56525
rect 36074 56513 36080 56525
rect 36979 56516 37037 56522
rect 36979 56513 36991 56516
rect 36074 56485 36991 56513
rect 36074 56473 36080 56485
rect 36979 56482 36991 56485
rect 37025 56482 37037 56516
rect 36979 56476 37037 56482
rect 37552 56473 37558 56525
rect 37610 56513 37616 56525
rect 37651 56516 37709 56522
rect 37651 56513 37663 56516
rect 37610 56485 37663 56513
rect 37610 56473 37616 56485
rect 37651 56482 37663 56485
rect 37697 56482 37709 56516
rect 37651 56476 37709 56482
rect 38608 56473 38614 56525
rect 38666 56513 38672 56525
rect 38803 56516 38861 56522
rect 38803 56513 38815 56516
rect 38666 56485 38815 56513
rect 38666 56473 38672 56485
rect 38803 56482 38815 56485
rect 38849 56482 38861 56516
rect 40144 56513 40150 56525
rect 40105 56485 40150 56513
rect 38803 56476 38861 56482
rect 40144 56473 40150 56485
rect 40202 56473 40208 56525
rect 41776 56473 41782 56525
rect 41834 56513 41840 56525
rect 41875 56516 41933 56522
rect 41875 56513 41887 56516
rect 41834 56485 41887 56513
rect 41834 56473 41840 56485
rect 41875 56482 41887 56485
rect 41921 56482 41933 56516
rect 41875 56476 41933 56482
rect 42256 56473 42262 56525
rect 42314 56513 42320 56525
rect 42739 56516 42797 56522
rect 42739 56513 42751 56516
rect 42314 56485 42751 56513
rect 42314 56473 42320 56485
rect 42739 56482 42751 56485
rect 42785 56482 42797 56516
rect 42739 56476 42797 56482
rect 43312 56473 43318 56525
rect 43370 56513 43376 56525
rect 43507 56516 43565 56522
rect 43507 56513 43519 56516
rect 43370 56485 43519 56513
rect 43370 56473 43376 56485
rect 43507 56482 43519 56485
rect 43553 56482 43565 56516
rect 43507 56476 43565 56482
rect 43888 56473 43894 56525
rect 43946 56513 43952 56525
rect 44275 56516 44333 56522
rect 44275 56513 44287 56516
rect 43946 56485 44287 56513
rect 43946 56473 43952 56485
rect 44275 56482 44287 56485
rect 44321 56482 44333 56516
rect 44275 56476 44333 56482
rect 44944 56473 44950 56525
rect 45002 56513 45008 56525
rect 45139 56516 45197 56522
rect 45139 56513 45151 56516
rect 45002 56485 45151 56513
rect 45002 56473 45008 56485
rect 45139 56482 45151 56485
rect 45185 56482 45197 56516
rect 45139 56476 45197 56482
rect 46480 56473 46486 56525
rect 46538 56513 46544 56525
rect 46675 56516 46733 56522
rect 46675 56513 46687 56516
rect 46538 56485 46687 56513
rect 46538 56473 46544 56485
rect 46675 56482 46687 56485
rect 46721 56482 46733 56516
rect 46675 56476 46733 56482
rect 48016 56473 48022 56525
rect 48074 56513 48080 56525
rect 48115 56516 48173 56522
rect 48115 56513 48127 56516
rect 48074 56485 48127 56513
rect 48074 56473 48080 56485
rect 48115 56482 48127 56485
rect 48161 56482 48173 56516
rect 48115 56476 48173 56482
rect 49648 56473 49654 56525
rect 49706 56513 49712 56525
rect 49747 56516 49805 56522
rect 49747 56513 49759 56516
rect 49706 56485 49759 56513
rect 49706 56473 49712 56485
rect 49747 56482 49759 56485
rect 49793 56482 49805 56516
rect 49747 56476 49805 56482
rect 50128 56473 50134 56525
rect 50186 56513 50192 56525
rect 50515 56516 50573 56522
rect 50515 56513 50527 56516
rect 50186 56485 50527 56513
rect 50186 56473 50192 56485
rect 50515 56482 50527 56485
rect 50561 56482 50573 56516
rect 50515 56476 50573 56482
rect 52912 56473 52918 56525
rect 52970 56513 52976 56525
rect 53011 56516 53069 56522
rect 53011 56513 53023 56516
rect 52970 56485 53023 56513
rect 52970 56473 52976 56485
rect 53011 56482 53023 56485
rect 53057 56482 53069 56516
rect 53011 56476 53069 56482
rect 53296 56473 53302 56525
rect 53354 56513 53360 56525
rect 53779 56516 53837 56522
rect 53779 56513 53791 56516
rect 53354 56485 53791 56513
rect 53354 56473 53360 56485
rect 53779 56482 53791 56485
rect 53825 56482 53837 56516
rect 53779 56476 53837 56482
rect 54352 56473 54358 56525
rect 54410 56513 54416 56525
rect 54451 56516 54509 56522
rect 54451 56513 54463 56516
rect 54410 56485 54463 56513
rect 54410 56473 54416 56485
rect 54451 56482 54463 56485
rect 54497 56482 54509 56516
rect 54451 56476 54509 56482
rect 54928 56473 54934 56525
rect 54986 56513 54992 56525
rect 55315 56516 55373 56522
rect 55315 56513 55327 56516
rect 54986 56485 55327 56513
rect 54986 56473 54992 56485
rect 55315 56482 55327 56485
rect 55361 56482 55373 56516
rect 55315 56476 55373 56482
rect 55984 56473 55990 56525
rect 56042 56513 56048 56525
rect 56083 56516 56141 56522
rect 56083 56513 56095 56516
rect 56042 56485 56095 56513
rect 56042 56473 56048 56485
rect 56083 56482 56095 56485
rect 56129 56482 56141 56516
rect 56083 56476 56141 56482
rect 26608 56399 26614 56451
rect 26666 56439 26672 56451
rect 56752 56439 56758 56451
rect 26666 56411 56758 56439
rect 26666 56399 26672 56411
rect 56752 56399 56758 56411
rect 56810 56399 56816 56451
rect 4531 56368 4589 56374
rect 4531 56334 4543 56368
rect 4577 56365 4589 56368
rect 11440 56365 11446 56377
rect 4577 56337 11446 56365
rect 4577 56334 4589 56337
rect 4531 56328 4589 56334
rect 11440 56325 11446 56337
rect 11498 56325 11504 56377
rect 12208 56325 12214 56377
rect 12266 56365 12272 56377
rect 15475 56368 15533 56374
rect 15475 56365 15487 56368
rect 12266 56337 15487 56365
rect 12266 56325 12272 56337
rect 15475 56334 15487 56337
rect 15521 56365 15533 56368
rect 15763 56368 15821 56374
rect 15763 56365 15775 56368
rect 15521 56337 15775 56365
rect 15521 56334 15533 56337
rect 15475 56328 15533 56334
rect 15763 56334 15775 56337
rect 15809 56334 15821 56368
rect 15763 56328 15821 56334
rect 19027 56368 19085 56374
rect 19027 56334 19039 56368
rect 19073 56365 19085 56368
rect 28720 56365 28726 56377
rect 19073 56337 28726 56365
rect 19073 56334 19085 56337
rect 19027 56328 19085 56334
rect 28720 56325 28726 56337
rect 28778 56325 28784 56377
rect 43888 56325 43894 56377
rect 43946 56365 43952 56377
rect 43946 56337 53294 56365
rect 43946 56325 43952 56337
rect 1747 56294 1805 56300
rect 1747 56260 1759 56294
rect 1793 56291 1805 56294
rect 2704 56291 2710 56303
rect 1793 56263 2710 56291
rect 1793 56260 1805 56263
rect 1747 56254 1805 56260
rect 2704 56251 2710 56263
rect 2762 56251 2768 56303
rect 2800 56251 2806 56303
rect 2858 56291 2864 56303
rect 24403 56294 24461 56300
rect 24403 56291 24415 56294
rect 2858 56263 24415 56291
rect 2858 56251 2864 56263
rect 24403 56260 24415 56263
rect 24449 56260 24461 56294
rect 24403 56254 24461 56260
rect 42544 56251 42550 56303
rect 42602 56291 42608 56303
rect 52627 56294 52685 56300
rect 52627 56291 52639 56294
rect 42602 56263 52639 56291
rect 42602 56251 42608 56263
rect 52627 56260 52639 56263
rect 52673 56291 52685 56294
rect 52915 56294 52973 56300
rect 52915 56291 52927 56294
rect 52673 56263 52927 56291
rect 52673 56260 52685 56263
rect 52627 56254 52685 56260
rect 52915 56260 52927 56263
rect 52961 56260 52973 56294
rect 53266 56291 53294 56337
rect 55699 56294 55757 56300
rect 55699 56291 55711 56294
rect 53266 56263 55711 56291
rect 52915 56254 52973 56260
rect 55699 56260 55711 56263
rect 55745 56291 55757 56294
rect 55987 56294 56045 56300
rect 55987 56291 55999 56294
rect 55745 56263 55999 56291
rect 55745 56260 55757 56263
rect 55699 56254 55757 56260
rect 55987 56260 55999 56263
rect 56033 56260 56045 56294
rect 55987 56254 56045 56260
rect 57811 56294 57869 56300
rect 57811 56260 57823 56294
rect 57857 56291 57869 56294
rect 58576 56291 58582 56303
rect 57857 56263 58582 56291
rect 57857 56260 57869 56263
rect 57811 56254 57869 56260
rect 58576 56251 58582 56263
rect 58634 56251 58640 56303
rect 2515 56220 2573 56226
rect 2515 56186 2527 56220
rect 2561 56217 2573 56220
rect 2608 56217 2614 56229
rect 2561 56189 2614 56217
rect 2561 56186 2573 56189
rect 2515 56180 2573 56186
rect 2608 56177 2614 56189
rect 2666 56177 2672 56229
rect 2995 56220 3053 56226
rect 2995 56186 3007 56220
rect 3041 56217 3053 56220
rect 3280 56217 3286 56229
rect 3041 56189 3286 56217
rect 3041 56186 3053 56189
rect 2995 56180 3053 56186
rect 3280 56177 3286 56189
rect 3338 56177 3344 56229
rect 5584 56217 5590 56229
rect 5545 56189 5590 56217
rect 5584 56177 5590 56189
rect 5642 56177 5648 56229
rect 5968 56217 5974 56229
rect 5929 56189 5974 56217
rect 5968 56177 5974 56189
rect 6026 56217 6032 56229
rect 6355 56220 6413 56226
rect 6355 56217 6367 56220
rect 6026 56189 6367 56217
rect 6026 56177 6032 56189
rect 6355 56186 6367 56189
rect 6401 56186 6413 56220
rect 6355 56180 6413 56186
rect 7216 56177 7222 56229
rect 7274 56217 7280 56229
rect 8176 56217 8182 56229
rect 7274 56189 7319 56217
rect 8137 56189 8182 56217
rect 7274 56177 7280 56189
rect 8176 56177 8182 56189
rect 8234 56217 8240 56229
rect 8467 56220 8525 56226
rect 8467 56217 8479 56220
rect 8234 56189 8479 56217
rect 8234 56177 8240 56189
rect 8467 56186 8479 56189
rect 8513 56186 8525 56220
rect 10096 56217 10102 56229
rect 10057 56189 10102 56217
rect 8467 56180 8525 56186
rect 10096 56177 10102 56189
rect 10154 56217 10160 56229
rect 10387 56220 10445 56226
rect 10387 56217 10399 56220
rect 10154 56189 10399 56217
rect 10154 56177 10160 56189
rect 10387 56186 10399 56189
rect 10433 56186 10445 56220
rect 11152 56217 11158 56229
rect 11113 56189 11158 56217
rect 10387 56180 10445 56186
rect 11152 56177 11158 56189
rect 11210 56177 11216 56229
rect 11920 56217 11926 56229
rect 11881 56189 11926 56217
rect 11920 56177 11926 56189
rect 11978 56177 11984 56229
rect 12688 56217 12694 56229
rect 12649 56189 12694 56217
rect 12688 56177 12694 56189
rect 12746 56177 12752 56229
rect 13264 56217 13270 56229
rect 13225 56189 13270 56217
rect 13264 56177 13270 56189
rect 13322 56217 13328 56229
rect 13459 56220 13517 56226
rect 13459 56217 13471 56220
rect 13322 56189 13471 56217
rect 13322 56177 13328 56189
rect 13459 56186 13471 56189
rect 13505 56186 13517 56220
rect 13459 56180 13517 56186
rect 15088 56177 15094 56229
rect 15146 56217 15152 56229
rect 15859 56220 15917 56226
rect 15146 56189 15191 56217
rect 15146 56177 15152 56189
rect 15859 56186 15871 56220
rect 15905 56186 15917 56220
rect 17200 56217 17206 56229
rect 17161 56189 17206 56217
rect 15859 56180 15917 56186
rect 15376 56103 15382 56155
rect 15434 56143 15440 56155
rect 15874 56143 15902 56180
rect 17200 56177 17206 56189
rect 17258 56177 17264 56229
rect 18256 56217 18262 56229
rect 18217 56189 18262 56217
rect 18256 56177 18262 56189
rect 18314 56177 18320 56229
rect 20368 56217 20374 56229
rect 20329 56189 20374 56217
rect 20368 56177 20374 56189
rect 20426 56177 20432 56229
rect 21139 56220 21197 56226
rect 21139 56186 21151 56220
rect 21185 56217 21197 56220
rect 21424 56217 21430 56229
rect 21185 56189 21430 56217
rect 21185 56186 21197 56189
rect 21139 56180 21197 56186
rect 21424 56177 21430 56189
rect 21482 56177 21488 56229
rect 21907 56220 21965 56226
rect 21907 56186 21919 56220
rect 21953 56217 21965 56220
rect 22192 56217 22198 56229
rect 21953 56189 22198 56217
rect 21953 56186 21965 56189
rect 21907 56180 21965 56186
rect 22192 56177 22198 56189
rect 22250 56177 22256 56229
rect 22960 56177 22966 56229
rect 23018 56217 23024 56229
rect 26128 56217 26134 56229
rect 23018 56189 23063 56217
rect 26089 56189 26134 56217
rect 23018 56177 23024 56189
rect 26128 56177 26134 56189
rect 26186 56177 26192 56229
rect 26611 56220 26669 56226
rect 26611 56186 26623 56220
rect 26657 56217 26669 56220
rect 26800 56217 26806 56229
rect 26657 56189 26806 56217
rect 26657 56186 26669 56189
rect 26611 56180 26669 56186
rect 26800 56177 26806 56189
rect 26858 56177 26864 56229
rect 27472 56217 27478 56229
rect 27433 56189 27478 56217
rect 27472 56177 27478 56189
rect 27530 56217 27536 56229
rect 27667 56220 27725 56226
rect 27667 56217 27679 56220
rect 27530 56189 27679 56217
rect 27530 56177 27536 56189
rect 27667 56186 27679 56189
rect 27713 56186 27725 56220
rect 28144 56217 28150 56229
rect 28105 56189 28150 56217
rect 27667 56180 27725 56186
rect 28144 56177 28150 56189
rect 28202 56217 28208 56229
rect 28435 56220 28493 56226
rect 28435 56217 28447 56220
rect 28202 56189 28447 56217
rect 28202 56177 28208 56189
rect 28435 56186 28447 56189
rect 28481 56186 28493 56220
rect 29296 56217 29302 56229
rect 29257 56189 29302 56217
rect 28435 56180 28493 56186
rect 29296 56177 29302 56189
rect 29354 56217 29360 56229
rect 29587 56220 29645 56226
rect 29587 56217 29599 56220
rect 29354 56189 29599 56217
rect 29354 56177 29360 56189
rect 29587 56186 29599 56189
rect 29633 56186 29645 56220
rect 30928 56217 30934 56229
rect 30889 56189 30934 56217
rect 29587 56180 29645 56186
rect 30928 56177 30934 56189
rect 30986 56177 30992 56229
rect 31411 56220 31469 56226
rect 31411 56186 31423 56220
rect 31457 56217 31469 56220
rect 31696 56217 31702 56229
rect 31457 56189 31702 56217
rect 31457 56186 31469 56189
rect 31411 56180 31469 56186
rect 31696 56177 31702 56189
rect 31754 56177 31760 56229
rect 32464 56217 32470 56229
rect 32425 56189 32470 56217
rect 32464 56177 32470 56189
rect 32522 56177 32528 56229
rect 32848 56217 32854 56229
rect 32809 56189 32854 56217
rect 32848 56177 32854 56189
rect 32906 56217 32912 56229
rect 33139 56220 33197 56226
rect 33139 56217 33151 56220
rect 32906 56189 33151 56217
rect 32906 56177 32912 56189
rect 33139 56186 33151 56189
rect 33185 56186 33197 56220
rect 33139 56180 33197 56186
rect 33235 56220 33293 56226
rect 33235 56186 33247 56220
rect 33281 56186 33293 56220
rect 33235 56180 33293 56186
rect 33715 56220 33773 56226
rect 33715 56186 33727 56220
rect 33761 56217 33773 56220
rect 34000 56217 34006 56229
rect 33761 56189 34006 56217
rect 33761 56186 33773 56189
rect 33715 56180 33773 56186
rect 15434 56115 15902 56143
rect 15434 56103 15440 56115
rect 32752 56103 32758 56155
rect 32810 56143 32816 56155
rect 33250 56143 33278 56180
rect 34000 56177 34006 56189
rect 34058 56177 34064 56229
rect 34384 56217 34390 56229
rect 34345 56189 34390 56217
rect 34384 56177 34390 56189
rect 34442 56217 34448 56229
rect 34675 56220 34733 56226
rect 34675 56217 34687 56220
rect 34442 56189 34687 56217
rect 34442 56177 34448 56189
rect 34675 56186 34687 56189
rect 34721 56186 34733 56220
rect 35824 56217 35830 56229
rect 35785 56189 35830 56217
rect 34675 56180 34733 56186
rect 35824 56177 35830 56189
rect 35882 56217 35888 56229
rect 36115 56220 36173 56226
rect 36115 56217 36127 56220
rect 35882 56189 36127 56217
rect 35882 56177 35888 56189
rect 36115 56186 36127 56189
rect 36161 56186 36173 56220
rect 36115 56180 36173 56186
rect 36211 56220 36269 56226
rect 36211 56186 36223 56220
rect 36257 56186 36269 56220
rect 36211 56180 36269 56186
rect 36691 56220 36749 56226
rect 36691 56186 36703 56220
rect 36737 56217 36749 56220
rect 36784 56217 36790 56229
rect 36737 56189 36790 56217
rect 36737 56186 36749 56189
rect 36691 56180 36749 56186
rect 32810 56115 33278 56143
rect 32810 56103 32816 56115
rect 35440 56103 35446 56155
rect 35498 56143 35504 56155
rect 36226 56143 36254 56180
rect 36784 56177 36790 56189
rect 36842 56217 36848 56229
rect 36883 56220 36941 56226
rect 36883 56217 36895 56220
rect 36842 56189 36895 56217
rect 36842 56177 36848 56189
rect 36883 56186 36895 56189
rect 36929 56186 36941 56220
rect 36883 56180 36941 56186
rect 37459 56220 37517 56226
rect 37459 56186 37471 56220
rect 37505 56217 37517 56220
rect 37744 56217 37750 56229
rect 37505 56189 37750 56217
rect 37505 56186 37517 56189
rect 37459 56180 37517 56186
rect 37744 56177 37750 56189
rect 37802 56177 37808 56229
rect 38515 56220 38573 56226
rect 38515 56186 38527 56220
rect 38561 56217 38573 56220
rect 38704 56217 38710 56229
rect 38561 56189 38710 56217
rect 38561 56186 38573 56189
rect 38515 56180 38573 56186
rect 38704 56177 38710 56189
rect 38762 56177 38768 56229
rect 39856 56217 39862 56229
rect 39817 56189 39862 56217
rect 39856 56177 39862 56189
rect 39914 56217 39920 56229
rect 40243 56220 40301 56226
rect 40243 56217 40255 56220
rect 39914 56189 40255 56217
rect 39914 56177 39920 56189
rect 40243 56186 40255 56189
rect 40289 56186 40301 56220
rect 40243 56180 40301 56186
rect 41968 56177 41974 56229
rect 42026 56217 42032 56229
rect 42451 56220 42509 56226
rect 42026 56189 42071 56217
rect 42026 56177 42032 56189
rect 42451 56186 42463 56220
rect 42497 56217 42509 56220
rect 42640 56217 42646 56229
rect 42497 56189 42646 56217
rect 42497 56186 42509 56189
rect 42451 56180 42509 56186
rect 42640 56177 42646 56189
rect 42698 56177 42704 56229
rect 43219 56220 43277 56226
rect 43219 56186 43231 56220
rect 43265 56217 43277 56220
rect 43411 56220 43469 56226
rect 43411 56217 43423 56220
rect 43265 56189 43423 56217
rect 43265 56186 43277 56189
rect 43219 56180 43277 56186
rect 43411 56186 43423 56189
rect 43457 56217 43469 56220
rect 43600 56217 43606 56229
rect 43457 56189 43606 56217
rect 43457 56186 43469 56189
rect 43411 56180 43469 56186
rect 43600 56177 43606 56189
rect 43658 56177 43664 56229
rect 43987 56220 44045 56226
rect 43987 56186 43999 56220
rect 44033 56217 44045 56220
rect 44176 56217 44182 56229
rect 44033 56189 44182 56217
rect 44033 56186 44045 56189
rect 43987 56180 44045 56186
rect 44176 56177 44182 56189
rect 44234 56177 44240 56229
rect 44851 56220 44909 56226
rect 44851 56186 44863 56220
rect 44897 56217 44909 56220
rect 45040 56217 45046 56229
rect 44897 56189 45046 56217
rect 44897 56186 44909 56189
rect 44851 56180 44909 56186
rect 45040 56177 45046 56189
rect 45098 56177 45104 56229
rect 46768 56217 46774 56229
rect 46729 56189 46774 56217
rect 46768 56177 46774 56189
rect 46826 56177 46832 56229
rect 48208 56217 48214 56229
rect 48169 56189 48214 56217
rect 48208 56177 48214 56189
rect 48266 56177 48272 56229
rect 48691 56220 48749 56226
rect 48691 56186 48703 56220
rect 48737 56217 48749 56220
rect 48784 56217 48790 56229
rect 48737 56189 48790 56217
rect 48737 56186 48749 56189
rect 48691 56180 48749 56186
rect 48784 56177 48790 56189
rect 48842 56217 48848 56229
rect 48883 56220 48941 56226
rect 48883 56217 48895 56220
rect 48842 56189 48895 56217
rect 48842 56177 48848 56189
rect 48883 56186 48895 56189
rect 48929 56186 48941 56220
rect 48883 56180 48941 56186
rect 48979 56220 49037 56226
rect 48979 56186 48991 56220
rect 49025 56186 49037 56220
rect 48979 56180 49037 56186
rect 49843 56220 49901 56226
rect 49843 56186 49855 56220
rect 49889 56186 49901 56220
rect 49843 56180 49901 56186
rect 35498 56115 36254 56143
rect 35498 56103 35504 56115
rect 37072 56103 37078 56155
rect 37130 56143 37136 56155
rect 40816 56143 40822 56155
rect 37130 56115 40822 56143
rect 37130 56103 37136 56115
rect 40816 56103 40822 56115
rect 40874 56103 40880 56155
rect 48592 56103 48598 56155
rect 48650 56143 48656 56155
rect 48994 56143 49022 56180
rect 48650 56115 49022 56143
rect 48650 56103 48656 56115
rect 38800 56029 38806 56081
rect 38858 56069 38864 56081
rect 49858 56069 49886 56180
rect 49936 56177 49942 56229
rect 49994 56217 50000 56229
rect 50611 56220 50669 56226
rect 50611 56217 50623 56220
rect 49994 56189 50623 56217
rect 49994 56177 50000 56189
rect 50611 56186 50623 56189
rect 50657 56186 50669 56220
rect 51664 56217 51670 56229
rect 51625 56189 51670 56217
rect 50611 56180 50669 56186
rect 51664 56177 51670 56189
rect 51722 56217 51728 56229
rect 51955 56220 52013 56226
rect 51955 56217 51967 56220
rect 51722 56189 51967 56217
rect 51722 56177 51728 56189
rect 51955 56186 51967 56189
rect 52001 56186 52013 56220
rect 51955 56180 52013 56186
rect 52051 56220 52109 56226
rect 52051 56186 52063 56220
rect 52097 56186 52109 56220
rect 52051 56180 52109 56186
rect 53491 56220 53549 56226
rect 53491 56186 53503 56220
rect 53537 56217 53549 56220
rect 53680 56217 53686 56229
rect 53537 56189 53686 56217
rect 53537 56186 53549 56189
rect 53491 56180 53549 56186
rect 51184 56103 51190 56155
rect 51242 56143 51248 56155
rect 52066 56143 52094 56180
rect 53680 56177 53686 56189
rect 53738 56177 53744 56229
rect 54544 56217 54550 56229
rect 54505 56189 54550 56217
rect 54544 56177 54550 56189
rect 54602 56177 54608 56229
rect 55027 56220 55085 56226
rect 55027 56186 55039 56220
rect 55073 56217 55085 56220
rect 55219 56220 55277 56226
rect 55219 56217 55231 56220
rect 55073 56189 55231 56217
rect 55073 56186 55085 56189
rect 55027 56180 55085 56186
rect 55219 56186 55231 56189
rect 55265 56217 55277 56220
rect 55504 56217 55510 56229
rect 55265 56189 55510 56217
rect 55265 56186 55277 56189
rect 55219 56180 55277 56186
rect 55504 56177 55510 56189
rect 55562 56177 55568 56229
rect 51242 56115 52094 56143
rect 51242 56103 51248 56115
rect 38858 56041 49886 56069
rect 38858 56029 38864 56041
rect 1152 55970 58848 55992
rect 1152 55918 4294 55970
rect 4346 55918 4358 55970
rect 4410 55918 4422 55970
rect 4474 55918 4486 55970
rect 4538 55918 35014 55970
rect 35066 55918 35078 55970
rect 35130 55918 35142 55970
rect 35194 55918 35206 55970
rect 35258 55918 58848 55970
rect 1152 55896 58848 55918
rect 3760 55733 3766 55785
rect 3818 55773 3824 55785
rect 9715 55776 9773 55782
rect 9715 55773 9727 55776
rect 3818 55745 9727 55773
rect 3818 55733 3824 55745
rect 9715 55742 9727 55745
rect 9761 55773 9773 55776
rect 9907 55776 9965 55782
rect 9907 55773 9919 55776
rect 9761 55745 9919 55773
rect 9761 55742 9773 55745
rect 9715 55736 9773 55742
rect 9907 55742 9919 55745
rect 9953 55742 9965 55776
rect 9907 55736 9965 55742
rect 11920 55733 11926 55785
rect 11978 55773 11984 55785
rect 11978 55745 17294 55773
rect 11978 55733 11984 55745
rect 1168 55659 1174 55711
rect 1226 55699 1232 55711
rect 1651 55702 1709 55708
rect 1651 55699 1663 55702
rect 1226 55671 1663 55699
rect 1226 55659 1232 55671
rect 1651 55668 1663 55671
rect 1697 55668 1709 55702
rect 1651 55662 1709 55668
rect 4435 55702 4493 55708
rect 4435 55668 4447 55702
rect 4481 55699 4493 55702
rect 4624 55699 4630 55711
rect 4481 55671 4630 55699
rect 4481 55668 4493 55671
rect 4435 55662 4493 55668
rect 4624 55659 4630 55671
rect 4682 55659 4688 55711
rect 7504 55659 7510 55711
rect 7562 55699 7568 55711
rect 7603 55702 7661 55708
rect 7603 55699 7615 55702
rect 7562 55671 7615 55699
rect 7562 55659 7568 55671
rect 7603 55668 7615 55671
rect 7649 55668 7661 55702
rect 7603 55662 7661 55668
rect 9136 55659 9142 55711
rect 9194 55699 9200 55711
rect 9331 55702 9389 55708
rect 9331 55699 9343 55702
rect 9194 55671 9343 55699
rect 9194 55659 9200 55671
rect 9331 55668 9343 55671
rect 9377 55668 9389 55702
rect 9331 55662 9389 55668
rect 13840 55659 13846 55711
rect 13898 55699 13904 55711
rect 13939 55702 13997 55708
rect 13939 55699 13951 55702
rect 13898 55671 13951 55699
rect 13898 55659 13904 55671
rect 13939 55668 13951 55671
rect 13985 55668 13997 55702
rect 13939 55662 13997 55668
rect 5008 55585 5014 55637
rect 5066 55625 5072 55637
rect 14035 55628 14093 55634
rect 14035 55625 14047 55628
rect 5066 55597 14047 55625
rect 5066 55585 5072 55597
rect 14035 55594 14047 55597
rect 14081 55594 14093 55628
rect 17266 55625 17294 55745
rect 27346 55745 48062 55773
rect 20176 55659 20182 55711
rect 20234 55699 20240 55711
rect 20275 55702 20333 55708
rect 20275 55699 20287 55702
rect 20234 55671 20287 55699
rect 20234 55659 20240 55671
rect 20275 55668 20287 55671
rect 20321 55668 20333 55702
rect 20275 55662 20333 55668
rect 23344 55659 23350 55711
rect 23402 55699 23408 55711
rect 23539 55702 23597 55708
rect 23539 55699 23551 55702
rect 23402 55671 23551 55699
rect 23402 55659 23408 55671
rect 23539 55668 23551 55671
rect 23585 55668 23597 55702
rect 23539 55662 23597 55668
rect 24880 55659 24886 55711
rect 24938 55699 24944 55711
rect 25075 55702 25133 55708
rect 25075 55699 25087 55702
rect 24938 55671 25087 55699
rect 24938 55659 24944 55671
rect 25075 55668 25087 55671
rect 25121 55668 25133 55702
rect 25075 55662 25133 55668
rect 27346 55625 27374 55745
rect 39088 55659 39094 55711
rect 39146 55699 39152 55711
rect 39283 55702 39341 55708
rect 39283 55699 39295 55702
rect 39146 55671 39295 55699
rect 39146 55659 39152 55671
rect 39283 55668 39295 55671
rect 39329 55668 39341 55702
rect 39283 55662 39341 55668
rect 40720 55659 40726 55711
rect 40778 55699 40784 55711
rect 40915 55702 40973 55708
rect 40915 55699 40927 55702
rect 40778 55671 40927 55699
rect 40778 55659 40784 55671
rect 40915 55668 40927 55671
rect 40961 55668 40973 55702
rect 40915 55662 40973 55668
rect 45424 55659 45430 55711
rect 45482 55699 45488 55711
rect 45619 55702 45677 55708
rect 45619 55699 45631 55702
rect 45482 55671 45631 55699
rect 45482 55659 45488 55671
rect 45619 55668 45631 55671
rect 45665 55668 45677 55702
rect 45619 55662 45677 55668
rect 46960 55659 46966 55711
rect 47018 55699 47024 55711
rect 48034 55708 48062 55745
rect 47155 55702 47213 55708
rect 47155 55699 47167 55702
rect 47018 55671 47167 55699
rect 47018 55659 47024 55671
rect 47155 55668 47167 55671
rect 47201 55668 47213 55702
rect 47155 55662 47213 55668
rect 48019 55702 48077 55708
rect 48019 55668 48031 55702
rect 48065 55668 48077 55702
rect 48019 55662 48077 55668
rect 51760 55659 51766 55711
rect 51818 55699 51824 55711
rect 51955 55702 52013 55708
rect 51955 55699 51967 55702
rect 51818 55671 51967 55699
rect 51818 55659 51824 55671
rect 51955 55668 51967 55671
rect 52001 55668 52013 55702
rect 51955 55662 52013 55668
rect 56464 55659 56470 55711
rect 56522 55699 56528 55711
rect 56659 55702 56717 55708
rect 56659 55699 56671 55702
rect 56522 55671 56671 55699
rect 56522 55659 56528 55671
rect 56659 55668 56671 55671
rect 56705 55668 56717 55702
rect 56659 55662 56717 55668
rect 57520 55659 57526 55711
rect 57578 55699 57584 55711
rect 57715 55702 57773 55708
rect 57715 55699 57727 55702
rect 57578 55671 57727 55699
rect 57578 55659 57584 55671
rect 57715 55668 57727 55671
rect 57761 55668 57773 55702
rect 57715 55662 57773 55668
rect 52624 55625 52630 55637
rect 17266 55597 27374 55625
rect 38818 55597 52630 55625
rect 14035 55588 14093 55594
rect 1744 55551 1750 55563
rect 1705 55523 1750 55551
rect 1744 55511 1750 55523
rect 1802 55551 1808 55563
rect 1939 55554 1997 55560
rect 1939 55551 1951 55554
rect 1802 55523 1951 55551
rect 1802 55511 1808 55523
rect 1939 55520 1951 55523
rect 1985 55520 1997 55554
rect 1939 55514 1997 55520
rect 4243 55554 4301 55560
rect 4243 55520 4255 55554
rect 4289 55551 4301 55554
rect 4531 55554 4589 55560
rect 4531 55551 4543 55554
rect 4289 55523 4543 55551
rect 4289 55520 4301 55523
rect 4243 55514 4301 55520
rect 4531 55520 4543 55523
rect 4577 55551 4589 55554
rect 4624 55551 4630 55563
rect 4577 55523 4630 55551
rect 4577 55520 4589 55523
rect 4531 55514 4589 55520
rect 4624 55511 4630 55523
rect 4682 55511 4688 55563
rect 7411 55554 7469 55560
rect 7411 55520 7423 55554
rect 7457 55551 7469 55554
rect 7696 55551 7702 55563
rect 7457 55523 7702 55551
rect 7457 55520 7469 55523
rect 7411 55514 7469 55520
rect 7696 55511 7702 55523
rect 7754 55511 7760 55563
rect 9235 55554 9293 55560
rect 9235 55551 9247 55554
rect 8962 55523 9247 55551
rect 8962 55415 8990 55523
rect 9235 55520 9247 55523
rect 9281 55520 9293 55554
rect 9235 55514 9293 55520
rect 12499 55554 12557 55560
rect 12499 55520 12511 55554
rect 12545 55551 12557 55554
rect 12784 55551 12790 55563
rect 12545 55523 12790 55551
rect 12545 55520 12557 55523
rect 12499 55514 12557 55520
rect 12784 55511 12790 55523
rect 12842 55511 12848 55563
rect 15283 55554 15341 55560
rect 15283 55520 15295 55554
rect 15329 55551 15341 55554
rect 15571 55554 15629 55560
rect 15571 55551 15583 55554
rect 15329 55523 15583 55551
rect 15329 55520 15341 55523
rect 15283 55514 15341 55520
rect 15571 55520 15583 55523
rect 15617 55551 15629 55554
rect 16528 55551 16534 55563
rect 15617 55523 16534 55551
rect 15617 55520 15629 55523
rect 15571 55514 15629 55520
rect 16528 55511 16534 55523
rect 16586 55511 16592 55563
rect 20272 55511 20278 55563
rect 20330 55551 20336 55563
rect 20371 55554 20429 55560
rect 20371 55551 20383 55554
rect 20330 55523 20383 55551
rect 20330 55511 20336 55523
rect 20371 55520 20383 55523
rect 20417 55520 20429 55554
rect 20371 55514 20429 55520
rect 23152 55511 23158 55563
rect 23210 55551 23216 55563
rect 23443 55554 23501 55560
rect 23443 55551 23455 55554
rect 23210 55523 23455 55551
rect 23210 55511 23216 55523
rect 23443 55520 23455 55523
rect 23489 55520 23501 55554
rect 23443 55514 23501 55520
rect 24880 55511 24886 55563
rect 24938 55551 24944 55563
rect 24979 55554 25037 55560
rect 24979 55551 24991 55554
rect 24938 55523 24991 55551
rect 24938 55511 24944 55523
rect 24979 55520 24991 55523
rect 25025 55520 25037 55554
rect 25648 55551 25654 55563
rect 25609 55523 25654 55551
rect 24979 55514 25037 55520
rect 25648 55511 25654 55523
rect 25706 55511 25712 55563
rect 29107 55554 29165 55560
rect 29107 55520 29119 55554
rect 29153 55551 29165 55554
rect 38818 55551 38846 55597
rect 52624 55585 52630 55597
rect 52682 55585 52688 55637
rect 39187 55554 39245 55560
rect 39187 55551 39199 55554
rect 29153 55523 38846 55551
rect 38914 55523 39199 55551
rect 29153 55520 29165 55523
rect 29107 55514 29165 55520
rect 14707 55480 14765 55486
rect 14707 55446 14719 55480
rect 14753 55477 14765 55480
rect 38800 55477 38806 55489
rect 14753 55449 38806 55477
rect 14753 55446 14765 55449
rect 14707 55440 14765 55446
rect 38800 55437 38806 55449
rect 38858 55437 38864 55489
rect 38914 55415 38942 55523
rect 39187 55520 39199 55523
rect 39233 55520 39245 55554
rect 40819 55554 40877 55560
rect 40819 55551 40831 55554
rect 39187 55514 39245 55520
rect 40546 55523 40831 55551
rect 8944 55403 8950 55415
rect 8905 55375 8950 55403
rect 8944 55363 8950 55375
rect 9002 55363 9008 55415
rect 23152 55403 23158 55415
rect 23113 55375 23158 55403
rect 23152 55363 23158 55375
rect 23210 55363 23216 55415
rect 24787 55406 24845 55412
rect 24787 55372 24799 55406
rect 24833 55403 24845 55406
rect 24880 55403 24886 55415
rect 24833 55375 24886 55403
rect 24833 55372 24845 55375
rect 24787 55366 24845 55372
rect 24880 55363 24886 55375
rect 24938 55363 24944 55415
rect 25555 55406 25613 55412
rect 25555 55372 25567 55406
rect 25601 55403 25613 55406
rect 25648 55403 25654 55415
rect 25601 55375 25654 55403
rect 25601 55372 25613 55375
rect 25555 55366 25613 55372
rect 25648 55363 25654 55375
rect 25706 55363 25712 55415
rect 38896 55403 38902 55415
rect 38857 55375 38902 55403
rect 38896 55363 38902 55375
rect 38954 55363 38960 55415
rect 40432 55363 40438 55415
rect 40490 55403 40496 55415
rect 40546 55412 40574 55523
rect 40819 55520 40831 55523
rect 40865 55551 40877 55554
rect 41107 55554 41165 55560
rect 41107 55551 41119 55554
rect 40865 55523 41119 55551
rect 40865 55520 40877 55523
rect 40819 55514 40877 55520
rect 41107 55520 41119 55523
rect 41153 55520 41165 55554
rect 41107 55514 41165 55520
rect 42547 55554 42605 55560
rect 42547 55520 42559 55554
rect 42593 55520 42605 55554
rect 45523 55554 45581 55560
rect 45523 55551 45535 55554
rect 42547 55514 42605 55520
rect 45250 55523 45535 55551
rect 40531 55406 40589 55412
rect 40531 55403 40543 55406
rect 40490 55375 40543 55403
rect 40490 55363 40496 55375
rect 40531 55372 40543 55375
rect 40577 55372 40589 55406
rect 42160 55403 42166 55415
rect 42121 55375 42166 55403
rect 40531 55366 40589 55372
rect 42160 55363 42166 55375
rect 42218 55403 42224 55415
rect 42562 55403 42590 55514
rect 45250 55415 45278 55523
rect 45523 55520 45535 55523
rect 45569 55520 45581 55554
rect 47059 55554 47117 55560
rect 47059 55551 47071 55554
rect 45523 55514 45581 55520
rect 46786 55523 47071 55551
rect 45232 55403 45238 55415
rect 42218 55375 42590 55403
rect 45193 55375 45238 55403
rect 42218 55363 42224 55375
rect 45232 55363 45238 55375
rect 45290 55363 45296 55415
rect 46576 55363 46582 55415
rect 46634 55403 46640 55415
rect 46786 55412 46814 55523
rect 47059 55520 47071 55523
rect 47105 55551 47117 55554
rect 47347 55554 47405 55560
rect 47347 55551 47359 55554
rect 47105 55523 47359 55551
rect 47105 55520 47117 55523
rect 47059 55514 47117 55520
rect 47347 55520 47359 55523
rect 47393 55520 47405 55554
rect 51859 55554 51917 55560
rect 51859 55551 51871 55554
rect 47347 55514 47405 55520
rect 51586 55523 51871 55551
rect 51586 55415 51614 55523
rect 51859 55520 51871 55523
rect 51905 55520 51917 55554
rect 55795 55554 55853 55560
rect 55795 55551 55807 55554
rect 51859 55514 51917 55520
rect 55618 55523 55807 55551
rect 55618 55415 55646 55523
rect 55795 55520 55807 55523
rect 55841 55520 55853 55554
rect 55795 55514 55853 55520
rect 56563 55554 56621 55560
rect 56563 55520 56575 55554
rect 56609 55520 56621 55554
rect 57619 55554 57677 55560
rect 57619 55551 57631 55554
rect 56563 55514 56621 55520
rect 57346 55523 57631 55551
rect 46771 55406 46829 55412
rect 46771 55403 46783 55406
rect 46634 55375 46783 55403
rect 46634 55363 46640 55375
rect 46771 55372 46783 55375
rect 46817 55372 46829 55406
rect 51568 55403 51574 55415
rect 51529 55375 51574 55403
rect 46771 55366 46829 55372
rect 51568 55363 51574 55375
rect 51626 55363 51632 55415
rect 55600 55403 55606 55415
rect 55561 55375 55606 55403
rect 55600 55363 55606 55375
rect 55658 55363 55664 55415
rect 56272 55403 56278 55415
rect 56233 55375 56278 55403
rect 56272 55363 56278 55375
rect 56330 55403 56336 55415
rect 56578 55403 56606 55514
rect 57346 55415 57374 55523
rect 57619 55520 57631 55523
rect 57665 55520 57677 55554
rect 57619 55514 57677 55520
rect 57328 55403 57334 55415
rect 56330 55375 56606 55403
rect 57289 55375 57334 55403
rect 56330 55363 56336 55375
rect 57328 55363 57334 55375
rect 57386 55363 57392 55415
rect 1152 55304 58848 55326
rect 1152 55252 19654 55304
rect 19706 55252 19718 55304
rect 19770 55252 19782 55304
rect 19834 55252 19846 55304
rect 19898 55252 50374 55304
rect 50426 55252 50438 55304
rect 50490 55252 50502 55304
rect 50554 55252 50566 55304
rect 50618 55252 58848 55304
rect 1152 55230 58848 55252
rect 19984 55141 19990 55193
rect 20042 55181 20048 55193
rect 55600 55181 55606 55193
rect 20042 55153 55606 55181
rect 20042 55141 20048 55153
rect 55600 55141 55606 55153
rect 55658 55141 55664 55193
rect 57811 55184 57869 55190
rect 57811 55150 57823 55184
rect 57857 55181 57869 55184
rect 59152 55181 59158 55193
rect 57857 55153 59158 55181
rect 57857 55150 57869 55153
rect 57811 55144 57869 55150
rect 59152 55141 59158 55153
rect 59210 55141 59216 55193
rect 11440 54993 11446 55045
rect 11498 55033 11504 55045
rect 12019 55036 12077 55042
rect 12019 55033 12031 55036
rect 11498 55005 12031 55033
rect 11498 54993 11504 55005
rect 12019 55002 12031 55005
rect 12065 55002 12077 55036
rect 12019 54996 12077 55002
rect 57619 54888 57677 54894
rect 57619 54854 57631 54888
rect 57665 54885 57677 54888
rect 57907 54888 57965 54894
rect 57907 54885 57919 54888
rect 57665 54857 57919 54885
rect 57665 54854 57677 54857
rect 57619 54848 57677 54854
rect 57907 54854 57919 54857
rect 57953 54885 57965 54888
rect 58000 54885 58006 54897
rect 57953 54857 58006 54885
rect 57953 54854 57965 54857
rect 57907 54848 57965 54854
rect 58000 54845 58006 54857
rect 58058 54845 58064 54897
rect 25843 54740 25901 54746
rect 25843 54706 25855 54740
rect 25889 54737 25901 54740
rect 26131 54740 26189 54746
rect 26131 54737 26143 54740
rect 25889 54709 26143 54737
rect 25889 54706 25901 54709
rect 25843 54700 25901 54706
rect 26131 54706 26143 54709
rect 26177 54737 26189 54740
rect 30064 54737 30070 54749
rect 26177 54709 30070 54737
rect 26177 54706 26189 54709
rect 26131 54700 26189 54706
rect 30064 54697 30070 54709
rect 30122 54697 30128 54749
rect 44656 54737 44662 54749
rect 44617 54709 44662 54737
rect 44656 54697 44662 54709
rect 44714 54737 44720 54749
rect 44851 54740 44909 54746
rect 44851 54737 44863 54740
rect 44714 54709 44863 54737
rect 44714 54697 44720 54709
rect 44851 54706 44863 54709
rect 44897 54706 44909 54740
rect 55792 54737 55798 54749
rect 55753 54709 55798 54737
rect 44851 54700 44909 54706
rect 55792 54697 55798 54709
rect 55850 54737 55856 54749
rect 55987 54740 56045 54746
rect 55987 54737 55999 54740
rect 55850 54709 55999 54737
rect 55850 54697 55856 54709
rect 55987 54706 55999 54709
rect 56033 54706 56045 54740
rect 55987 54700 56045 54706
rect 1152 54638 58848 54660
rect 1152 54586 4294 54638
rect 4346 54586 4358 54638
rect 4410 54586 4422 54638
rect 4474 54586 4486 54638
rect 4538 54586 35014 54638
rect 35066 54586 35078 54638
rect 35130 54586 35142 54638
rect 35194 54586 35206 54638
rect 35258 54586 58848 54638
rect 1152 54564 58848 54586
rect 57907 54370 57965 54376
rect 57907 54336 57919 54370
rect 57953 54367 57965 54370
rect 58096 54367 58102 54379
rect 57953 54339 58102 54367
rect 57953 54336 57965 54339
rect 57907 54330 57965 54336
rect 58096 54327 58102 54339
rect 58154 54327 58160 54379
rect 14131 54222 14189 54228
rect 14131 54188 14143 54222
rect 14177 54188 14189 54222
rect 14131 54182 14189 54188
rect 49075 54222 49133 54228
rect 49075 54188 49087 54222
rect 49121 54219 49133 54222
rect 49363 54222 49421 54228
rect 49363 54219 49375 54222
rect 49121 54191 49375 54219
rect 49121 54188 49133 54191
rect 49075 54182 49133 54188
rect 49363 54188 49375 54191
rect 49409 54219 49421 54222
rect 53008 54219 53014 54231
rect 49409 54191 53014 54219
rect 49409 54188 49421 54191
rect 49363 54182 49421 54188
rect 13843 54148 13901 54154
rect 13843 54114 13855 54148
rect 13889 54145 13901 54148
rect 14146 54145 14174 54182
rect 53008 54179 53014 54191
rect 53066 54179 53072 54231
rect 57616 54179 57622 54231
rect 57674 54219 57680 54231
rect 57811 54222 57869 54228
rect 57811 54219 57823 54222
rect 57674 54191 57823 54219
rect 57674 54179 57680 54191
rect 57811 54188 57823 54191
rect 57857 54188 57869 54222
rect 57811 54182 57869 54188
rect 36496 54145 36502 54157
rect 13889 54117 36502 54145
rect 13889 54114 13901 54117
rect 13843 54108 13901 54114
rect 36496 54105 36502 54117
rect 36554 54105 36560 54157
rect 36880 54105 36886 54157
rect 36938 54145 36944 54157
rect 55792 54145 55798 54157
rect 36938 54117 55798 54145
rect 36938 54105 36944 54117
rect 55792 54105 55798 54117
rect 55850 54105 55856 54157
rect 1152 53972 58848 53994
rect 1152 53920 19654 53972
rect 19706 53920 19718 53972
rect 19770 53920 19782 53972
rect 19834 53920 19846 53972
rect 19898 53920 50374 53972
rect 50426 53920 50438 53972
rect 50490 53920 50502 53972
rect 50554 53920 50566 53972
rect 50618 53920 58848 53972
rect 1152 53898 58848 53920
rect 10864 53809 10870 53861
rect 10922 53849 10928 53861
rect 57616 53849 57622 53861
rect 10922 53821 57622 53849
rect 10922 53809 10928 53821
rect 57616 53809 57622 53821
rect 57674 53809 57680 53861
rect 57907 53852 57965 53858
rect 57907 53818 57919 53852
rect 57953 53849 57965 53852
rect 59632 53849 59638 53861
rect 57953 53821 59638 53849
rect 57953 53818 57965 53821
rect 57907 53812 57965 53818
rect 59632 53809 59638 53821
rect 59690 53809 59696 53861
rect 57811 53556 57869 53562
rect 57811 53553 57823 53556
rect 57634 53525 57823 53553
rect 57634 53417 57662 53525
rect 57811 53522 57823 53525
rect 57857 53522 57869 53556
rect 57811 53516 57869 53522
rect 6448 53365 6454 53417
rect 6506 53405 6512 53417
rect 26803 53408 26861 53414
rect 26803 53405 26815 53408
rect 6506 53377 26815 53405
rect 6506 53365 6512 53377
rect 26803 53374 26815 53377
rect 26849 53405 26861 53408
rect 26995 53408 27053 53414
rect 26995 53405 27007 53408
rect 26849 53377 27007 53405
rect 26849 53374 26861 53377
rect 26803 53368 26861 53374
rect 26995 53374 27007 53377
rect 27041 53374 27053 53408
rect 26995 53368 27053 53374
rect 57616 53365 57622 53417
rect 57674 53405 57680 53417
rect 57674 53377 57719 53405
rect 57674 53365 57680 53377
rect 1152 53306 58848 53328
rect 1152 53254 4294 53306
rect 4346 53254 4358 53306
rect 4410 53254 4422 53306
rect 4474 53254 4486 53306
rect 4538 53254 35014 53306
rect 35066 53254 35078 53306
rect 35130 53254 35142 53306
rect 35194 53254 35206 53306
rect 35258 53254 58848 53306
rect 1152 53232 58848 53254
rect 23923 52890 23981 52896
rect 23923 52856 23935 52890
rect 23969 52887 23981 52890
rect 24211 52890 24269 52896
rect 24211 52887 24223 52890
rect 23969 52859 24223 52887
rect 23969 52856 23981 52859
rect 23923 52850 23981 52856
rect 24211 52856 24223 52859
rect 24257 52856 24269 52890
rect 24211 52850 24269 52856
rect 40819 52890 40877 52896
rect 40819 52856 40831 52890
rect 40865 52887 40877 52890
rect 41107 52890 41165 52896
rect 41107 52887 41119 52890
rect 40865 52859 41119 52887
rect 40865 52856 40877 52859
rect 40819 52850 40877 52856
rect 41107 52856 41119 52859
rect 41153 52887 41165 52890
rect 48880 52887 48886 52899
rect 41153 52859 48886 52887
rect 41153 52856 41165 52859
rect 41107 52850 41165 52856
rect 48880 52847 48886 52859
rect 48938 52847 48944 52899
rect 21331 52816 21389 52822
rect 21331 52782 21343 52816
rect 21377 52813 21389 52816
rect 30928 52813 30934 52825
rect 21377 52785 30934 52813
rect 21377 52782 21389 52785
rect 21331 52776 21389 52782
rect 30928 52773 30934 52785
rect 30986 52773 30992 52825
rect 22672 52699 22678 52751
rect 22730 52739 22736 52751
rect 23923 52742 23981 52748
rect 23923 52739 23935 52742
rect 22730 52711 23935 52739
rect 22730 52699 22736 52711
rect 23923 52708 23935 52711
rect 23969 52739 23981 52742
rect 24019 52742 24077 52748
rect 24019 52739 24031 52742
rect 23969 52711 24031 52739
rect 23969 52708 23981 52711
rect 23923 52702 23981 52708
rect 24019 52708 24031 52711
rect 24065 52708 24077 52742
rect 24019 52702 24077 52708
rect 1152 52640 58848 52662
rect 1152 52588 19654 52640
rect 19706 52588 19718 52640
rect 19770 52588 19782 52640
rect 19834 52588 19846 52640
rect 19898 52588 50374 52640
rect 50426 52588 50438 52640
rect 50490 52588 50502 52640
rect 50554 52588 50566 52640
rect 50618 52588 58848 52640
rect 1152 52566 58848 52588
rect 37075 52224 37133 52230
rect 37075 52190 37087 52224
rect 37121 52221 37133 52224
rect 46768 52221 46774 52233
rect 37121 52193 46774 52221
rect 37121 52190 37133 52193
rect 37075 52184 37133 52190
rect 46768 52181 46774 52193
rect 46826 52181 46832 52233
rect 42832 52073 42838 52085
rect 42793 52045 42838 52073
rect 42832 52033 42838 52045
rect 42890 52073 42896 52085
rect 43027 52076 43085 52082
rect 43027 52073 43039 52076
rect 42890 52045 43039 52073
rect 42890 52033 42896 52045
rect 43027 52042 43039 52045
rect 43073 52042 43085 52076
rect 43027 52036 43085 52042
rect 1152 51974 58848 51996
rect 1152 51922 4294 51974
rect 4346 51922 4358 51974
rect 4410 51922 4422 51974
rect 4474 51922 4486 51974
rect 4538 51922 35014 51974
rect 35066 51922 35078 51974
rect 35130 51922 35142 51974
rect 35194 51922 35206 51974
rect 35258 51922 58848 51974
rect 1152 51900 58848 51922
rect 7186 51601 27374 51629
rect 1651 51558 1709 51564
rect 1651 51524 1663 51558
rect 1697 51555 1709 51558
rect 1936 51555 1942 51567
rect 1697 51527 1942 51555
rect 1697 51524 1709 51527
rect 1651 51518 1709 51524
rect 1936 51515 1942 51527
rect 1994 51515 2000 51567
rect 5683 51558 5741 51564
rect 5683 51524 5695 51558
rect 5729 51555 5741 51558
rect 5971 51558 6029 51564
rect 5971 51555 5983 51558
rect 5729 51527 5983 51555
rect 5729 51524 5741 51527
rect 5683 51518 5741 51524
rect 5971 51524 5983 51527
rect 6017 51555 6029 51558
rect 7186 51555 7214 51601
rect 6017 51527 7214 51555
rect 20083 51558 20141 51564
rect 6017 51524 6029 51527
rect 5971 51518 6029 51524
rect 20083 51524 20095 51558
rect 20129 51524 20141 51558
rect 27346 51555 27374 51601
rect 52912 51555 52918 51567
rect 27346 51527 52918 51555
rect 20083 51518 20141 51524
rect 19795 51484 19853 51490
rect 19795 51450 19807 51484
rect 19841 51481 19853 51484
rect 20098 51481 20126 51518
rect 52912 51515 52918 51527
rect 52970 51515 52976 51567
rect 48592 51481 48598 51493
rect 19841 51453 48598 51481
rect 19841 51450 19853 51453
rect 19795 51444 19853 51450
rect 48592 51441 48598 51453
rect 48650 51441 48656 51493
rect 1152 51308 58848 51330
rect 1152 51256 19654 51308
rect 19706 51256 19718 51308
rect 19770 51256 19782 51308
rect 19834 51256 19846 51308
rect 19898 51256 50374 51308
rect 50426 51256 50438 51308
rect 50490 51256 50502 51308
rect 50554 51256 50566 51308
rect 50618 51256 58848 51308
rect 1152 51234 58848 51256
rect 1936 51145 1942 51197
rect 1994 51185 2000 51197
rect 32368 51185 32374 51197
rect 1994 51157 32374 51185
rect 1994 51145 2000 51157
rect 32368 51145 32374 51157
rect 32426 51145 32432 51197
rect 25363 50744 25421 50750
rect 25363 50710 25375 50744
rect 25409 50741 25421 50744
rect 25651 50744 25709 50750
rect 25651 50741 25663 50744
rect 25409 50713 25663 50741
rect 25409 50710 25421 50713
rect 25363 50704 25421 50710
rect 25651 50710 25663 50713
rect 25697 50741 25709 50744
rect 31312 50741 31318 50753
rect 25697 50713 31318 50741
rect 25697 50710 25709 50713
rect 25651 50704 25709 50710
rect 31312 50701 31318 50713
rect 31370 50701 31376 50753
rect 31504 50741 31510 50753
rect 31465 50713 31510 50741
rect 31504 50701 31510 50713
rect 31562 50741 31568 50753
rect 31699 50744 31757 50750
rect 31699 50741 31711 50744
rect 31562 50713 31711 50741
rect 31562 50701 31568 50713
rect 31699 50710 31711 50713
rect 31745 50710 31757 50744
rect 31699 50704 31757 50710
rect 1152 50642 58848 50664
rect 1152 50590 4294 50642
rect 4346 50590 4358 50642
rect 4410 50590 4422 50642
rect 4474 50590 4486 50642
rect 4538 50590 35014 50642
rect 35066 50590 35078 50642
rect 35130 50590 35142 50642
rect 35194 50590 35206 50642
rect 35258 50590 58848 50642
rect 1152 50568 58848 50590
rect 23824 50479 23830 50531
rect 23882 50519 23888 50531
rect 31504 50519 31510 50531
rect 23882 50491 31510 50519
rect 23882 50479 23888 50491
rect 31504 50479 31510 50491
rect 31562 50479 31568 50531
rect 31312 50405 31318 50457
rect 31370 50445 31376 50457
rect 42256 50445 42262 50457
rect 31370 50417 42262 50445
rect 31370 50405 31376 50417
rect 42256 50405 42262 50417
rect 42314 50405 42320 50457
rect 29779 50300 29837 50306
rect 29779 50266 29791 50300
rect 29825 50297 29837 50300
rect 30067 50300 30125 50306
rect 30067 50297 30079 50300
rect 29825 50269 30079 50297
rect 29825 50266 29837 50269
rect 29779 50260 29837 50266
rect 30067 50266 30079 50269
rect 30113 50297 30125 50300
rect 56848 50297 56854 50309
rect 30113 50269 56854 50297
rect 30113 50266 30125 50269
rect 30067 50260 30125 50266
rect 56848 50257 56854 50269
rect 56906 50257 56912 50309
rect 49168 50223 49174 50235
rect 49129 50195 49174 50223
rect 49168 50183 49174 50195
rect 49226 50183 49232 50235
rect 57715 50226 57773 50232
rect 57715 50223 57727 50226
rect 57586 50195 57727 50223
rect 31792 50109 31798 50161
rect 31850 50149 31856 50161
rect 57586 50149 57614 50195
rect 57715 50192 57727 50195
rect 57761 50223 57773 50226
rect 57811 50226 57869 50232
rect 57811 50223 57823 50226
rect 57761 50195 57823 50223
rect 57761 50192 57773 50195
rect 57715 50186 57773 50192
rect 57811 50192 57823 50195
rect 57857 50192 57869 50226
rect 57811 50186 57869 50192
rect 31850 50121 57614 50149
rect 31850 50109 31856 50121
rect 49075 50078 49133 50084
rect 49075 50044 49087 50078
rect 49121 50075 49133 50078
rect 49168 50075 49174 50087
rect 49121 50047 49174 50075
rect 49121 50044 49133 50047
rect 49075 50038 49133 50044
rect 49168 50035 49174 50047
rect 49226 50035 49232 50087
rect 1152 49976 58848 49998
rect 1152 49924 19654 49976
rect 19706 49924 19718 49976
rect 19770 49924 19782 49976
rect 19834 49924 19846 49976
rect 19898 49924 50374 49976
rect 50426 49924 50438 49976
rect 50490 49924 50502 49976
rect 50554 49924 50566 49976
rect 50618 49924 58848 49976
rect 1152 49902 58848 49924
rect 38131 49412 38189 49418
rect 38131 49378 38143 49412
rect 38177 49409 38189 49412
rect 38416 49409 38422 49421
rect 38177 49381 38422 49409
rect 38177 49378 38189 49381
rect 38131 49372 38189 49378
rect 38416 49369 38422 49381
rect 38474 49369 38480 49421
rect 50323 49412 50381 49418
rect 50323 49378 50335 49412
rect 50369 49409 50381 49412
rect 50611 49412 50669 49418
rect 50611 49409 50623 49412
rect 50369 49381 50623 49409
rect 50369 49378 50381 49381
rect 50323 49372 50381 49378
rect 50611 49378 50623 49381
rect 50657 49409 50669 49412
rect 51280 49409 51286 49421
rect 50657 49381 51286 49409
rect 50657 49378 50669 49381
rect 50611 49372 50669 49378
rect 51280 49369 51286 49381
rect 51338 49369 51344 49421
rect 52048 49409 52054 49421
rect 52009 49381 52054 49409
rect 52048 49369 52054 49381
rect 52106 49369 52112 49421
rect 1152 49310 58848 49332
rect 1152 49258 4294 49310
rect 4346 49258 4358 49310
rect 4410 49258 4422 49310
rect 4474 49258 4486 49310
rect 4538 49258 35014 49310
rect 35066 49258 35078 49310
rect 35130 49258 35142 49310
rect 35194 49258 35206 49310
rect 35258 49258 58848 49310
rect 1152 49236 58848 49258
rect 40336 49147 40342 49199
rect 40394 49187 40400 49199
rect 40531 49190 40589 49196
rect 40531 49187 40543 49190
rect 40394 49159 40543 49187
rect 40394 49147 40400 49159
rect 40531 49156 40543 49159
rect 40577 49156 40589 49190
rect 40531 49150 40589 49156
rect 30928 49073 30934 49125
rect 30986 49113 30992 49125
rect 52048 49113 52054 49125
rect 30986 49085 52054 49113
rect 30986 49073 30992 49085
rect 52048 49073 52054 49085
rect 52106 49073 52112 49125
rect 38416 48999 38422 49051
rect 38474 49039 38480 49051
rect 48976 49039 48982 49051
rect 38474 49011 48982 49039
rect 38474 48999 38480 49011
rect 48976 48999 48982 49011
rect 49034 48999 49040 49051
rect 55600 48965 55606 48977
rect 27346 48937 55606 48965
rect 19123 48894 19181 48900
rect 19123 48860 19135 48894
rect 19169 48891 19181 48894
rect 19411 48894 19469 48900
rect 19411 48891 19423 48894
rect 19169 48863 19423 48891
rect 19169 48860 19181 48863
rect 19123 48854 19181 48860
rect 19411 48860 19423 48863
rect 19457 48891 19469 48894
rect 27346 48891 27374 48937
rect 55600 48925 55606 48937
rect 55658 48925 55664 48977
rect 19457 48863 27374 48891
rect 47827 48894 47885 48900
rect 19457 48860 19469 48863
rect 19411 48854 19469 48860
rect 47827 48860 47839 48894
rect 47873 48860 47885 48894
rect 47827 48854 47885 48860
rect 47842 48755 47870 48854
rect 47731 48746 47789 48752
rect 47731 48712 47743 48746
rect 47777 48743 47789 48746
rect 47824 48743 47830 48755
rect 47777 48715 47830 48743
rect 47777 48712 47789 48715
rect 47731 48706 47789 48712
rect 47824 48703 47830 48715
rect 47882 48703 47888 48755
rect 1152 48644 58848 48666
rect 1152 48592 19654 48644
rect 19706 48592 19718 48644
rect 19770 48592 19782 48644
rect 19834 48592 19846 48644
rect 19898 48592 50374 48644
rect 50426 48592 50438 48644
rect 50490 48592 50502 48644
rect 50554 48592 50566 48644
rect 50618 48592 58848 48644
rect 1152 48570 58848 48592
rect 10960 48037 10966 48089
rect 11018 48077 11024 48089
rect 54931 48080 54989 48086
rect 54931 48077 54943 48080
rect 11018 48049 54943 48077
rect 11018 48037 11024 48049
rect 54931 48046 54943 48049
rect 54977 48077 54989 48080
rect 55123 48080 55181 48086
rect 55123 48077 55135 48080
rect 54977 48049 55135 48077
rect 54977 48046 54989 48049
rect 54931 48040 54989 48046
rect 55123 48046 55135 48049
rect 55169 48046 55181 48080
rect 55123 48040 55181 48046
rect 1152 47978 58848 48000
rect 1152 47926 4294 47978
rect 4346 47926 4358 47978
rect 4410 47926 4422 47978
rect 4474 47926 4486 47978
rect 4538 47926 35014 47978
rect 35066 47926 35078 47978
rect 35130 47926 35142 47978
rect 35194 47926 35206 47978
rect 35258 47926 58848 47978
rect 1152 47904 58848 47926
rect 28720 47815 28726 47867
rect 28778 47855 28784 47867
rect 31411 47858 31469 47864
rect 31411 47855 31423 47858
rect 28778 47827 31423 47855
rect 28778 47815 28784 47827
rect 31411 47824 31423 47827
rect 31457 47824 31469 47858
rect 31411 47818 31469 47824
rect 27955 47636 28013 47642
rect 27955 47602 27967 47636
rect 28001 47633 28013 47636
rect 28243 47636 28301 47642
rect 28243 47633 28255 47636
rect 28001 47605 28255 47633
rect 28001 47602 28013 47605
rect 27955 47596 28013 47602
rect 28243 47602 28255 47605
rect 28289 47633 28301 47636
rect 34192 47633 34198 47645
rect 28289 47605 34198 47633
rect 28289 47602 28301 47605
rect 28243 47596 28301 47602
rect 34192 47593 34198 47605
rect 34250 47593 34256 47645
rect 54256 47519 54262 47571
rect 54314 47559 54320 47571
rect 54355 47562 54413 47568
rect 54355 47559 54367 47562
rect 54314 47531 54367 47559
rect 54314 47519 54320 47531
rect 54355 47528 54367 47531
rect 54401 47559 54413 47562
rect 54451 47562 54509 47568
rect 54451 47559 54463 47562
rect 54401 47531 54463 47559
rect 54401 47528 54413 47531
rect 54355 47522 54413 47528
rect 54451 47528 54463 47531
rect 54497 47528 54509 47562
rect 54451 47522 54509 47528
rect 1152 47312 58848 47334
rect 1152 47260 19654 47312
rect 19706 47260 19718 47312
rect 19770 47260 19782 47312
rect 19834 47260 19846 47312
rect 19898 47260 50374 47312
rect 50426 47260 50438 47312
rect 50490 47260 50502 47312
rect 50554 47260 50566 47312
rect 50618 47260 58848 47312
rect 1152 47238 58848 47260
rect 2608 47149 2614 47201
rect 2666 47189 2672 47201
rect 6643 47192 6701 47198
rect 6643 47189 6655 47192
rect 2666 47161 6655 47189
rect 2666 47149 2672 47161
rect 6643 47158 6655 47161
rect 6689 47158 6701 47192
rect 6643 47152 6701 47158
rect 19120 46819 19126 46831
rect 7186 46791 19126 46819
rect 2707 46748 2765 46754
rect 2707 46714 2719 46748
rect 2753 46745 2765 46748
rect 2995 46748 3053 46754
rect 2995 46745 3007 46748
rect 2753 46717 3007 46745
rect 2753 46714 2765 46717
rect 2707 46708 2765 46714
rect 2995 46714 3007 46717
rect 3041 46745 3053 46748
rect 7186 46745 7214 46791
rect 19120 46779 19126 46791
rect 19178 46779 19184 46831
rect 3041 46717 7214 46745
rect 3041 46714 3053 46717
rect 2995 46708 3053 46714
rect 10672 46705 10678 46757
rect 10730 46745 10736 46757
rect 13075 46748 13133 46754
rect 13075 46745 13087 46748
rect 10730 46717 13087 46745
rect 10730 46705 10736 46717
rect 13075 46714 13087 46717
rect 13121 46745 13133 46748
rect 13267 46748 13325 46754
rect 13267 46745 13279 46748
rect 13121 46717 13279 46745
rect 13121 46714 13133 46717
rect 13075 46708 13133 46714
rect 13267 46714 13279 46717
rect 13313 46714 13325 46748
rect 13267 46708 13325 46714
rect 1152 46646 58848 46668
rect 1152 46594 4294 46646
rect 4346 46594 4358 46646
rect 4410 46594 4422 46646
rect 4474 46594 4486 46646
rect 4538 46594 35014 46646
rect 35066 46594 35078 46646
rect 35130 46594 35142 46646
rect 35194 46594 35206 46646
rect 35258 46594 58848 46646
rect 1152 46572 58848 46594
rect 6064 46483 6070 46535
rect 6122 46523 6128 46535
rect 10672 46523 10678 46535
rect 6122 46495 10678 46523
rect 6122 46483 6128 46495
rect 10672 46483 10678 46495
rect 10730 46483 10736 46535
rect 10864 46523 10870 46535
rect 10825 46495 10870 46523
rect 10864 46483 10870 46495
rect 10922 46483 10928 46535
rect 24787 46304 24845 46310
rect 24787 46270 24799 46304
rect 24833 46301 24845 46304
rect 24833 46273 31262 46301
rect 24833 46270 24845 46273
rect 24787 46264 24845 46270
rect 27955 46230 28013 46236
rect 27955 46196 27967 46230
rect 28001 46227 28013 46230
rect 28243 46230 28301 46236
rect 28243 46227 28255 46230
rect 28001 46199 28255 46227
rect 28001 46196 28013 46199
rect 27955 46190 28013 46196
rect 28243 46196 28255 46199
rect 28289 46196 28301 46230
rect 31234 46227 31262 46273
rect 33808 46261 33814 46313
rect 33866 46301 33872 46313
rect 43699 46304 43757 46310
rect 43699 46301 43711 46304
rect 33866 46273 43711 46301
rect 33866 46261 33872 46273
rect 43699 46270 43711 46273
rect 43745 46301 43757 46304
rect 43891 46304 43949 46310
rect 43891 46301 43903 46304
rect 43745 46273 43903 46301
rect 43745 46270 43757 46273
rect 43699 46264 43757 46270
rect 43891 46270 43903 46273
rect 43937 46270 43949 46304
rect 43891 46264 43949 46270
rect 41968 46227 41974 46239
rect 31234 46199 41974 46227
rect 28243 46190 28301 46196
rect 28258 46153 28286 46190
rect 41968 46187 41974 46199
rect 42026 46187 42032 46239
rect 41104 46153 41110 46165
rect 27778 46125 27998 46153
rect 28258 46125 41110 46153
rect 7216 46039 7222 46091
rect 7274 46079 7280 46091
rect 27778 46079 27806 46125
rect 7274 46051 27806 46079
rect 27970 46079 27998 46125
rect 41104 46113 41110 46125
rect 41162 46113 41168 46165
rect 31411 46082 31469 46088
rect 31411 46079 31423 46082
rect 27970 46051 31423 46079
rect 7274 46039 7280 46051
rect 31411 46048 31423 46051
rect 31457 46048 31469 46082
rect 31411 46042 31469 46048
rect 1152 45980 58848 46002
rect 1152 45928 19654 45980
rect 19706 45928 19718 45980
rect 19770 45928 19782 45980
rect 19834 45928 19846 45980
rect 19898 45928 50374 45980
rect 50426 45928 50438 45980
rect 50490 45928 50502 45980
rect 50554 45928 50566 45980
rect 50618 45928 58848 45980
rect 1152 45906 58848 45928
rect 6259 45416 6317 45422
rect 6259 45382 6271 45416
rect 6305 45413 6317 45416
rect 6544 45413 6550 45425
rect 6305 45385 6550 45413
rect 6305 45382 6317 45385
rect 6259 45376 6317 45382
rect 6544 45373 6550 45385
rect 6602 45373 6608 45425
rect 41008 45373 41014 45425
rect 41066 45413 41072 45425
rect 41107 45416 41165 45422
rect 41107 45413 41119 45416
rect 41066 45385 41119 45413
rect 41066 45373 41072 45385
rect 41107 45382 41119 45385
rect 41153 45413 41165 45416
rect 41299 45416 41357 45422
rect 41299 45413 41311 45416
rect 41153 45385 41311 45413
rect 41153 45382 41165 45385
rect 41107 45376 41165 45382
rect 41299 45382 41311 45385
rect 41345 45382 41357 45416
rect 41299 45376 41357 45382
rect 1152 45314 58848 45336
rect 1152 45262 4294 45314
rect 4346 45262 4358 45314
rect 4410 45262 4422 45314
rect 4474 45262 4486 45314
rect 4538 45262 35014 45314
rect 35066 45262 35078 45314
rect 35130 45262 35142 45314
rect 35194 45262 35206 45314
rect 35258 45262 58848 45314
rect 1152 45240 58848 45262
rect 6544 45151 6550 45203
rect 6602 45191 6608 45203
rect 53200 45191 53206 45203
rect 6602 45163 53206 45191
rect 6602 45151 6608 45163
rect 53200 45151 53206 45163
rect 53258 45151 53264 45203
rect 44083 44898 44141 44904
rect 44083 44864 44095 44898
rect 44129 44864 44141 44898
rect 44083 44858 44141 44864
rect 47539 44898 47597 44904
rect 47539 44864 47551 44898
rect 47585 44895 47597 44898
rect 47635 44898 47693 44904
rect 47635 44895 47647 44898
rect 47585 44867 47647 44895
rect 47585 44864 47597 44867
rect 47539 44858 47597 44864
rect 47635 44864 47647 44867
rect 47681 44864 47693 44898
rect 47635 44858 47693 44864
rect 37456 44707 37462 44759
rect 37514 44747 37520 44759
rect 43891 44750 43949 44756
rect 43891 44747 43903 44750
rect 37514 44719 43903 44747
rect 37514 44707 37520 44719
rect 43891 44716 43903 44719
rect 43937 44747 43949 44750
rect 44098 44747 44126 44858
rect 43937 44719 44126 44747
rect 43937 44716 43949 44719
rect 43891 44710 43949 44716
rect 44848 44707 44854 44759
rect 44906 44747 44912 44759
rect 47554 44747 47582 44858
rect 44906 44719 47582 44747
rect 44906 44707 44912 44719
rect 1152 44648 58848 44670
rect 1152 44596 19654 44648
rect 19706 44596 19718 44648
rect 19770 44596 19782 44648
rect 19834 44596 19846 44648
rect 19898 44596 50374 44648
rect 50426 44596 50438 44648
rect 50490 44596 50502 44648
rect 50554 44596 50566 44648
rect 50618 44596 58848 44648
rect 1152 44574 58848 44596
rect 12019 44158 12077 44164
rect 12019 44124 12031 44158
rect 12065 44155 12077 44158
rect 26128 44155 26134 44167
rect 12065 44127 26134 44155
rect 12065 44124 12077 44127
rect 12019 44118 12077 44124
rect 26128 44115 26134 44127
rect 26186 44115 26192 44167
rect 17104 44081 17110 44093
rect 17017 44053 17110 44081
rect 17104 44041 17110 44053
rect 17162 44081 17168 44093
rect 17299 44084 17357 44090
rect 17299 44081 17311 44084
rect 17162 44053 17311 44081
rect 17162 44041 17168 44053
rect 17299 44050 17311 44053
rect 17345 44050 17357 44084
rect 17299 44044 17357 44050
rect 1152 43982 58848 44004
rect 1152 43930 4294 43982
rect 4346 43930 4358 43982
rect 4410 43930 4422 43982
rect 4474 43930 4486 43982
rect 4538 43930 35014 43982
rect 35066 43930 35078 43982
rect 35130 43930 35142 43982
rect 35194 43930 35206 43982
rect 35258 43930 58848 43982
rect 1152 43908 58848 43930
rect 21619 43566 21677 43572
rect 21619 43532 21631 43566
rect 21665 43532 21677 43566
rect 21619 43526 21677 43532
rect 12304 43375 12310 43427
rect 12362 43415 12368 43427
rect 21427 43418 21485 43424
rect 21427 43415 21439 43418
rect 12362 43387 21439 43415
rect 12362 43375 12368 43387
rect 21427 43384 21439 43387
rect 21473 43415 21485 43418
rect 21634 43415 21662 43526
rect 21473 43387 21662 43415
rect 21473 43384 21485 43387
rect 21427 43378 21485 43384
rect 1152 43316 58848 43338
rect 1152 43264 19654 43316
rect 19706 43264 19718 43316
rect 19770 43264 19782 43316
rect 19834 43264 19846 43316
rect 19898 43264 50374 43316
rect 50426 43264 50438 43316
rect 50490 43264 50502 43316
rect 50554 43264 50566 43316
rect 50618 43264 58848 43316
rect 1152 43242 58848 43264
rect 1840 42709 1846 42761
rect 1898 42749 1904 42761
rect 2131 42752 2189 42758
rect 2131 42749 2143 42752
rect 1898 42721 2143 42749
rect 1898 42709 1904 42721
rect 2131 42718 2143 42721
rect 2177 42749 2189 42752
rect 2323 42752 2381 42758
rect 2323 42749 2335 42752
rect 2177 42721 2335 42749
rect 2177 42718 2189 42721
rect 2131 42712 2189 42718
rect 2323 42718 2335 42721
rect 2369 42718 2381 42752
rect 2323 42712 2381 42718
rect 1152 42650 58848 42672
rect 1152 42598 4294 42650
rect 4346 42598 4358 42650
rect 4410 42598 4422 42650
rect 4474 42598 4486 42650
rect 4538 42598 35014 42650
rect 35066 42598 35078 42650
rect 35130 42598 35142 42650
rect 35194 42598 35206 42650
rect 35258 42598 58848 42650
rect 1152 42576 58848 42598
rect 33235 42234 33293 42240
rect 33235 42200 33247 42234
rect 33281 42231 33293 42234
rect 33523 42234 33581 42240
rect 33523 42231 33535 42234
rect 33281 42203 33535 42231
rect 33281 42200 33293 42203
rect 33235 42194 33293 42200
rect 33523 42200 33535 42203
rect 33569 42231 33581 42234
rect 39664 42231 39670 42243
rect 33569 42203 39670 42231
rect 33569 42200 33581 42203
rect 33523 42194 33581 42200
rect 39664 42191 39670 42203
rect 39722 42191 39728 42243
rect 46483 42234 46541 42240
rect 46483 42231 46495 42234
rect 46306 42203 46495 42231
rect 18256 42117 18262 42169
rect 18314 42157 18320 42169
rect 30931 42160 30989 42166
rect 30931 42157 30943 42160
rect 18314 42129 30943 42157
rect 18314 42117 18320 42129
rect 30931 42126 30943 42129
rect 30977 42126 30989 42160
rect 40147 42160 40205 42166
rect 40147 42157 40159 42160
rect 30931 42120 30989 42126
rect 37426 42129 40159 42157
rect 5584 42043 5590 42095
rect 5642 42083 5648 42095
rect 37426 42083 37454 42129
rect 40147 42126 40159 42129
rect 40193 42126 40205 42160
rect 40147 42120 40205 42126
rect 46306 42095 46334 42203
rect 46483 42200 46495 42203
rect 46529 42200 46541 42234
rect 46483 42194 46541 42200
rect 46288 42083 46294 42095
rect 5642 42055 37454 42083
rect 46249 42055 46294 42083
rect 5642 42043 5648 42055
rect 46288 42043 46294 42055
rect 46346 42043 46352 42095
rect 1152 41984 58848 42006
rect 1152 41932 19654 41984
rect 19706 41932 19718 41984
rect 19770 41932 19782 41984
rect 19834 41932 19846 41984
rect 19898 41932 50374 41984
rect 50426 41932 50438 41984
rect 50490 41932 50502 41984
rect 50554 41932 50566 41984
rect 50618 41932 58848 41984
rect 1152 41910 58848 41932
rect 22306 41463 27374 41491
rect 17200 41377 17206 41429
rect 17258 41417 17264 41429
rect 22306 41417 22334 41463
rect 17258 41389 22334 41417
rect 25363 41420 25421 41426
rect 17258 41377 17264 41389
rect 25363 41386 25375 41420
rect 25409 41417 25421 41420
rect 25651 41420 25709 41426
rect 25651 41417 25663 41420
rect 25409 41389 25663 41417
rect 25409 41386 25421 41389
rect 25363 41380 25421 41386
rect 25651 41386 25663 41389
rect 25697 41417 25709 41420
rect 25744 41417 25750 41429
rect 25697 41389 25750 41417
rect 25697 41386 25709 41389
rect 25651 41380 25709 41386
rect 25744 41377 25750 41389
rect 25802 41377 25808 41429
rect 27346 41417 27374 41463
rect 48307 41420 48365 41426
rect 48307 41417 48319 41420
rect 27346 41389 48319 41417
rect 48307 41386 48319 41389
rect 48353 41386 48365 41420
rect 48307 41380 48365 41386
rect 1152 41318 58848 41340
rect 1152 41266 4294 41318
rect 4346 41266 4358 41318
rect 4410 41266 4422 41318
rect 4474 41266 4486 41318
rect 4538 41266 35014 41318
rect 35066 41266 35078 41318
rect 35130 41266 35142 41318
rect 35194 41266 35206 41318
rect 35258 41266 58848 41318
rect 1152 41244 58848 41266
rect 25744 41155 25750 41207
rect 25802 41195 25808 41207
rect 46192 41195 46198 41207
rect 25802 41167 46198 41195
rect 25802 41155 25808 41167
rect 46192 41155 46198 41167
rect 46250 41155 46256 41207
rect 15379 40976 15437 40982
rect 15379 40942 15391 40976
rect 15425 40973 15437 40976
rect 15667 40976 15725 40982
rect 15667 40973 15679 40976
rect 15425 40945 15679 40973
rect 15425 40942 15437 40945
rect 15379 40936 15437 40942
rect 15667 40942 15679 40945
rect 15713 40973 15725 40976
rect 22387 40976 22445 40982
rect 22387 40973 22399 40976
rect 15713 40945 22399 40973
rect 15713 40942 15725 40945
rect 15667 40936 15725 40942
rect 22387 40942 22399 40945
rect 22433 40942 22445 40976
rect 22387 40936 22445 40942
rect 1747 40902 1805 40908
rect 1747 40868 1759 40902
rect 1793 40868 1805 40902
rect 1747 40862 1805 40868
rect 17395 40902 17453 40908
rect 17395 40868 17407 40902
rect 17441 40899 17453 40902
rect 17683 40902 17741 40908
rect 17683 40899 17695 40902
rect 17441 40871 17695 40899
rect 17441 40868 17453 40871
rect 17395 40862 17453 40868
rect 17683 40868 17695 40871
rect 17729 40899 17741 40902
rect 42736 40899 42742 40911
rect 17729 40871 42742 40899
rect 17729 40868 17741 40871
rect 17683 40862 17741 40868
rect 1762 40751 1790 40862
rect 42736 40859 42742 40871
rect 42794 40859 42800 40911
rect 22387 40828 22445 40834
rect 7186 40797 22334 40825
rect 1939 40754 1997 40760
rect 1939 40751 1951 40754
rect 1762 40723 1951 40751
rect 1939 40720 1951 40723
rect 1985 40751 1997 40754
rect 7186 40751 7214 40797
rect 1985 40723 7214 40751
rect 22306 40751 22334 40797
rect 22387 40794 22399 40828
rect 22433 40825 22445 40828
rect 29104 40825 29110 40837
rect 22433 40797 29110 40825
rect 22433 40794 22445 40797
rect 22387 40788 22445 40794
rect 29104 40785 29110 40797
rect 29162 40785 29168 40837
rect 45136 40751 45142 40763
rect 22306 40723 45142 40751
rect 1985 40720 1997 40723
rect 1939 40714 1997 40720
rect 45136 40711 45142 40723
rect 45194 40711 45200 40763
rect 1152 40652 58848 40674
rect 1152 40600 19654 40652
rect 19706 40600 19718 40652
rect 19770 40600 19782 40652
rect 19834 40600 19846 40652
rect 19898 40600 50374 40652
rect 50426 40600 50438 40652
rect 50490 40600 50502 40652
rect 50554 40600 50566 40652
rect 50618 40600 58848 40652
rect 1152 40578 58848 40600
rect 2803 40384 2861 40390
rect 2803 40350 2815 40384
rect 2849 40381 2861 40384
rect 57328 40381 57334 40393
rect 2849 40353 57334 40381
rect 2849 40350 2861 40353
rect 2803 40344 2861 40350
rect 57328 40341 57334 40353
rect 57386 40341 57392 40393
rect 32944 40085 32950 40097
rect 32905 40057 32950 40085
rect 32944 40045 32950 40057
rect 33002 40085 33008 40097
rect 33139 40088 33197 40094
rect 33139 40085 33151 40088
rect 33002 40057 33151 40085
rect 33002 40045 33008 40057
rect 33139 40054 33151 40057
rect 33185 40054 33197 40088
rect 33139 40048 33197 40054
rect 1152 39986 58848 40008
rect 1152 39934 4294 39986
rect 4346 39934 4358 39986
rect 4410 39934 4422 39986
rect 4474 39934 4486 39986
rect 4538 39934 35014 39986
rect 35066 39934 35078 39986
rect 35130 39934 35142 39986
rect 35194 39934 35206 39986
rect 35258 39934 58848 39986
rect 1152 39912 58848 39934
rect 49171 39570 49229 39576
rect 49171 39567 49183 39570
rect 48994 39539 49183 39567
rect 23920 39379 23926 39431
rect 23978 39419 23984 39431
rect 48994 39428 49022 39539
rect 49171 39536 49183 39539
rect 49217 39536 49229 39570
rect 49171 39530 49229 39536
rect 48979 39422 49037 39428
rect 48979 39419 48991 39422
rect 23978 39391 48991 39419
rect 23978 39379 23984 39391
rect 48979 39388 48991 39391
rect 49025 39388 49037 39422
rect 48979 39382 49037 39388
rect 1152 39320 58848 39342
rect 1152 39268 19654 39320
rect 19706 39268 19718 39320
rect 19770 39268 19782 39320
rect 19834 39268 19846 39320
rect 19898 39268 50374 39320
rect 50426 39268 50438 39320
rect 50490 39268 50502 39320
rect 50554 39268 50566 39320
rect 50618 39268 58848 39320
rect 1152 39246 58848 39268
rect 11152 38787 11158 38839
rect 11210 38827 11216 38839
rect 58003 38830 58061 38836
rect 58003 38827 58015 38830
rect 11210 38799 27374 38827
rect 11210 38787 11216 38799
rect 12307 38756 12365 38762
rect 12307 38722 12319 38756
rect 12353 38753 12365 38756
rect 12592 38753 12598 38765
rect 12353 38725 12598 38753
rect 12353 38722 12365 38725
rect 12307 38716 12365 38722
rect 12592 38713 12598 38725
rect 12650 38713 12656 38765
rect 24112 38753 24118 38765
rect 24073 38725 24118 38753
rect 24112 38713 24118 38725
rect 24170 38713 24176 38765
rect 27346 38753 27374 38799
rect 47506 38799 58015 38827
rect 47506 38753 47534 38799
rect 58003 38796 58015 38799
rect 58049 38796 58061 38830
rect 58003 38790 58061 38796
rect 52336 38753 52342 38765
rect 27346 38725 47534 38753
rect 52297 38725 52342 38753
rect 52336 38713 52342 38725
rect 52394 38753 52400 38765
rect 52531 38756 52589 38762
rect 52531 38753 52543 38756
rect 52394 38725 52543 38753
rect 52394 38713 52400 38725
rect 52531 38722 52543 38725
rect 52577 38722 52589 38756
rect 52531 38716 52589 38722
rect 1152 38654 58848 38676
rect 1152 38602 4294 38654
rect 4346 38602 4358 38654
rect 4410 38602 4422 38654
rect 4474 38602 4486 38654
rect 4538 38602 35014 38654
rect 35066 38602 35078 38654
rect 35130 38602 35142 38654
rect 35194 38602 35206 38654
rect 35258 38602 58848 38654
rect 1152 38580 58848 38602
rect 12592 38491 12598 38543
rect 12650 38531 12656 38543
rect 55984 38531 55990 38543
rect 12650 38503 55990 38531
rect 12650 38491 12656 38503
rect 55984 38491 55990 38503
rect 56042 38491 56048 38543
rect 11344 38417 11350 38469
rect 11402 38457 11408 38469
rect 52336 38457 52342 38469
rect 11402 38429 52342 38457
rect 11402 38417 11408 38429
rect 52336 38417 52342 38429
rect 52394 38417 52400 38469
rect 10867 38238 10925 38244
rect 10867 38204 10879 38238
rect 10913 38204 10925 38238
rect 10867 38198 10925 38204
rect 12787 38238 12845 38244
rect 12787 38204 12799 38238
rect 12833 38235 12845 38238
rect 13075 38238 13133 38244
rect 13075 38235 13087 38238
rect 12833 38207 13087 38235
rect 12833 38204 12845 38207
rect 12787 38198 12845 38204
rect 13075 38204 13087 38207
rect 13121 38235 13133 38238
rect 50224 38235 50230 38247
rect 13121 38207 50230 38235
rect 13121 38204 13133 38207
rect 13075 38198 13133 38204
rect 4048 38047 4054 38099
rect 4106 38087 4112 38099
rect 10675 38090 10733 38096
rect 10675 38087 10687 38090
rect 4106 38059 10687 38087
rect 4106 38047 4112 38059
rect 10675 38056 10687 38059
rect 10721 38087 10733 38090
rect 10882 38087 10910 38198
rect 50224 38195 50230 38207
rect 50282 38195 50288 38247
rect 10721 38059 10910 38087
rect 10721 38056 10733 38059
rect 10675 38050 10733 38056
rect 1152 37988 58848 38010
rect 1152 37936 19654 37988
rect 19706 37936 19718 37988
rect 19770 37936 19782 37988
rect 19834 37936 19846 37988
rect 19898 37936 50374 37988
rect 50426 37936 50438 37988
rect 50490 37936 50502 37988
rect 50554 37936 50566 37988
rect 50618 37936 58848 37988
rect 1152 37914 58848 37936
rect 10003 37572 10061 37578
rect 10003 37538 10015 37572
rect 10049 37569 10061 37572
rect 10049 37541 10142 37569
rect 10049 37538 10061 37541
rect 10003 37532 10061 37538
rect 10114 37421 10142 37541
rect 10291 37424 10349 37430
rect 10291 37421 10303 37424
rect 10114 37393 10303 37421
rect 10291 37390 10303 37393
rect 10337 37421 10349 37424
rect 11152 37421 11158 37433
rect 10337 37393 11158 37421
rect 10337 37390 10349 37393
rect 10291 37384 10349 37390
rect 11152 37381 11158 37393
rect 11210 37381 11216 37433
rect 11443 37424 11501 37430
rect 11443 37390 11455 37424
rect 11489 37421 11501 37424
rect 20272 37421 20278 37433
rect 11489 37393 20278 37421
rect 11489 37390 11501 37393
rect 11443 37384 11501 37390
rect 20272 37381 20278 37393
rect 20330 37381 20336 37433
rect 29491 37424 29549 37430
rect 29491 37390 29503 37424
rect 29537 37421 29549 37424
rect 29584 37421 29590 37433
rect 29537 37393 29590 37421
rect 29537 37390 29549 37393
rect 29491 37384 29549 37390
rect 29584 37381 29590 37393
rect 29642 37381 29648 37433
rect 1152 37322 58848 37344
rect 1152 37270 4294 37322
rect 4346 37270 4358 37322
rect 4410 37270 4422 37322
rect 4474 37270 4486 37322
rect 4538 37270 35014 37322
rect 35066 37270 35078 37322
rect 35130 37270 35142 37322
rect 35194 37270 35206 37322
rect 35258 37270 58848 37322
rect 1152 37248 58848 37270
rect 5008 37199 5014 37211
rect 4969 37171 5014 37199
rect 5008 37159 5014 37171
rect 5066 37159 5072 37211
rect 11152 37159 11158 37211
rect 11210 37199 11216 37211
rect 30256 37199 30262 37211
rect 11210 37171 30262 37199
rect 11210 37159 11216 37171
rect 30256 37159 30262 37171
rect 30314 37159 30320 37211
rect 33811 36906 33869 36912
rect 33811 36872 33823 36906
rect 33857 36903 33869 36906
rect 34099 36906 34157 36912
rect 34099 36903 34111 36906
rect 33857 36875 34111 36903
rect 33857 36872 33869 36875
rect 33811 36866 33869 36872
rect 34099 36872 34111 36875
rect 34145 36903 34157 36906
rect 51760 36903 51766 36915
rect 34145 36875 51766 36903
rect 34145 36872 34157 36875
rect 34099 36866 34157 36872
rect 51760 36863 51766 36875
rect 51818 36863 51824 36915
rect 1152 36656 58848 36678
rect 1152 36604 19654 36656
rect 19706 36604 19718 36656
rect 19770 36604 19782 36656
rect 19834 36604 19846 36656
rect 19898 36604 50374 36656
rect 50426 36604 50438 36656
rect 50490 36604 50502 36656
rect 50554 36604 50566 36656
rect 50618 36604 58848 36656
rect 1152 36582 58848 36604
rect 2419 36536 2477 36542
rect 2419 36502 2431 36536
rect 2465 36533 2477 36536
rect 2800 36533 2806 36545
rect 2465 36505 2806 36533
rect 2465 36502 2477 36505
rect 2419 36496 2477 36502
rect 2800 36493 2806 36505
rect 2858 36493 2864 36545
rect 7315 36166 7373 36172
rect 7315 36132 7327 36166
rect 7361 36163 7373 36166
rect 7361 36135 17294 36163
rect 7361 36132 7373 36135
rect 7315 36126 7373 36132
rect 16432 36089 16438 36101
rect 16393 36061 16438 36089
rect 16432 36049 16438 36061
rect 16490 36089 16496 36101
rect 16819 36092 16877 36098
rect 16819 36089 16831 36092
rect 16490 36061 16831 36089
rect 16490 36049 16496 36061
rect 16819 36058 16831 36061
rect 16865 36058 16877 36092
rect 17266 36089 17294 36135
rect 56272 36089 56278 36101
rect 17266 36061 56278 36089
rect 16819 36052 16877 36058
rect 56272 36049 56278 36061
rect 56330 36049 56336 36101
rect 1152 35990 58848 36012
rect 1152 35938 4294 35990
rect 4346 35938 4358 35990
rect 4410 35938 4422 35990
rect 4474 35938 4486 35990
rect 4538 35938 35014 35990
rect 35066 35938 35078 35990
rect 35130 35938 35142 35990
rect 35194 35938 35206 35990
rect 35258 35938 58848 35990
rect 1152 35916 58848 35938
rect 13072 35531 13078 35583
rect 13130 35571 13136 35583
rect 13267 35574 13325 35580
rect 13267 35571 13279 35574
rect 13130 35543 13279 35571
rect 13130 35531 13136 35543
rect 13267 35540 13279 35543
rect 13313 35540 13325 35574
rect 13267 35534 13325 35540
rect 22960 35531 22966 35583
rect 23018 35571 23024 35583
rect 39091 35574 39149 35580
rect 39091 35571 39103 35574
rect 23018 35543 39103 35571
rect 23018 35531 23024 35543
rect 39091 35540 39103 35543
rect 39137 35540 39149 35574
rect 39091 35534 39149 35540
rect 43891 35574 43949 35580
rect 43891 35540 43903 35574
rect 43937 35540 43949 35574
rect 43891 35534 43949 35540
rect 7186 35469 17294 35497
rect 5296 35383 5302 35435
rect 5354 35423 5360 35435
rect 7186 35423 7214 35469
rect 13072 35423 13078 35435
rect 5354 35395 7214 35423
rect 13033 35395 13078 35423
rect 5354 35383 5360 35395
rect 13072 35383 13078 35395
rect 13130 35383 13136 35435
rect 17266 35423 17294 35469
rect 43699 35426 43757 35432
rect 43699 35423 43711 35426
rect 17266 35395 43711 35423
rect 43699 35392 43711 35395
rect 43745 35423 43757 35426
rect 43906 35423 43934 35534
rect 43745 35395 43934 35423
rect 43745 35392 43757 35395
rect 43699 35386 43757 35392
rect 1152 35324 58848 35346
rect 1152 35272 19654 35324
rect 19706 35272 19718 35324
rect 19770 35272 19782 35324
rect 19834 35272 19846 35324
rect 19898 35272 50374 35324
rect 50426 35272 50438 35324
rect 50490 35272 50502 35324
rect 50554 35272 50566 35324
rect 50618 35272 58848 35324
rect 1152 35250 58848 35272
rect 32464 35013 32470 35065
rect 32522 35053 32528 35065
rect 33139 35056 33197 35062
rect 33139 35053 33151 35056
rect 32522 35025 33151 35053
rect 32522 35013 32528 35025
rect 33139 35022 33151 35025
rect 33185 35022 33197 35056
rect 33139 35016 33197 35022
rect 22288 34865 22294 34917
rect 22346 34905 22352 34917
rect 51667 34908 51725 34914
rect 51667 34905 51679 34908
rect 22346 34877 51679 34905
rect 22346 34865 22352 34877
rect 51667 34874 51679 34877
rect 51713 34905 51725 34908
rect 51859 34908 51917 34914
rect 51859 34905 51871 34908
rect 51713 34877 51871 34905
rect 51713 34874 51725 34877
rect 51667 34868 51725 34874
rect 51859 34874 51871 34877
rect 51905 34874 51917 34908
rect 51859 34868 51917 34874
rect 6067 34834 6125 34840
rect 6067 34800 6079 34834
rect 6113 34831 6125 34834
rect 12688 34831 12694 34843
rect 6113 34803 12694 34831
rect 6113 34800 6125 34803
rect 6067 34794 6125 34800
rect 12688 34791 12694 34803
rect 12746 34791 12752 34843
rect 22771 34834 22829 34840
rect 22771 34831 22783 34834
rect 17266 34803 22783 34831
rect 12592 34717 12598 34769
rect 12650 34757 12656 34769
rect 17266 34757 17294 34803
rect 22771 34800 22783 34803
rect 22817 34831 22829 34834
rect 22963 34834 23021 34840
rect 22963 34831 22975 34834
rect 22817 34803 22975 34831
rect 22817 34800 22829 34803
rect 22771 34794 22829 34800
rect 22963 34800 22975 34803
rect 23009 34800 23021 34834
rect 36592 34831 36598 34843
rect 22963 34794 23021 34800
rect 27346 34803 36598 34831
rect 12650 34729 17294 34757
rect 21043 34760 21101 34766
rect 12650 34717 12656 34729
rect 21043 34726 21055 34760
rect 21089 34757 21101 34760
rect 21331 34760 21389 34766
rect 21331 34757 21343 34760
rect 21089 34729 21343 34757
rect 21089 34726 21101 34729
rect 21043 34720 21101 34726
rect 21331 34726 21343 34729
rect 21377 34757 21389 34760
rect 27346 34757 27374 34803
rect 36592 34791 36598 34803
rect 36650 34791 36656 34843
rect 43408 34791 43414 34843
rect 43466 34831 43472 34843
rect 52339 34834 52397 34840
rect 52339 34831 52351 34834
rect 43466 34803 52351 34831
rect 43466 34791 43472 34803
rect 52339 34800 52351 34803
rect 52385 34831 52397 34834
rect 52531 34834 52589 34840
rect 52531 34831 52543 34834
rect 52385 34803 52543 34831
rect 52385 34800 52397 34803
rect 52339 34794 52397 34800
rect 52531 34800 52543 34803
rect 52577 34800 52589 34834
rect 52531 34794 52589 34800
rect 28528 34757 28534 34769
rect 21377 34729 27374 34757
rect 28489 34729 28534 34757
rect 21377 34726 21389 34729
rect 21331 34720 21389 34726
rect 28528 34717 28534 34729
rect 28586 34757 28592 34769
rect 28723 34760 28781 34766
rect 28723 34757 28735 34760
rect 28586 34729 28735 34757
rect 28586 34717 28592 34729
rect 28723 34726 28735 34729
rect 28769 34726 28781 34760
rect 28723 34720 28781 34726
rect 1152 34658 58848 34680
rect 1152 34606 4294 34658
rect 4346 34606 4358 34658
rect 4410 34606 4422 34658
rect 4474 34606 4486 34658
rect 4538 34606 35014 34658
rect 35066 34606 35078 34658
rect 35130 34606 35142 34658
rect 35194 34606 35206 34658
rect 35258 34606 58848 34658
rect 1152 34584 58848 34606
rect 22960 34239 22966 34251
rect 22921 34211 22966 34239
rect 22960 34199 22966 34211
rect 23018 34199 23024 34251
rect 55795 34242 55853 34248
rect 55795 34208 55807 34242
rect 55841 34239 55853 34242
rect 56944 34239 56950 34251
rect 55841 34211 56950 34239
rect 55841 34208 55853 34211
rect 55795 34202 55853 34208
rect 56944 34199 56950 34211
rect 57002 34199 57008 34251
rect 1152 33992 58848 34014
rect 1152 33940 19654 33992
rect 19706 33940 19718 33992
rect 19770 33940 19782 33992
rect 19834 33940 19846 33992
rect 19898 33940 50374 33992
rect 50426 33940 50438 33992
rect 50490 33940 50502 33992
rect 50554 33940 50566 33992
rect 50618 33940 58848 33992
rect 1152 33918 58848 33940
rect 34576 33607 34582 33659
rect 34634 33647 34640 33659
rect 34634 33619 52574 33647
rect 34634 33607 34640 33619
rect 12496 33533 12502 33585
rect 12554 33573 12560 33585
rect 28147 33576 28205 33582
rect 28147 33573 28159 33576
rect 12554 33545 28159 33573
rect 12554 33533 12560 33545
rect 28147 33542 28159 33545
rect 28193 33573 28205 33576
rect 28339 33576 28397 33582
rect 28339 33573 28351 33576
rect 28193 33545 28351 33573
rect 28193 33542 28205 33545
rect 28147 33536 28205 33542
rect 28339 33542 28351 33545
rect 28385 33542 28397 33576
rect 48208 33573 48214 33585
rect 28339 33536 28397 33542
rect 42370 33545 48214 33573
rect 27346 33471 37454 33499
rect 15952 33385 15958 33437
rect 16010 33425 16016 33437
rect 17107 33428 17165 33434
rect 17107 33425 17119 33428
rect 16010 33397 17119 33425
rect 16010 33385 16016 33397
rect 17107 33394 17119 33397
rect 17153 33425 17165 33428
rect 17299 33428 17357 33434
rect 17299 33425 17311 33428
rect 17153 33397 17311 33425
rect 17153 33394 17165 33397
rect 17107 33388 17165 33394
rect 17299 33394 17311 33397
rect 17345 33394 17357 33428
rect 17299 33388 17357 33394
rect 18739 33428 18797 33434
rect 18739 33394 18751 33428
rect 18785 33425 18797 33428
rect 27346 33425 27374 33471
rect 18785 33397 27374 33425
rect 37426 33425 37454 33471
rect 42370 33425 42398 33545
rect 48208 33533 48214 33545
rect 48266 33533 48272 33585
rect 52546 33499 52574 33619
rect 57619 33502 57677 33508
rect 57619 33499 57631 33502
rect 52546 33471 57631 33499
rect 57619 33468 57631 33471
rect 57665 33468 57677 33502
rect 57619 33462 57677 33468
rect 43120 33425 43126 33437
rect 37426 33397 42398 33425
rect 43081 33397 43126 33425
rect 18785 33394 18797 33397
rect 18739 33388 18797 33394
rect 43120 33385 43126 33397
rect 43178 33385 43184 33437
rect 1152 33326 58848 33348
rect 1152 33274 4294 33326
rect 4346 33274 4358 33326
rect 4410 33274 4422 33326
rect 4474 33274 4486 33326
rect 4538 33274 35014 33326
rect 35066 33274 35078 33326
rect 35130 33274 35142 33326
rect 35194 33274 35206 33326
rect 35258 33274 58848 33326
rect 1152 33252 58848 33274
rect 13744 33163 13750 33215
rect 13802 33203 13808 33215
rect 43120 33203 43126 33215
rect 13802 33175 43126 33203
rect 13802 33163 13808 33175
rect 43120 33163 43126 33175
rect 43178 33163 43184 33215
rect 44755 33206 44813 33212
rect 44755 33172 44767 33206
rect 44801 33203 44813 33206
rect 49648 33203 49654 33215
rect 44801 33175 49654 33203
rect 44801 33172 44813 33175
rect 44755 33166 44813 33172
rect 49648 33163 49654 33175
rect 49706 33163 49712 33215
rect 2515 33058 2573 33064
rect 2515 33024 2527 33058
rect 2561 33055 2573 33058
rect 2704 33055 2710 33067
rect 2561 33027 2710 33055
rect 2561 33024 2573 33027
rect 2515 33018 2573 33024
rect 2704 33015 2710 33027
rect 2762 33015 2768 33067
rect 29488 32941 29494 32993
rect 29546 32981 29552 32993
rect 46771 32984 46829 32990
rect 46771 32981 46783 32984
rect 29546 32953 46783 32981
rect 29546 32941 29552 32953
rect 46771 32950 46783 32953
rect 46817 32981 46829 32984
rect 46963 32984 47021 32990
rect 46963 32981 46975 32984
rect 46817 32953 46975 32981
rect 46817 32950 46829 32953
rect 46771 32944 46829 32950
rect 46963 32950 46975 32953
rect 47009 32950 47021 32984
rect 46963 32944 47021 32950
rect 40051 32910 40109 32916
rect 40051 32876 40063 32910
rect 40097 32876 40109 32910
rect 40051 32870 40109 32876
rect 33232 32719 33238 32771
rect 33290 32759 33296 32771
rect 39859 32762 39917 32768
rect 39859 32759 39871 32762
rect 33290 32731 39871 32759
rect 33290 32719 33296 32731
rect 39859 32728 39871 32731
rect 39905 32759 39917 32762
rect 40066 32759 40094 32870
rect 39905 32731 40094 32759
rect 39905 32728 39917 32731
rect 39859 32722 39917 32728
rect 1152 32660 58848 32682
rect 1152 32608 19654 32660
rect 19706 32608 19718 32660
rect 19770 32608 19782 32660
rect 19834 32608 19846 32660
rect 19898 32608 50374 32660
rect 50426 32608 50438 32660
rect 50490 32608 50502 32660
rect 50554 32608 50566 32660
rect 50618 32608 58848 32660
rect 1152 32586 58848 32608
rect 8467 32170 8525 32176
rect 8467 32136 8479 32170
rect 8513 32167 8525 32170
rect 53680 32167 53686 32179
rect 8513 32139 53686 32167
rect 8513 32136 8525 32139
rect 8467 32130 8525 32136
rect 53680 32127 53686 32139
rect 53738 32127 53744 32179
rect 32176 32093 32182 32105
rect 32137 32065 32182 32093
rect 32176 32053 32182 32065
rect 32234 32053 32240 32105
rect 39280 32053 39286 32105
rect 39338 32093 39344 32105
rect 43027 32096 43085 32102
rect 43027 32093 43039 32096
rect 39338 32065 43039 32093
rect 39338 32053 39344 32065
rect 43027 32062 43039 32065
rect 43073 32062 43085 32096
rect 43027 32056 43085 32062
rect 1152 31994 58848 32016
rect 1152 31942 4294 31994
rect 4346 31942 4358 31994
rect 4410 31942 4422 31994
rect 4474 31942 4486 31994
rect 4538 31942 35014 31994
rect 35066 31942 35078 31994
rect 35130 31942 35142 31994
rect 35194 31942 35206 31994
rect 35258 31942 58848 31994
rect 1152 31920 58848 31942
rect 32176 31831 32182 31883
rect 32234 31871 32240 31883
rect 52048 31871 52054 31883
rect 32234 31843 52054 31871
rect 32234 31831 32240 31843
rect 52048 31831 52054 31843
rect 52106 31831 52112 31883
rect 21232 31683 21238 31735
rect 21290 31723 21296 31735
rect 21331 31726 21389 31732
rect 21331 31723 21343 31726
rect 21290 31695 21343 31723
rect 21290 31683 21296 31695
rect 21331 31692 21343 31695
rect 21377 31692 21389 31726
rect 21331 31686 21389 31692
rect 34675 31726 34733 31732
rect 34675 31692 34687 31726
rect 34721 31723 34733 31726
rect 36112 31723 36118 31735
rect 34721 31695 36118 31723
rect 34721 31692 34733 31695
rect 34675 31686 34733 31692
rect 36112 31683 36118 31695
rect 36170 31683 36176 31735
rect 20368 31609 20374 31661
rect 20426 31649 20432 31661
rect 29011 31652 29069 31658
rect 29011 31649 29023 31652
rect 20426 31621 29023 31649
rect 20426 31609 20432 31621
rect 29011 31618 29023 31621
rect 29057 31618 29069 31652
rect 29011 31612 29069 31618
rect 1152 31328 58848 31350
rect 1152 31276 19654 31328
rect 19706 31276 19718 31328
rect 19770 31276 19782 31328
rect 19834 31276 19846 31328
rect 19898 31276 50374 31328
rect 50426 31276 50438 31328
rect 50490 31276 50502 31328
rect 50554 31276 50566 31328
rect 50618 31276 58848 31328
rect 1152 31254 58848 31276
rect 54544 31017 54550 31069
rect 54602 31057 54608 31069
rect 54739 31060 54797 31066
rect 54739 31057 54751 31060
rect 54602 31029 54751 31057
rect 54602 31017 54608 31029
rect 54739 31026 54751 31029
rect 54785 31026 54797 31060
rect 54739 31020 54797 31026
rect 7987 30764 8045 30770
rect 7987 30730 7999 30764
rect 8033 30761 8045 30764
rect 8275 30764 8333 30770
rect 8275 30761 8287 30764
rect 8033 30733 8287 30761
rect 8033 30730 8045 30733
rect 7987 30724 8045 30730
rect 8275 30730 8287 30733
rect 8321 30761 8333 30764
rect 35440 30761 35446 30773
rect 8321 30733 35446 30761
rect 8321 30730 8333 30733
rect 8275 30724 8333 30730
rect 35440 30721 35446 30733
rect 35498 30721 35504 30773
rect 1152 30662 58848 30684
rect 1152 30610 4294 30662
rect 4346 30610 4358 30662
rect 4410 30610 4422 30662
rect 4474 30610 4486 30662
rect 4538 30610 35014 30662
rect 35066 30610 35078 30662
rect 35130 30610 35142 30662
rect 35194 30610 35206 30662
rect 35258 30610 58848 30662
rect 1152 30588 58848 30610
rect 16147 30320 16205 30326
rect 16147 30286 16159 30320
rect 16193 30317 16205 30320
rect 16240 30317 16246 30329
rect 16193 30289 16246 30317
rect 16193 30286 16205 30289
rect 16147 30280 16205 30286
rect 16240 30277 16246 30289
rect 16298 30277 16304 30329
rect 1152 29996 58848 30018
rect 1152 29944 19654 29996
rect 19706 29944 19718 29996
rect 19770 29944 19782 29996
rect 19834 29944 19846 29996
rect 19898 29944 50374 29996
rect 50426 29944 50438 29996
rect 50490 29944 50502 29996
rect 50554 29944 50566 29996
rect 50618 29944 58848 29996
rect 1152 29922 58848 29944
rect 5779 29654 5837 29660
rect 5779 29620 5791 29654
rect 5825 29651 5837 29654
rect 6067 29654 6125 29660
rect 6067 29651 6079 29654
rect 5825 29623 6079 29651
rect 5825 29620 5837 29623
rect 5779 29614 5837 29620
rect 6067 29620 6079 29623
rect 6113 29651 6125 29654
rect 13264 29651 13270 29663
rect 6113 29623 13270 29651
rect 6113 29620 6125 29623
rect 6067 29614 6125 29620
rect 13264 29611 13270 29623
rect 13322 29611 13328 29663
rect 8656 29537 8662 29589
rect 8714 29577 8720 29589
rect 18832 29577 18838 29589
rect 8714 29549 18838 29577
rect 8714 29537 8720 29549
rect 18832 29537 18838 29549
rect 18890 29537 18896 29589
rect 8272 29463 8278 29515
rect 8330 29503 8336 29515
rect 17872 29503 17878 29515
rect 8330 29475 17878 29503
rect 8330 29463 8336 29475
rect 17872 29463 17878 29475
rect 17930 29463 17936 29515
rect 18352 29429 18358 29441
rect 18313 29401 18358 29429
rect 18352 29389 18358 29401
rect 18410 29389 18416 29441
rect 1152 29330 58848 29352
rect 1152 29278 4294 29330
rect 4346 29278 4358 29330
rect 4410 29278 4422 29330
rect 4474 29278 4486 29330
rect 4538 29278 35014 29330
rect 35066 29278 35078 29330
rect 35130 29278 35142 29330
rect 35194 29278 35206 29330
rect 35258 29278 58848 29330
rect 1152 29256 58848 29278
rect 8230 28923 8282 28929
rect 8674 28923 8702 29024
rect 8656 28871 8662 28923
rect 8714 28871 8720 28923
rect 8230 28865 8282 28871
rect 10096 28797 10102 28849
rect 10154 28837 10160 28849
rect 47347 28840 47405 28846
rect 10154 28809 46142 28837
rect 10154 28797 10160 28809
rect 8609 28723 8615 28775
rect 8667 28723 8673 28775
rect 46114 28763 46142 28809
rect 47347 28806 47359 28840
rect 47393 28806 47405 28840
rect 47347 28800 47405 28806
rect 47362 28763 47390 28800
rect 47539 28766 47597 28772
rect 47539 28763 47551 28766
rect 46114 28735 47551 28763
rect 47539 28732 47551 28735
rect 47585 28732 47597 28766
rect 47539 28726 47597 28732
rect 1152 28664 58848 28686
rect 1152 28612 19654 28664
rect 19706 28612 19718 28664
rect 19770 28612 19782 28664
rect 19834 28612 19846 28664
rect 19898 28612 50374 28664
rect 50426 28612 50438 28664
rect 50490 28612 50502 28664
rect 50554 28612 50566 28664
rect 50618 28612 58848 28664
rect 1152 28590 58848 28612
rect 8609 28501 8615 28553
rect 8667 28541 8673 28553
rect 18928 28541 18934 28553
rect 8667 28513 18934 28541
rect 8667 28501 8673 28513
rect 18928 28501 18934 28513
rect 18986 28501 18992 28553
rect 5968 28279 5974 28331
rect 6026 28319 6032 28331
rect 14416 28319 14422 28331
rect 6026 28291 14422 28319
rect 6026 28279 6032 28291
rect 14416 28279 14422 28291
rect 14474 28279 14480 28331
rect 3280 28205 3286 28257
rect 3338 28245 3344 28257
rect 31027 28248 31085 28254
rect 31027 28245 31039 28248
rect 3338 28217 31039 28245
rect 3338 28205 3344 28217
rect 31027 28214 31039 28217
rect 31073 28245 31085 28248
rect 31219 28248 31277 28254
rect 31219 28245 31231 28248
rect 31073 28217 31231 28245
rect 31073 28214 31085 28217
rect 31027 28208 31085 28214
rect 31219 28214 31231 28217
rect 31265 28214 31277 28248
rect 31219 28208 31277 28214
rect 8176 28131 8182 28183
rect 8234 28171 8240 28183
rect 18064 28171 18070 28183
rect 8234 28143 18070 28171
rect 8234 28131 8240 28143
rect 18064 28131 18070 28143
rect 18122 28131 18128 28183
rect 6544 28057 6550 28109
rect 6602 28097 6608 28109
rect 9907 28100 9965 28106
rect 9907 28097 9919 28100
rect 6602 28069 9919 28097
rect 6602 28057 6608 28069
rect 9907 28066 9919 28069
rect 9953 28066 9965 28100
rect 21328 28097 21334 28109
rect 21289 28069 21334 28097
rect 9907 28060 9965 28066
rect 21328 28057 21334 28069
rect 21386 28057 21392 28109
rect 29008 28057 29014 28109
rect 29066 28097 29072 28109
rect 57331 28100 57389 28106
rect 57331 28097 57343 28100
rect 29066 28069 57343 28097
rect 29066 28057 29072 28069
rect 57331 28066 57343 28069
rect 57377 28066 57389 28100
rect 57331 28060 57389 28066
rect 1152 27998 58848 28020
rect 1152 27946 4294 27998
rect 4346 27946 4358 27998
rect 4410 27946 4422 27998
rect 4474 27946 4486 27998
rect 4538 27946 35014 27998
rect 35066 27946 35078 27998
rect 35130 27946 35142 27998
rect 35194 27946 35206 27998
rect 35258 27946 58848 27998
rect 1152 27924 58848 27946
rect 9328 27835 9334 27887
rect 9386 27875 9392 27887
rect 12688 27875 12694 27887
rect 9386 27847 12694 27875
rect 9386 27835 9392 27847
rect 12688 27835 12694 27847
rect 12746 27835 12752 27887
rect 14416 27875 14422 27887
rect 14377 27847 14422 27875
rect 14416 27835 14422 27847
rect 14474 27875 14480 27887
rect 14611 27878 14669 27884
rect 14611 27875 14623 27878
rect 14474 27847 14623 27875
rect 14474 27835 14480 27847
rect 14611 27844 14623 27847
rect 14657 27844 14669 27878
rect 14611 27838 14669 27844
rect 21328 27835 21334 27887
rect 21386 27875 21392 27887
rect 48112 27875 48118 27887
rect 21386 27847 48118 27875
rect 21386 27835 21392 27847
rect 48112 27835 48118 27847
rect 48170 27835 48176 27887
rect 5299 27582 5357 27588
rect 5299 27548 5311 27582
rect 5345 27579 5357 27582
rect 5392 27579 5398 27591
rect 5345 27551 5398 27579
rect 5345 27548 5357 27551
rect 5299 27542 5357 27548
rect 5392 27539 5398 27551
rect 5450 27539 5456 27591
rect 26224 27539 26230 27591
rect 26282 27579 26288 27591
rect 57715 27582 57773 27588
rect 57715 27579 57727 27582
rect 26282 27551 57727 27579
rect 26282 27539 26288 27551
rect 57715 27548 57727 27551
rect 57761 27548 57773 27582
rect 57715 27542 57773 27548
rect 8176 27465 8182 27517
rect 8234 27465 8240 27517
rect 9328 27465 9334 27517
rect 9386 27465 9392 27517
rect 9040 27431 9046 27443
rect 8641 27403 9046 27431
rect 9040 27391 9046 27403
rect 9098 27391 9104 27443
rect 9616 27391 9622 27443
rect 9674 27431 9680 27443
rect 16816 27431 16822 27443
rect 9674 27403 16822 27431
rect 9674 27391 9680 27403
rect 16816 27391 16822 27403
rect 16874 27391 16880 27443
rect 1152 27332 58848 27354
rect 1152 27280 19654 27332
rect 19706 27280 19718 27332
rect 19770 27280 19782 27332
rect 19834 27280 19846 27332
rect 19898 27280 50374 27332
rect 50426 27280 50438 27332
rect 50490 27280 50502 27332
rect 50554 27280 50566 27332
rect 50618 27280 58848 27332
rect 1152 27258 58848 27280
rect 31696 27169 31702 27221
rect 31754 27209 31760 27221
rect 38611 27212 38669 27218
rect 38611 27209 38623 27212
rect 31754 27181 38623 27209
rect 31754 27169 31760 27181
rect 38611 27178 38623 27181
rect 38657 27178 38669 27212
rect 38611 27172 38669 27178
rect 38626 27061 38654 27172
rect 38803 27064 38861 27070
rect 38803 27061 38815 27064
rect 38626 27033 38815 27061
rect 38803 27030 38815 27033
rect 38849 27030 38861 27064
rect 38803 27024 38861 27030
rect 1936 26873 1942 26925
rect 1994 26913 2000 26925
rect 34864 26913 34870 26925
rect 1994 26885 34870 26913
rect 1994 26873 2000 26885
rect 34864 26873 34870 26885
rect 34922 26873 34928 26925
rect 18160 26799 18166 26851
rect 18218 26839 18224 26851
rect 42259 26842 42317 26848
rect 42259 26839 42271 26842
rect 18218 26811 42271 26839
rect 18218 26799 18224 26811
rect 42259 26808 42271 26811
rect 42305 26808 42317 26842
rect 42259 26802 42317 26808
rect 15091 26768 15149 26774
rect 15091 26734 15103 26768
rect 15137 26765 15149 26768
rect 26416 26765 26422 26777
rect 15137 26737 26422 26765
rect 15137 26734 15149 26737
rect 15091 26728 15149 26734
rect 26416 26725 26422 26737
rect 26474 26725 26480 26777
rect 36208 26765 36214 26777
rect 36169 26737 36214 26765
rect 36208 26725 36214 26737
rect 36266 26725 36272 26777
rect 1152 26666 58848 26688
rect 1152 26614 4294 26666
rect 4346 26614 4358 26666
rect 4410 26614 4422 26666
rect 4474 26614 4486 26666
rect 4538 26614 35014 26666
rect 35066 26614 35078 26666
rect 35130 26614 35142 26666
rect 35194 26614 35206 26666
rect 35258 26614 58848 26666
rect 1152 26592 58848 26614
rect 1936 26543 1942 26555
rect 1897 26515 1942 26543
rect 1936 26503 1942 26515
rect 1994 26503 2000 26555
rect 10864 26543 10870 26555
rect 8530 26515 10870 26543
rect 8530 26469 8558 26515
rect 10864 26503 10870 26515
rect 10922 26503 10928 26555
rect 7954 26441 8558 26469
rect 8755 26472 8813 26478
rect 7954 26381 7982 26441
rect 8755 26438 8767 26472
rect 8801 26469 8813 26472
rect 12112 26469 12118 26481
rect 8801 26441 12118 26469
rect 8801 26438 8813 26441
rect 8755 26432 8813 26438
rect 12112 26429 12118 26441
rect 12170 26429 12176 26481
rect 8371 26398 8429 26404
rect 8371 26395 8383 26398
rect 8256 26367 8383 26395
rect 8371 26364 8383 26367
rect 8417 26364 8429 26398
rect 8371 26358 8429 26364
rect 37744 26207 37750 26259
rect 37802 26247 37808 26259
rect 57715 26250 57773 26256
rect 57715 26247 57727 26250
rect 37802 26219 57727 26247
rect 37802 26207 37808 26219
rect 57715 26216 57727 26219
rect 57761 26247 57773 26250
rect 57811 26250 57869 26256
rect 57811 26247 57823 26250
rect 57761 26219 57823 26247
rect 57761 26216 57773 26219
rect 57715 26210 57773 26216
rect 57811 26216 57823 26219
rect 57857 26216 57869 26250
rect 57811 26210 57869 26216
rect 17008 26099 17014 26111
rect 8640 26071 17014 26099
rect 17008 26059 17014 26071
rect 17066 26059 17072 26111
rect 1152 26000 58848 26022
rect 1152 25948 19654 26000
rect 19706 25948 19718 26000
rect 19770 25948 19782 26000
rect 19834 25948 19846 26000
rect 19898 25948 50374 26000
rect 50426 25948 50438 26000
rect 50490 25948 50502 26000
rect 50554 25948 50566 26000
rect 50618 25948 58848 26000
rect 1152 25926 58848 25948
rect 25363 25584 25421 25590
rect 25363 25550 25375 25584
rect 25409 25581 25421 25584
rect 25651 25584 25709 25590
rect 25651 25581 25663 25584
rect 25409 25553 25663 25581
rect 25409 25550 25421 25553
rect 25363 25544 25421 25550
rect 25651 25550 25663 25553
rect 25697 25581 25709 25584
rect 40720 25581 40726 25593
rect 25697 25553 40726 25581
rect 25697 25550 25709 25553
rect 25651 25544 25709 25550
rect 40720 25541 40726 25553
rect 40778 25541 40784 25593
rect 12016 25467 12022 25519
rect 12074 25507 12080 25519
rect 33523 25510 33581 25516
rect 33523 25507 33535 25510
rect 12074 25479 33535 25507
rect 12074 25467 12080 25479
rect 33523 25476 33535 25479
rect 33569 25476 33581 25510
rect 33523 25470 33581 25476
rect 1152 25334 58848 25356
rect 1152 25282 4294 25334
rect 4346 25282 4358 25334
rect 4410 25282 4422 25334
rect 4474 25282 4486 25334
rect 4538 25282 35014 25334
rect 35066 25282 35078 25334
rect 35130 25282 35142 25334
rect 35194 25282 35206 25334
rect 35258 25282 58848 25334
rect 1152 25260 58848 25282
rect 11056 25211 11062 25223
rect 8530 25183 11062 25211
rect 8530 25137 8558 25183
rect 11056 25171 11062 25183
rect 11114 25171 11120 25223
rect 7954 25109 8558 25137
rect 7954 25049 7982 25109
rect 8098 25035 8256 25063
rect 8098 25001 8126 25035
rect 8080 24949 8086 25001
rect 8138 24949 8144 25001
rect 26803 24918 26861 24924
rect 26803 24884 26815 24918
rect 26849 24915 26861 24918
rect 26896 24915 26902 24927
rect 26849 24887 26902 24915
rect 26849 24884 26861 24887
rect 26803 24878 26861 24884
rect 26896 24875 26902 24887
rect 26954 24875 26960 24927
rect 31696 24875 31702 24927
rect 31754 24915 31760 24927
rect 33523 24918 33581 24924
rect 33523 24915 33535 24918
rect 31754 24887 33535 24915
rect 31754 24875 31760 24887
rect 33523 24884 33535 24887
rect 33569 24884 33581 24918
rect 33523 24878 33581 24884
rect 51184 24875 51190 24927
rect 51242 24915 51248 24927
rect 51283 24918 51341 24924
rect 51283 24915 51295 24918
rect 51242 24887 51295 24915
rect 51242 24875 51248 24887
rect 51283 24884 51295 24887
rect 51329 24884 51341 24918
rect 51283 24878 51341 24884
rect 8752 24767 8758 24779
rect 8640 24739 8758 24767
rect 8752 24727 8758 24739
rect 8810 24727 8816 24779
rect 1152 24668 58848 24690
rect 1152 24616 19654 24668
rect 19706 24616 19718 24668
rect 19770 24616 19782 24668
rect 19834 24616 19846 24668
rect 19898 24616 50374 24668
rect 50426 24616 50438 24668
rect 50490 24616 50502 24668
rect 50554 24616 50566 24668
rect 50618 24616 58848 24668
rect 1152 24594 58848 24616
rect 8080 24505 8086 24557
rect 8138 24545 8144 24557
rect 14128 24545 14134 24557
rect 8138 24517 14134 24545
rect 8138 24505 8144 24517
rect 14128 24505 14134 24517
rect 14186 24505 14192 24557
rect 35344 24175 35350 24187
rect 27346 24147 35350 24175
rect 10483 24104 10541 24110
rect 10483 24070 10495 24104
rect 10529 24101 10541 24104
rect 27346 24101 27374 24147
rect 35344 24135 35350 24147
rect 35402 24135 35408 24187
rect 10529 24073 27374 24101
rect 10529 24070 10541 24073
rect 10483 24064 10541 24070
rect 31984 24061 31990 24113
rect 32042 24101 32048 24113
rect 36595 24104 36653 24110
rect 36595 24101 36607 24104
rect 32042 24073 36607 24101
rect 32042 24061 32048 24073
rect 36595 24070 36607 24073
rect 36641 24070 36653 24104
rect 36595 24064 36653 24070
rect 41491 24104 41549 24110
rect 41491 24070 41503 24104
rect 41537 24101 41549 24104
rect 44752 24101 44758 24113
rect 41537 24073 44758 24101
rect 41537 24070 41549 24073
rect 41491 24064 41549 24070
rect 44752 24061 44758 24073
rect 44810 24061 44816 24113
rect 1152 24002 58848 24024
rect 1152 23950 4294 24002
rect 4346 23950 4358 24002
rect 4410 23950 4422 24002
rect 4474 23950 4486 24002
rect 4538 23950 35014 24002
rect 35066 23950 35078 24002
rect 35130 23950 35142 24002
rect 35194 23950 35206 24002
rect 35258 23950 58848 24002
rect 1152 23928 58848 23950
rect 8194 23851 8558 23879
rect 8194 23791 8222 23851
rect 8530 23805 8558 23851
rect 25456 23839 25462 23891
rect 25514 23879 25520 23891
rect 31984 23879 31990 23891
rect 25514 23851 31990 23879
rect 25514 23839 25520 23851
rect 31984 23839 31990 23851
rect 32042 23839 32048 23891
rect 15472 23805 15478 23817
rect 8530 23777 15478 23805
rect 15472 23765 15478 23777
rect 15530 23765 15536 23817
rect 19891 23660 19949 23666
rect 19891 23626 19903 23660
rect 19937 23657 19949 23660
rect 20179 23660 20237 23666
rect 20179 23657 20191 23660
rect 19937 23629 20191 23657
rect 19937 23626 19949 23629
rect 19891 23620 19949 23626
rect 20179 23626 20191 23629
rect 20225 23657 20237 23660
rect 34384 23657 34390 23669
rect 20225 23629 34390 23657
rect 20225 23626 20237 23629
rect 20179 23620 20237 23626
rect 34384 23617 34390 23629
rect 34442 23617 34448 23669
rect 29971 23586 30029 23592
rect 29971 23552 29983 23586
rect 30017 23583 30029 23586
rect 30067 23586 30125 23592
rect 30067 23583 30079 23586
rect 30017 23555 30079 23583
rect 30017 23552 30029 23555
rect 29971 23546 30029 23552
rect 30067 23552 30079 23555
rect 30113 23552 30125 23586
rect 30067 23546 30125 23552
rect 41779 23586 41837 23592
rect 41779 23552 41791 23586
rect 41825 23583 41837 23586
rect 41872 23583 41878 23595
rect 41825 23555 41878 23583
rect 41825 23552 41837 23555
rect 41779 23546 41837 23552
rect 41872 23543 41878 23555
rect 41930 23543 41936 23595
rect 44659 23586 44717 23592
rect 44659 23552 44671 23586
rect 44705 23552 44717 23586
rect 46960 23583 46966 23595
rect 46921 23555 46966 23583
rect 44659 23546 44717 23552
rect 8080 23509 8086 23521
rect 7968 23481 8086 23509
rect 8080 23469 8086 23481
rect 8138 23469 8144 23521
rect 13264 23509 13270 23521
rect 8242 23435 8270 23495
rect 8544 23481 13270 23509
rect 13264 23469 13270 23481
rect 13322 23469 13328 23521
rect 29392 23469 29398 23521
rect 29450 23509 29456 23521
rect 44674 23509 44702 23546
rect 46960 23543 46966 23555
rect 47018 23543 47024 23595
rect 29450 23481 44702 23509
rect 29450 23469 29456 23481
rect 8464 23435 8470 23447
rect 8242 23407 8470 23435
rect 8464 23395 8470 23407
rect 8522 23395 8528 23447
rect 30067 23438 30125 23444
rect 30067 23404 30079 23438
rect 30113 23435 30125 23438
rect 49744 23435 49750 23447
rect 30113 23407 49750 23435
rect 30113 23404 30125 23407
rect 30067 23398 30125 23404
rect 49744 23395 49750 23407
rect 49802 23395 49808 23447
rect 1152 23336 58848 23358
rect 1152 23284 19654 23336
rect 19706 23284 19718 23336
rect 19770 23284 19782 23336
rect 19834 23284 19846 23336
rect 19898 23284 50374 23336
rect 50426 23284 50438 23336
rect 50490 23284 50502 23336
rect 50554 23284 50566 23336
rect 50618 23284 58848 23336
rect 1152 23262 58848 23284
rect 8080 23173 8086 23225
rect 8138 23213 8144 23225
rect 13168 23213 13174 23225
rect 8138 23185 13174 23213
rect 8138 23173 8144 23185
rect 13168 23173 13174 23185
rect 13226 23173 13232 23225
rect 8464 23099 8470 23151
rect 8522 23139 8528 23151
rect 14032 23139 14038 23151
rect 8522 23111 14038 23139
rect 8522 23099 8528 23111
rect 14032 23099 14038 23111
rect 14090 23099 14096 23151
rect 10576 22877 10582 22929
rect 10634 22917 10640 22929
rect 55408 22917 55414 22929
rect 10634 22889 55414 22917
rect 10634 22877 10640 22889
rect 55408 22877 55414 22889
rect 55466 22877 55472 22929
rect 8080 22803 8086 22855
rect 8138 22843 8144 22855
rect 26608 22843 26614 22855
rect 8138 22815 26614 22843
rect 8138 22803 8144 22815
rect 26608 22803 26614 22815
rect 26666 22803 26672 22855
rect 46672 22843 46678 22855
rect 27346 22815 46678 22843
rect 10195 22772 10253 22778
rect 10195 22738 10207 22772
rect 10241 22769 10253 22772
rect 27346 22769 27374 22815
rect 46672 22803 46678 22815
rect 46730 22803 46736 22855
rect 37552 22769 37558 22781
rect 10241 22741 27374 22769
rect 37513 22741 37558 22769
rect 10241 22738 10253 22741
rect 10195 22732 10253 22738
rect 37552 22729 37558 22741
rect 37610 22729 37616 22781
rect 1152 22670 58848 22692
rect 1152 22618 4294 22670
rect 4346 22618 4358 22670
rect 4410 22618 4422 22670
rect 4474 22618 4486 22670
rect 4538 22618 35014 22670
rect 35066 22618 35078 22670
rect 35130 22618 35142 22670
rect 35194 22618 35206 22670
rect 35258 22618 58848 22670
rect 1152 22596 58848 22618
rect 8179 22550 8237 22556
rect 8179 22516 8191 22550
rect 8225 22547 8237 22550
rect 8225 22519 17294 22547
rect 8225 22516 8237 22519
rect 8179 22510 8237 22516
rect 8194 22459 8222 22510
rect 17266 22473 17294 22519
rect 25744 22507 25750 22559
rect 25802 22547 25808 22559
rect 37552 22547 37558 22559
rect 25802 22519 37558 22547
rect 25802 22507 25808 22519
rect 37552 22507 37558 22519
rect 37610 22507 37616 22559
rect 57616 22473 57622 22485
rect 17266 22445 57622 22473
rect 57616 22433 57622 22445
rect 57674 22433 57680 22485
rect 7968 22371 8126 22399
rect 8098 22337 8126 22371
rect 8080 22285 8086 22337
rect 8138 22285 8144 22337
rect 10576 22177 10582 22189
rect 8256 22149 10582 22177
rect 10576 22137 10582 22149
rect 10634 22137 10640 22189
rect 7603 22106 7661 22112
rect 7603 22072 7615 22106
rect 7649 22103 7661 22106
rect 8083 22106 8141 22112
rect 8083 22103 8095 22106
rect 7649 22075 8095 22103
rect 7649 22072 7661 22075
rect 7603 22066 7661 22072
rect 8083 22072 8095 22075
rect 8129 22072 8141 22106
rect 8083 22066 8141 22072
rect 1152 22004 58848 22026
rect 1152 21952 19654 22004
rect 19706 21952 19718 22004
rect 19770 21952 19782 22004
rect 19834 21952 19846 22004
rect 19898 21952 50374 22004
rect 50426 21952 50438 22004
rect 50490 21952 50502 22004
rect 50554 21952 50566 22004
rect 50618 21952 58848 22004
rect 1152 21930 58848 21952
rect 7987 21662 8045 21668
rect 7987 21628 7999 21662
rect 8033 21659 8045 21662
rect 8275 21662 8333 21668
rect 8275 21659 8287 21662
rect 8033 21631 8287 21659
rect 8033 21628 8045 21631
rect 7987 21622 8045 21628
rect 8275 21628 8287 21631
rect 8321 21659 8333 21662
rect 43888 21659 43894 21671
rect 8321 21631 43894 21659
rect 8321 21628 8333 21631
rect 8275 21622 8333 21628
rect 43888 21619 43894 21631
rect 43946 21619 43952 21671
rect 8080 21545 8086 21597
rect 8138 21585 8144 21597
rect 48688 21585 48694 21597
rect 8138 21557 48694 21585
rect 8138 21545 8144 21557
rect 48688 21545 48694 21557
rect 48746 21545 48752 21597
rect 52816 21511 52822 21523
rect 17266 21483 52822 21511
rect 8560 21397 8566 21449
rect 8618 21437 8624 21449
rect 17266 21437 17294 21483
rect 52816 21471 52822 21483
rect 52874 21471 52880 21523
rect 8618 21409 17294 21437
rect 32851 21440 32909 21446
rect 8618 21397 8624 21409
rect 32851 21406 32863 21440
rect 32897 21437 32909 21440
rect 33040 21437 33046 21449
rect 32897 21409 33046 21437
rect 32897 21406 32909 21409
rect 32851 21400 32909 21406
rect 33040 21397 33046 21409
rect 33098 21397 33104 21449
rect 1152 21338 58848 21360
rect 1152 21286 4294 21338
rect 4346 21286 4358 21338
rect 4410 21286 4422 21338
rect 4474 21286 4486 21338
rect 4538 21286 35014 21338
rect 35066 21286 35078 21338
rect 35130 21286 35142 21338
rect 35194 21286 35206 21338
rect 35258 21286 58848 21338
rect 1152 21264 58848 21286
rect 8080 20899 8086 20951
rect 8138 20919 8144 20951
rect 50800 20919 50806 20931
rect 8138 20899 8256 20919
rect 8098 20891 8256 20899
rect 17266 20891 50806 20919
rect 17266 20845 17294 20891
rect 50800 20879 50806 20891
rect 50858 20879 50864 20931
rect 7600 20771 7606 20783
rect 7561 20743 7606 20771
rect 7600 20731 7606 20743
rect 7658 20731 7664 20783
rect 8194 20771 8222 20831
rect 9120 20817 17294 20845
rect 8560 20771 8566 20783
rect 8194 20743 8566 20771
rect 8560 20731 8566 20743
rect 8618 20731 8624 20783
rect 8752 20731 8758 20783
rect 8810 20731 8816 20783
rect 9328 20731 9334 20783
rect 9386 20771 9392 20783
rect 55504 20771 55510 20783
rect 9386 20743 55510 20771
rect 9386 20731 9392 20743
rect 55504 20731 55510 20743
rect 55562 20731 55568 20783
rect 1152 20672 58848 20694
rect 1152 20620 19654 20672
rect 19706 20620 19718 20672
rect 19770 20620 19782 20672
rect 19834 20620 19846 20672
rect 19898 20620 50374 20672
rect 50426 20620 50438 20672
rect 50490 20620 50502 20672
rect 50554 20620 50566 20672
rect 50618 20620 58848 20672
rect 1152 20598 58848 20620
rect 7600 20509 7606 20561
rect 7658 20549 7664 20561
rect 8752 20549 8758 20561
rect 7658 20521 8758 20549
rect 7658 20509 7664 20521
rect 8752 20509 8758 20521
rect 8810 20549 8816 20561
rect 9328 20549 9334 20561
rect 8810 20521 9334 20549
rect 8810 20509 8816 20521
rect 9328 20509 9334 20521
rect 9386 20509 9392 20561
rect 24019 20182 24077 20188
rect 24019 20148 24031 20182
rect 24065 20179 24077 20182
rect 24307 20182 24365 20188
rect 24307 20179 24319 20182
rect 24065 20151 24319 20179
rect 24065 20148 24077 20151
rect 24019 20142 24077 20148
rect 24307 20148 24319 20151
rect 24353 20179 24365 20182
rect 44176 20179 44182 20191
rect 24353 20151 44182 20179
rect 24353 20148 24365 20151
rect 24307 20142 24365 20148
rect 44176 20139 44182 20151
rect 44234 20139 44240 20191
rect 7600 20065 7606 20117
rect 7658 20105 7664 20117
rect 8752 20105 8758 20117
rect 7658 20077 8758 20105
rect 7658 20065 7664 20077
rect 8752 20065 8758 20077
rect 8810 20065 8816 20117
rect 16147 20108 16205 20114
rect 16147 20074 16159 20108
rect 16193 20105 16205 20108
rect 16720 20105 16726 20117
rect 16193 20077 16726 20105
rect 16193 20074 16205 20077
rect 16147 20068 16205 20074
rect 16720 20065 16726 20077
rect 16778 20065 16784 20117
rect 27571 20108 27629 20114
rect 27571 20074 27583 20108
rect 27617 20105 27629 20108
rect 32560 20105 32566 20117
rect 27617 20077 32566 20105
rect 27617 20074 27629 20077
rect 27571 20068 27629 20074
rect 32560 20065 32566 20077
rect 32618 20065 32624 20117
rect 1152 20006 58848 20028
rect 1152 19954 4294 20006
rect 4346 19954 4358 20006
rect 4410 19954 4422 20006
rect 4474 19954 4486 20006
rect 4538 19954 35014 20006
rect 35066 19954 35078 20006
rect 35130 19954 35142 20006
rect 35194 19954 35206 20006
rect 35258 19954 58848 20006
rect 1152 19932 58848 19954
rect 7600 19883 7606 19895
rect 7561 19855 7606 19883
rect 7600 19843 7606 19855
rect 7658 19843 7664 19895
rect 8752 19843 8758 19895
rect 8810 19883 8816 19895
rect 48784 19883 48790 19895
rect 8810 19855 48790 19883
rect 8810 19843 8816 19855
rect 48784 19843 48790 19855
rect 48842 19843 48848 19895
rect 8770 19795 8798 19843
rect 16720 19769 16726 19821
rect 16778 19809 16784 19821
rect 40336 19809 40342 19821
rect 16778 19781 40342 19809
rect 16778 19769 16784 19781
rect 40336 19769 40342 19781
rect 40394 19769 40400 19821
rect 6835 19590 6893 19596
rect 6835 19556 6847 19590
rect 6881 19587 6893 19590
rect 7120 19587 7126 19599
rect 6881 19559 7126 19587
rect 6881 19556 6893 19559
rect 6835 19550 6893 19556
rect 7120 19547 7126 19559
rect 7178 19547 7184 19599
rect 34768 19587 34774 19599
rect 34729 19559 34774 19587
rect 34768 19547 34774 19559
rect 34826 19547 34832 19599
rect 8272 19473 8278 19525
rect 8330 19473 8336 19525
rect 9040 19473 9046 19525
rect 9098 19513 9104 19525
rect 46096 19513 46102 19525
rect 9098 19485 46102 19513
rect 9098 19473 9104 19485
rect 46096 19473 46102 19485
rect 46154 19473 46160 19525
rect 1152 19340 58848 19362
rect 1152 19288 19654 19340
rect 19706 19288 19718 19340
rect 19770 19288 19782 19340
rect 19834 19288 19846 19340
rect 19898 19288 50374 19340
rect 50426 19288 50438 19340
rect 50490 19288 50502 19340
rect 50554 19288 50566 19340
rect 50618 19288 58848 19340
rect 1152 19266 58848 19288
rect 7120 19177 7126 19229
rect 7178 19217 7184 19229
rect 49840 19217 49846 19229
rect 7178 19189 49846 19217
rect 7178 19177 7184 19189
rect 49840 19177 49846 19189
rect 49898 19177 49904 19229
rect 2512 19103 2518 19155
rect 2570 19143 2576 19155
rect 34768 19143 34774 19155
rect 2570 19115 34774 19143
rect 2570 19103 2576 19115
rect 34768 19103 34774 19115
rect 34826 19103 34832 19155
rect 39856 18881 39862 18933
rect 39914 18921 39920 18933
rect 48691 18924 48749 18930
rect 48691 18921 48703 18924
rect 39914 18893 48703 18921
rect 39914 18881 39920 18893
rect 48691 18890 48703 18893
rect 48737 18921 48749 18924
rect 48883 18924 48941 18930
rect 48883 18921 48895 18924
rect 48737 18893 48895 18921
rect 48737 18890 48749 18893
rect 48691 18884 48749 18890
rect 48883 18890 48895 18893
rect 48929 18890 48941 18924
rect 48883 18884 48941 18890
rect 21232 18773 21238 18785
rect 21193 18745 21238 18773
rect 21232 18733 21238 18745
rect 21290 18733 21296 18785
rect 47632 18733 47638 18785
rect 47690 18773 47696 18785
rect 52051 18776 52109 18782
rect 52051 18773 52063 18776
rect 47690 18745 52063 18773
rect 47690 18733 47696 18745
rect 52051 18742 52063 18745
rect 52097 18742 52109 18776
rect 52051 18736 52109 18742
rect 1152 18674 58848 18696
rect 1152 18622 4294 18674
rect 4346 18622 4358 18674
rect 4410 18622 4422 18674
rect 4474 18622 4486 18674
rect 4538 18622 35014 18674
rect 35066 18622 35078 18674
rect 35130 18622 35142 18674
rect 35194 18622 35206 18674
rect 35258 18622 58848 18674
rect 1152 18600 58848 18622
rect 7603 18554 7661 18560
rect 7603 18520 7615 18554
rect 7649 18551 7661 18554
rect 7891 18554 7949 18560
rect 7891 18551 7903 18554
rect 7649 18523 7903 18551
rect 7649 18520 7661 18523
rect 7603 18514 7661 18520
rect 7891 18520 7903 18523
rect 7937 18520 7949 18554
rect 7891 18514 7949 18520
rect 8179 18554 8237 18560
rect 8179 18520 8191 18554
rect 8225 18551 8237 18554
rect 8225 18523 17294 18551
rect 8225 18520 8237 18523
rect 8179 18514 8237 18520
rect 8194 18463 8222 18514
rect 17266 18477 17294 18523
rect 45232 18477 45238 18489
rect 17266 18449 45238 18477
rect 45232 18437 45238 18449
rect 45290 18437 45296 18489
rect 8098 18267 8126 18368
rect 47152 18329 47158 18341
rect 27346 18301 47158 18329
rect 1747 18258 1805 18264
rect 1747 18224 1759 18258
rect 1793 18255 1805 18258
rect 7408 18255 7414 18267
rect 1793 18227 7414 18255
rect 1793 18224 1805 18227
rect 1747 18218 1805 18224
rect 7408 18215 7414 18227
rect 7466 18215 7472 18267
rect 8080 18215 8086 18267
rect 8138 18215 8144 18267
rect 24499 18258 24557 18264
rect 24499 18224 24511 18258
rect 24545 18255 24557 18258
rect 27346 18255 27374 18301
rect 47152 18289 47158 18301
rect 47210 18289 47216 18341
rect 51664 18329 51670 18341
rect 47506 18301 51670 18329
rect 40720 18255 40726 18267
rect 24545 18227 27374 18255
rect 40681 18227 40726 18255
rect 24545 18224 24557 18227
rect 24499 18218 24557 18224
rect 40720 18215 40726 18227
rect 40778 18215 40784 18267
rect 47506 18181 47534 18301
rect 51664 18289 51670 18301
rect 51722 18289 51728 18341
rect 51187 18258 51245 18264
rect 51187 18224 51199 18258
rect 51233 18224 51245 18258
rect 51187 18218 51245 18224
rect 27346 18153 47534 18181
rect 26131 18110 26189 18116
rect 26131 18076 26143 18110
rect 26177 18107 26189 18110
rect 26419 18110 26477 18116
rect 26419 18107 26431 18110
rect 26177 18079 26431 18107
rect 26177 18076 26189 18079
rect 26131 18070 26189 18076
rect 26419 18076 26431 18079
rect 26465 18107 26477 18110
rect 27346 18107 27374 18153
rect 50992 18107 50998 18119
rect 26465 18079 27374 18107
rect 50953 18079 50998 18107
rect 26465 18076 26477 18079
rect 26419 18070 26477 18076
rect 50992 18067 50998 18079
rect 51050 18107 51056 18119
rect 51202 18107 51230 18218
rect 51050 18079 51230 18107
rect 51050 18067 51056 18079
rect 1152 18008 58848 18030
rect 1152 17956 19654 18008
rect 19706 17956 19718 18008
rect 19770 17956 19782 18008
rect 19834 17956 19846 18008
rect 19898 17956 50374 18008
rect 50426 17956 50438 18008
rect 50490 17956 50502 18008
rect 50554 17956 50566 18008
rect 50618 17956 58848 18008
rect 1152 17934 58848 17956
rect 7792 17845 7798 17897
rect 7850 17885 7856 17897
rect 7850 17857 17294 17885
rect 7850 17845 7856 17857
rect 17266 17811 17294 17857
rect 50992 17811 50998 17823
rect 17266 17783 50998 17811
rect 50992 17771 50998 17783
rect 51050 17771 51056 17823
rect 8080 17697 8086 17749
rect 8138 17737 8144 17749
rect 42928 17737 42934 17749
rect 8138 17709 42934 17737
rect 8138 17697 8144 17709
rect 42928 17697 42934 17709
rect 42986 17697 42992 17749
rect 30643 17666 30701 17672
rect 30643 17632 30655 17666
rect 30689 17663 30701 17666
rect 30931 17666 30989 17672
rect 30931 17663 30943 17666
rect 30689 17635 30943 17663
rect 30689 17632 30701 17635
rect 30643 17626 30701 17632
rect 30931 17632 30943 17635
rect 30977 17663 30989 17666
rect 35824 17663 35830 17675
rect 30977 17635 35830 17663
rect 30977 17632 30989 17635
rect 30931 17626 30989 17632
rect 35824 17623 35830 17635
rect 35882 17623 35888 17675
rect 7408 17475 7414 17527
rect 7466 17515 7472 17527
rect 8560 17515 8566 17527
rect 7466 17487 8566 17515
rect 7466 17475 7472 17487
rect 8560 17475 8566 17487
rect 8618 17475 8624 17527
rect 1939 17444 1997 17450
rect 1939 17410 1951 17444
rect 1985 17441 1997 17444
rect 23728 17441 23734 17453
rect 1985 17413 23734 17441
rect 1985 17410 1997 17413
rect 1939 17404 1997 17410
rect 23728 17401 23734 17413
rect 23786 17401 23792 17453
rect 1152 17342 58848 17364
rect 1152 17290 4294 17342
rect 4346 17290 4358 17342
rect 4410 17290 4422 17342
rect 4474 17290 4486 17342
rect 4538 17290 35014 17342
rect 35066 17290 35078 17342
rect 35130 17290 35142 17342
rect 35194 17290 35206 17342
rect 35258 17290 58848 17342
rect 1152 17268 58848 17290
rect 15088 16957 15094 17009
rect 15146 16997 15152 17009
rect 56755 17000 56813 17006
rect 56755 16997 56767 17000
rect 15146 16969 56767 16997
rect 15146 16957 15152 16969
rect 56755 16966 56767 16969
rect 56801 16966 56813 17000
rect 56755 16960 56813 16966
rect 5968 16923 5974 16935
rect 5929 16895 5974 16923
rect 5968 16883 5974 16895
rect 6026 16883 6032 16935
rect 7120 16923 7126 16935
rect 7081 16895 7126 16923
rect 7120 16883 7126 16895
rect 7178 16883 7184 16935
rect 46864 16923 46870 16935
rect 46825 16895 46870 16923
rect 46864 16883 46870 16895
rect 46922 16883 46928 16935
rect 55984 16923 55990 16935
rect 55945 16895 55990 16923
rect 55984 16883 55990 16895
rect 56042 16883 56048 16935
rect 39760 16849 39766 16861
rect 7968 16821 39766 16849
rect 39760 16809 39766 16821
rect 39818 16809 39824 16861
rect 7603 16778 7661 16784
rect 7603 16744 7615 16778
rect 7649 16775 7661 16778
rect 42640 16775 42646 16787
rect 7649 16747 42646 16775
rect 7649 16744 7661 16747
rect 7603 16738 7661 16744
rect 42640 16735 42646 16747
rect 42698 16735 42704 16787
rect 1152 16676 58848 16698
rect 1152 16624 19654 16676
rect 19706 16624 19718 16676
rect 19770 16624 19782 16676
rect 19834 16624 19846 16676
rect 19898 16624 50374 16676
rect 50426 16624 50438 16676
rect 50490 16624 50502 16676
rect 50554 16624 50566 16676
rect 50618 16624 58848 16676
rect 1152 16602 58848 16624
rect 5968 16513 5974 16565
rect 6026 16553 6032 16565
rect 13552 16553 13558 16565
rect 6026 16525 13558 16553
rect 6026 16513 6032 16525
rect 13552 16513 13558 16525
rect 13610 16513 13616 16565
rect 30160 16513 30166 16565
rect 30218 16553 30224 16565
rect 46864 16553 46870 16565
rect 30218 16525 46870 16553
rect 30218 16513 30224 16525
rect 46864 16513 46870 16525
rect 46922 16513 46928 16565
rect 7120 16439 7126 16491
rect 7178 16479 7184 16491
rect 54064 16479 54070 16491
rect 7178 16451 54070 16479
rect 7178 16439 7184 16451
rect 54064 16439 54070 16451
rect 54122 16439 54128 16491
rect 27091 16112 27149 16118
rect 27091 16078 27103 16112
rect 27137 16109 27149 16112
rect 52432 16109 52438 16121
rect 27137 16081 52438 16109
rect 27137 16078 27149 16081
rect 27091 16072 27149 16078
rect 52432 16069 52438 16081
rect 52490 16069 52496 16121
rect 1152 16010 58848 16032
rect 1152 15958 4294 16010
rect 4346 15958 4358 16010
rect 4410 15958 4422 16010
rect 4474 15958 4486 16010
rect 4538 15958 35014 16010
rect 35066 15958 35078 16010
rect 35130 15958 35142 16010
rect 35194 15958 35206 16010
rect 35258 15958 58848 16010
rect 1152 15936 58848 15958
rect 21424 15551 21430 15603
rect 21482 15591 21488 15603
rect 46867 15594 46925 15600
rect 46867 15591 46879 15594
rect 21482 15563 46879 15591
rect 21482 15551 21488 15563
rect 46867 15560 46879 15563
rect 46913 15591 46925 15594
rect 47059 15594 47117 15600
rect 47059 15591 47071 15594
rect 46913 15563 47071 15591
rect 46913 15560 46925 15563
rect 46867 15554 46925 15560
rect 47059 15560 47071 15563
rect 47105 15560 47117 15594
rect 47059 15554 47117 15560
rect 36688 15517 36694 15529
rect 7968 15489 36694 15517
rect 36688 15477 36694 15489
rect 36746 15477 36752 15529
rect 7603 15446 7661 15452
rect 7603 15412 7615 15446
rect 7649 15443 7661 15446
rect 38896 15443 38902 15455
rect 7649 15415 38902 15443
rect 7649 15412 7661 15415
rect 7603 15406 7661 15412
rect 38896 15403 38902 15415
rect 38954 15403 38960 15455
rect 1152 15344 58848 15366
rect 1152 15292 19654 15344
rect 19706 15292 19718 15344
rect 19770 15292 19782 15344
rect 19834 15292 19846 15344
rect 19898 15292 50374 15344
rect 50426 15292 50438 15344
rect 50490 15292 50502 15344
rect 50554 15292 50566 15344
rect 50618 15292 58848 15344
rect 1152 15270 58848 15292
rect 12307 15224 12365 15230
rect 12307 15190 12319 15224
rect 12353 15221 12365 15224
rect 12595 15224 12653 15230
rect 12595 15221 12607 15224
rect 12353 15193 12607 15221
rect 12353 15190 12365 15193
rect 12307 15184 12365 15190
rect 12595 15190 12607 15193
rect 12641 15221 12653 15224
rect 13648 15221 13654 15233
rect 12641 15193 13654 15221
rect 12641 15190 12653 15193
rect 12595 15184 12653 15190
rect 13648 15181 13654 15193
rect 13706 15181 13712 15233
rect 22192 15181 22198 15233
rect 22250 15221 22256 15233
rect 24019 15224 24077 15230
rect 24019 15221 24031 15224
rect 22250 15193 24031 15221
rect 22250 15181 22256 15193
rect 24019 15190 24031 15193
rect 24065 15190 24077 15224
rect 24019 15184 24077 15190
rect 24034 15073 24062 15184
rect 24211 15076 24269 15082
rect 24211 15073 24223 15076
rect 24034 15045 24223 15073
rect 24211 15042 24223 15045
rect 24257 15042 24269 15076
rect 24211 15036 24269 15042
rect 57715 15076 57773 15082
rect 57715 15042 57727 15076
rect 57761 15073 57773 15076
rect 58000 15073 58006 15085
rect 57761 15045 58006 15073
rect 57761 15042 57773 15045
rect 57715 15036 57773 15042
rect 58000 15033 58006 15045
rect 58058 15033 58064 15085
rect 17776 14885 17782 14937
rect 17834 14925 17840 14937
rect 46576 14925 46582 14937
rect 17834 14897 46582 14925
rect 17834 14885 17840 14897
rect 46576 14885 46582 14897
rect 46634 14885 46640 14937
rect 7696 14811 7702 14863
rect 7754 14851 7760 14863
rect 23731 14854 23789 14860
rect 23731 14851 23743 14854
rect 7754 14823 23743 14851
rect 7754 14811 7760 14823
rect 23731 14820 23743 14823
rect 23777 14820 23789 14854
rect 23731 14814 23789 14820
rect 1152 14678 58848 14700
rect 1152 14626 4294 14678
rect 4346 14626 4358 14678
rect 4410 14626 4422 14678
rect 4474 14626 4486 14678
rect 4538 14626 35014 14678
rect 35066 14626 35078 14678
rect 35130 14626 35142 14678
rect 35194 14626 35206 14678
rect 35258 14626 58848 14678
rect 1152 14604 58848 14626
rect 3571 14558 3629 14564
rect 3571 14524 3583 14558
rect 3617 14555 3629 14558
rect 3859 14558 3917 14564
rect 3859 14555 3871 14558
rect 3617 14527 3871 14555
rect 3617 14524 3629 14527
rect 3571 14518 3629 14524
rect 3859 14524 3871 14527
rect 3905 14555 3917 14558
rect 45040 14555 45046 14567
rect 3905 14527 45046 14555
rect 3905 14524 3917 14527
rect 3859 14518 3917 14524
rect 45040 14515 45046 14527
rect 45098 14515 45104 14567
rect 12691 14484 12749 14490
rect 12691 14450 12703 14484
rect 12737 14481 12749 14484
rect 45232 14481 45238 14493
rect 12737 14453 45238 14481
rect 12737 14450 12749 14453
rect 12691 14444 12749 14450
rect 45232 14441 45238 14453
rect 45290 14441 45296 14493
rect 17491 14410 17549 14416
rect 17491 14376 17503 14410
rect 17537 14407 17549 14410
rect 17776 14407 17782 14419
rect 17537 14379 17782 14407
rect 17537 14376 17549 14379
rect 17491 14370 17549 14376
rect 17776 14367 17782 14379
rect 17834 14367 17840 14419
rect 34096 14185 34102 14197
rect 7968 14157 34102 14185
rect 34096 14145 34102 14157
rect 34154 14145 34160 14197
rect 4435 14114 4493 14120
rect 4435 14080 4447 14114
rect 4481 14111 4493 14114
rect 4720 14111 4726 14123
rect 4481 14083 4726 14111
rect 4481 14080 4493 14083
rect 4435 14074 4493 14080
rect 4720 14071 4726 14083
rect 4778 14071 4784 14123
rect 7603 14114 7661 14120
rect 7603 14080 7615 14114
rect 7649 14111 7661 14114
rect 36784 14111 36790 14123
rect 7649 14083 36790 14111
rect 7649 14080 7661 14083
rect 7603 14074 7661 14080
rect 36784 14071 36790 14083
rect 36842 14071 36848 14123
rect 1152 14012 58848 14034
rect 1152 13960 19654 14012
rect 19706 13960 19718 14012
rect 19770 13960 19782 14012
rect 19834 13960 19846 14012
rect 19898 13960 50374 14012
rect 50426 13960 50438 14012
rect 50490 13960 50502 14012
rect 50554 13960 50566 14012
rect 50618 13960 58848 14012
rect 1152 13938 58848 13960
rect 4720 13849 4726 13901
rect 4778 13889 4784 13901
rect 27472 13889 27478 13901
rect 4778 13861 27478 13889
rect 4778 13849 4784 13861
rect 27472 13849 27478 13861
rect 27530 13849 27536 13901
rect 9232 13701 9238 13753
rect 9290 13741 9296 13753
rect 25648 13741 25654 13753
rect 9290 13713 25654 13741
rect 9290 13701 9296 13713
rect 25648 13701 25654 13713
rect 25706 13701 25712 13753
rect 47635 13744 47693 13750
rect 47635 13741 47647 13744
rect 47506 13713 47647 13741
rect 7600 13627 7606 13679
rect 7658 13667 7664 13679
rect 9904 13667 9910 13679
rect 7658 13639 9910 13667
rect 7658 13627 7664 13639
rect 9904 13627 9910 13639
rect 9962 13667 9968 13679
rect 32848 13667 32854 13679
rect 9962 13639 32854 13667
rect 9962 13627 9968 13639
rect 32848 13627 32854 13639
rect 32906 13627 32912 13679
rect 8368 13479 8374 13531
rect 8426 13519 8432 13531
rect 29968 13519 29974 13531
rect 8426 13491 29974 13519
rect 8426 13479 8432 13491
rect 29968 13479 29974 13491
rect 30026 13479 30032 13531
rect 8560 13405 8566 13457
rect 8618 13445 8624 13457
rect 9808 13445 9814 13457
rect 8618 13417 9814 13445
rect 8618 13405 8624 13417
rect 9808 13405 9814 13417
rect 9866 13405 9872 13457
rect 15088 13445 15094 13457
rect 15049 13417 15094 13445
rect 15088 13405 15094 13417
rect 15146 13405 15152 13457
rect 47347 13448 47405 13454
rect 47347 13414 47359 13448
rect 47393 13445 47405 13448
rect 47506 13445 47534 13713
rect 47635 13710 47647 13713
rect 47681 13741 47693 13744
rect 51568 13741 51574 13753
rect 47681 13713 51574 13741
rect 47681 13710 47693 13713
rect 47635 13704 47693 13710
rect 51568 13701 51574 13713
rect 51626 13701 51632 13753
rect 47393 13417 47534 13445
rect 47393 13414 47405 13417
rect 47347 13408 47405 13414
rect 1152 13346 58848 13368
rect 1152 13294 4294 13346
rect 4346 13294 4358 13346
rect 4410 13294 4422 13346
rect 4474 13294 4486 13346
rect 4538 13294 35014 13346
rect 35066 13294 35078 13346
rect 35130 13294 35142 13346
rect 35194 13294 35206 13346
rect 35258 13294 58848 13346
rect 1152 13272 58848 13294
rect 7600 13223 7606 13235
rect 7561 13195 7606 13223
rect 7600 13183 7606 13195
rect 7658 13183 7664 13235
rect 15088 13183 15094 13235
rect 15146 13223 15152 13235
rect 48304 13223 48310 13235
rect 15146 13195 48310 13223
rect 15146 13183 15152 13195
rect 48304 13183 48310 13195
rect 48362 13183 48368 13235
rect 8368 13149 8374 13161
rect 8256 13121 8374 13149
rect 8368 13109 8374 13121
rect 8426 13109 8432 13161
rect 26707 13152 26765 13158
rect 26707 13118 26719 13152
rect 26753 13149 26765 13152
rect 36208 13149 36214 13161
rect 26753 13121 36214 13149
rect 26753 13118 26765 13121
rect 26707 13112 26765 13118
rect 36208 13109 36214 13121
rect 36266 13109 36272 13161
rect 34000 13035 34006 13087
rect 34058 13075 34064 13087
rect 48979 13078 49037 13084
rect 48979 13075 48991 13078
rect 34058 13047 48991 13075
rect 34058 13035 34064 13047
rect 48979 13044 48991 13047
rect 49025 13075 49037 13078
rect 49171 13078 49229 13084
rect 49171 13075 49183 13078
rect 49025 13047 49183 13075
rect 49025 13044 49037 13047
rect 48979 13038 49037 13044
rect 49171 13044 49183 13047
rect 49217 13044 49229 13078
rect 49171 13038 49229 13044
rect 28144 12961 28150 13013
rect 28202 13001 28208 13013
rect 58003 13004 58061 13010
rect 58003 13001 58015 13004
rect 28202 12973 58015 13001
rect 28202 12961 28208 12973
rect 58003 12970 58015 12973
rect 58049 12970 58061 13004
rect 58003 12964 58061 12970
rect 9904 12779 9910 12791
rect 9793 12751 9910 12779
rect 9904 12739 9910 12751
rect 9962 12739 9968 12791
rect 1152 12680 58848 12702
rect 1152 12628 19654 12680
rect 19706 12628 19718 12680
rect 19770 12628 19782 12680
rect 19834 12628 19846 12680
rect 19898 12628 50374 12680
rect 50426 12628 50438 12680
rect 50490 12628 50502 12680
rect 50554 12628 50566 12680
rect 50618 12628 58848 12680
rect 1152 12606 58848 12628
rect 8560 12517 8566 12569
rect 8618 12557 8624 12569
rect 29296 12557 29302 12569
rect 8618 12529 29302 12557
rect 8618 12517 8624 12529
rect 29296 12517 29302 12529
rect 29354 12517 29360 12569
rect 6832 12369 6838 12421
rect 6890 12409 6896 12421
rect 13072 12409 13078 12421
rect 6890 12381 13078 12409
rect 6890 12369 6896 12381
rect 13072 12369 13078 12381
rect 13130 12369 13136 12421
rect 56944 12369 56950 12421
rect 57002 12409 57008 12421
rect 57715 12412 57773 12418
rect 57715 12409 57727 12412
rect 57002 12381 57727 12409
rect 57002 12369 57008 12381
rect 57715 12378 57727 12381
rect 57761 12378 57773 12412
rect 57715 12372 57773 12378
rect 8080 12295 8086 12347
rect 8138 12335 8144 12347
rect 27184 12335 27190 12347
rect 8138 12307 27190 12335
rect 8138 12295 8144 12307
rect 27184 12295 27190 12307
rect 27242 12295 27248 12347
rect 27346 12307 37454 12335
rect 12496 12261 12502 12273
rect 5746 12233 12502 12261
rect 5200 12147 5206 12199
rect 5258 12187 5264 12199
rect 5746 12187 5774 12233
rect 12496 12221 12502 12233
rect 12554 12221 12560 12273
rect 12784 12221 12790 12273
rect 12842 12261 12848 12273
rect 27346 12261 27374 12307
rect 12842 12233 27374 12261
rect 31315 12264 31373 12270
rect 12842 12221 12848 12233
rect 31315 12230 31327 12264
rect 31361 12230 31373 12264
rect 37426 12261 37454 12307
rect 47536 12261 47542 12273
rect 37426 12233 47542 12261
rect 31315 12224 31373 12230
rect 15856 12187 15862 12199
rect 5258 12159 5774 12187
rect 10786 12159 15862 12187
rect 5258 12147 5264 12159
rect 5011 12116 5069 12122
rect 5011 12082 5023 12116
rect 5057 12113 5069 12116
rect 10786 12113 10814 12159
rect 15856 12147 15862 12159
rect 15914 12147 15920 12199
rect 31027 12190 31085 12196
rect 31027 12156 31039 12190
rect 31073 12187 31085 12190
rect 31330 12187 31358 12224
rect 47536 12221 47542 12233
rect 47594 12221 47600 12273
rect 57520 12221 57526 12273
rect 57578 12261 57584 12273
rect 57619 12264 57677 12270
rect 57619 12261 57631 12264
rect 57578 12233 57631 12261
rect 57578 12221 57584 12233
rect 57619 12230 57631 12233
rect 57665 12230 57677 12264
rect 57619 12224 57677 12230
rect 42448 12187 42454 12199
rect 31073 12159 42454 12187
rect 31073 12156 31085 12159
rect 31027 12150 31085 12156
rect 42448 12147 42454 12159
rect 42506 12147 42512 12199
rect 15184 12113 15190 12125
rect 5057 12085 10814 12113
rect 15145 12085 15190 12113
rect 5057 12082 5069 12085
rect 5011 12076 5069 12082
rect 15184 12073 15190 12085
rect 15242 12073 15248 12125
rect 18736 12113 18742 12125
rect 18697 12085 18742 12113
rect 18736 12073 18742 12085
rect 18794 12073 18800 12125
rect 29587 12116 29645 12122
rect 29587 12082 29599 12116
rect 29633 12113 29645 12116
rect 33520 12113 33526 12125
rect 29633 12085 33526 12113
rect 29633 12082 29645 12085
rect 29587 12076 29645 12082
rect 33520 12073 33526 12085
rect 33578 12073 33584 12125
rect 1152 12014 58848 12036
rect 1152 11962 4294 12014
rect 4346 11962 4358 12014
rect 4410 11962 4422 12014
rect 4474 11962 4486 12014
rect 4538 11962 35014 12014
rect 35066 11962 35078 12014
rect 35130 11962 35142 12014
rect 35194 11962 35206 12014
rect 35258 11962 58848 12014
rect 1152 11940 58848 11962
rect 1744 11891 1750 11903
rect 1705 11863 1750 11891
rect 1744 11851 1750 11863
rect 1802 11891 1808 11903
rect 1843 11894 1901 11900
rect 1843 11891 1855 11894
rect 1802 11863 1855 11891
rect 1802 11851 1808 11863
rect 1843 11860 1855 11863
rect 1889 11860 1901 11894
rect 5200 11891 5206 11903
rect 5161 11863 5206 11891
rect 1843 11854 1901 11860
rect 5200 11851 5206 11863
rect 5258 11851 5264 11903
rect 7603 11894 7661 11900
rect 7603 11860 7615 11894
rect 7649 11891 7661 11894
rect 8368 11891 8374 11903
rect 7649 11863 7934 11891
rect 7649 11860 7661 11863
rect 7603 11854 7661 11860
rect 7906 11817 7934 11863
rect 8290 11863 8374 11891
rect 8290 11817 8318 11863
rect 8368 11851 8374 11863
rect 8426 11851 8432 11903
rect 15184 11851 15190 11903
rect 15242 11891 15248 11903
rect 42928 11891 42934 11903
rect 15242 11863 42934 11891
rect 15242 11851 15248 11863
rect 42928 11851 42934 11863
rect 42986 11851 42992 11903
rect 7906 11789 8318 11817
rect 8560 11777 8566 11829
rect 8618 11777 8624 11829
rect 8080 11743 8086 11755
rect 7968 11715 8086 11743
rect 8080 11703 8086 11715
rect 8138 11703 8144 11755
rect 24304 11703 24310 11755
rect 24362 11743 24368 11755
rect 56467 11746 56525 11752
rect 24362 11715 47534 11743
rect 24362 11703 24368 11715
rect 9235 11672 9293 11678
rect 9235 11638 9247 11672
rect 9281 11669 9293 11672
rect 9523 11672 9581 11678
rect 9523 11669 9535 11672
rect 9281 11641 9535 11669
rect 9281 11638 9293 11641
rect 9235 11632 9293 11638
rect 9523 11638 9535 11641
rect 9569 11669 9581 11672
rect 40432 11669 40438 11681
rect 9569 11641 40438 11669
rect 9569 11638 9581 11641
rect 9523 11632 9581 11638
rect 40432 11629 40438 11641
rect 40490 11629 40496 11681
rect 47506 11669 47534 11715
rect 56467 11712 56479 11746
rect 56513 11743 56525 11746
rect 56513 11715 57614 11743
rect 56513 11712 56525 11715
rect 56467 11706 56525 11712
rect 56947 11672 57005 11678
rect 56947 11669 56959 11672
rect 47506 11641 56959 11669
rect 56947 11638 56959 11641
rect 56993 11669 57005 11672
rect 57235 11672 57293 11678
rect 57235 11669 57247 11672
rect 56993 11641 57247 11669
rect 56993 11638 57005 11641
rect 56947 11632 57005 11638
rect 57235 11638 57247 11641
rect 57281 11638 57293 11672
rect 57235 11632 57293 11638
rect 37651 11598 37709 11604
rect 37651 11564 37663 11598
rect 37697 11595 37709 11598
rect 38512 11595 38518 11607
rect 37697 11567 38518 11595
rect 37697 11564 37709 11567
rect 37651 11558 37709 11564
rect 38512 11555 38518 11567
rect 38570 11555 38576 11607
rect 52528 11555 52534 11607
rect 52586 11595 52592 11607
rect 54640 11595 54646 11607
rect 52586 11567 54494 11595
rect 54601 11567 54646 11595
rect 52586 11555 52592 11567
rect 54466 11521 54494 11567
rect 54640 11555 54646 11567
rect 54698 11555 54704 11607
rect 56563 11598 56621 11604
rect 56563 11595 56575 11598
rect 54754 11567 56575 11595
rect 54754 11521 54782 11567
rect 56563 11564 56575 11567
rect 56609 11564 56621 11598
rect 57586 11595 57614 11715
rect 58192 11595 58198 11607
rect 57586 11567 58198 11595
rect 56563 11558 56621 11564
rect 58192 11555 58198 11567
rect 58250 11555 58256 11607
rect 54466 11493 54782 11521
rect 57136 11407 57142 11459
rect 57194 11447 57200 11459
rect 57331 11450 57389 11456
rect 57331 11447 57343 11450
rect 57194 11419 57343 11447
rect 57194 11407 57200 11419
rect 57331 11416 57343 11419
rect 57377 11416 57389 11450
rect 57331 11410 57389 11416
rect 1152 11348 58848 11370
rect 1152 11296 19654 11348
rect 19706 11296 19718 11348
rect 19770 11296 19782 11348
rect 19834 11296 19846 11348
rect 19898 11296 50374 11348
rect 50426 11296 50438 11348
rect 50490 11296 50502 11348
rect 50554 11296 50566 11348
rect 50618 11296 58848 11348
rect 1152 11274 58848 11296
rect 8656 11185 8662 11237
rect 8714 11225 8720 11237
rect 16048 11225 16054 11237
rect 8714 11197 16054 11225
rect 8714 11185 8720 11197
rect 16048 11185 16054 11197
rect 16106 11185 16112 11237
rect 21328 11037 21334 11089
rect 21386 11077 21392 11089
rect 55795 11080 55853 11086
rect 21386 11049 47534 11077
rect 21386 11037 21392 11049
rect 8080 10963 8086 11015
rect 8138 11003 8144 11015
rect 24208 11003 24214 11015
rect 8138 10975 24214 11003
rect 8138 10963 8144 10975
rect 24208 10963 24214 10975
rect 24266 10963 24272 11015
rect 24496 10963 24502 11015
rect 24554 11003 24560 11015
rect 33808 11003 33814 11015
rect 24554 10975 33814 11003
rect 24554 10963 24560 10975
rect 33808 10963 33814 10975
rect 33866 10963 33872 11015
rect 47506 11003 47534 11049
rect 55795 11046 55807 11080
rect 55841 11077 55853 11080
rect 55987 11080 56045 11086
rect 55987 11077 55999 11080
rect 55841 11049 55999 11077
rect 55841 11046 55853 11049
rect 55795 11040 55853 11046
rect 55987 11046 55999 11049
rect 56033 11077 56045 11080
rect 56080 11077 56086 11089
rect 56033 11049 56086 11077
rect 56033 11046 56045 11049
rect 55987 11040 56045 11046
rect 56080 11037 56086 11049
rect 56138 11077 56144 11089
rect 56275 11080 56333 11086
rect 56275 11077 56287 11080
rect 56138 11049 56287 11077
rect 56138 11037 56144 11049
rect 56275 11046 56287 11049
rect 56321 11046 56333 11080
rect 56275 11040 56333 11046
rect 56947 11006 57005 11012
rect 56947 11003 56959 11006
rect 47506 10975 56959 11003
rect 56947 10972 56959 10975
rect 56993 11003 57005 11006
rect 57235 11006 57293 11012
rect 57235 11003 57247 11006
rect 56993 10975 57247 11003
rect 56993 10972 57005 10975
rect 56947 10966 57005 10972
rect 57235 10972 57247 10975
rect 57281 10972 57293 11006
rect 57235 10966 57293 10972
rect 56083 10932 56141 10938
rect 56083 10898 56095 10932
rect 56129 10898 56141 10932
rect 56083 10892 56141 10898
rect 10576 10815 10582 10867
rect 10634 10855 10640 10867
rect 26800 10855 26806 10867
rect 10634 10827 26806 10855
rect 10634 10815 10640 10827
rect 26800 10815 26806 10827
rect 26858 10815 26864 10867
rect 28432 10815 28438 10867
rect 28490 10855 28496 10867
rect 29584 10855 29590 10867
rect 28490 10827 29590 10855
rect 28490 10815 28496 10827
rect 29584 10815 29590 10827
rect 29642 10815 29648 10867
rect 56098 10855 56126 10892
rect 56752 10889 56758 10941
rect 56810 10929 56816 10941
rect 57331 10932 57389 10938
rect 57331 10929 57343 10932
rect 56810 10901 57343 10929
rect 56810 10889 56816 10901
rect 57331 10898 57343 10901
rect 57377 10898 57389 10932
rect 57331 10892 57389 10898
rect 58288 10855 58294 10867
rect 56098 10827 58294 10855
rect 58288 10815 58294 10827
rect 58346 10815 58352 10867
rect 10864 10741 10870 10793
rect 10922 10781 10928 10793
rect 11152 10781 11158 10793
rect 10922 10753 11158 10781
rect 10922 10741 10928 10753
rect 11152 10741 11158 10753
rect 11210 10741 11216 10793
rect 12115 10784 12173 10790
rect 12115 10750 12127 10784
rect 12161 10781 12173 10784
rect 36016 10781 36022 10793
rect 12161 10753 36022 10781
rect 12161 10750 12173 10753
rect 12115 10744 12173 10750
rect 36016 10741 36022 10753
rect 36074 10741 36080 10793
rect 40720 10741 40726 10793
rect 40778 10781 40784 10793
rect 50896 10781 50902 10793
rect 40778 10753 50902 10781
rect 40778 10741 40784 10753
rect 50896 10741 50902 10753
rect 50954 10741 50960 10793
rect 1152 10682 58848 10704
rect 1152 10630 4294 10682
rect 4346 10630 4358 10682
rect 4410 10630 4422 10682
rect 4474 10630 4486 10682
rect 4538 10630 35014 10682
rect 35066 10630 35078 10682
rect 35130 10630 35142 10682
rect 35194 10630 35206 10682
rect 35258 10630 58848 10682
rect 1152 10608 58848 10630
rect 7603 10562 7661 10568
rect 7603 10528 7615 10562
rect 7649 10559 7661 10562
rect 56371 10562 56429 10568
rect 7649 10531 7934 10559
rect 7649 10528 7661 10531
rect 7603 10522 7661 10528
rect 7906 10485 7934 10531
rect 56371 10528 56383 10562
rect 56417 10559 56429 10562
rect 56848 10559 56854 10571
rect 56417 10531 56854 10559
rect 56417 10528 56429 10531
rect 56371 10522 56429 10528
rect 56848 10519 56854 10531
rect 56906 10519 56912 10571
rect 10576 10485 10582 10497
rect 7906 10457 10582 10485
rect 10576 10445 10582 10457
rect 10634 10445 10640 10497
rect 57043 10488 57101 10494
rect 57043 10485 57055 10488
rect 47506 10457 57055 10485
rect 12880 10371 12886 10423
rect 12938 10411 12944 10423
rect 47506 10411 47534 10457
rect 57043 10454 57055 10457
rect 57089 10485 57101 10488
rect 57089 10457 57374 10485
rect 57089 10454 57101 10457
rect 57043 10448 57101 10454
rect 12938 10383 47534 10411
rect 55027 10414 55085 10420
rect 12938 10371 12944 10383
rect 55027 10380 55039 10414
rect 55073 10380 55085 10414
rect 55027 10374 55085 10380
rect 55123 10414 55181 10420
rect 55123 10380 55135 10414
rect 55169 10411 55181 10414
rect 55984 10411 55990 10423
rect 55169 10383 55990 10411
rect 55169 10380 55181 10383
rect 55123 10374 55181 10380
rect 25168 10297 25174 10349
rect 25226 10337 25232 10349
rect 29203 10340 29261 10346
rect 29203 10337 29215 10340
rect 25226 10309 29215 10337
rect 25226 10297 25232 10309
rect 29203 10306 29215 10309
rect 29249 10306 29261 10340
rect 55042 10337 55070 10374
rect 55984 10371 55990 10383
rect 56042 10371 56048 10423
rect 56080 10371 56086 10423
rect 56138 10411 56144 10423
rect 57346 10420 57374 10457
rect 56659 10414 56717 10420
rect 56659 10411 56671 10414
rect 56138 10383 56671 10411
rect 56138 10371 56144 10383
rect 56659 10380 56671 10383
rect 56705 10380 56717 10414
rect 56659 10374 56717 10380
rect 57331 10414 57389 10420
rect 57331 10380 57343 10414
rect 57377 10380 57389 10414
rect 57331 10374 57389 10380
rect 55042 10309 57614 10337
rect 29203 10300 29261 10306
rect 26608 10223 26614 10275
rect 26666 10263 26672 10275
rect 28435 10266 28493 10272
rect 28435 10263 28447 10266
rect 26666 10235 28447 10263
rect 26666 10223 26672 10235
rect 28435 10232 28447 10235
rect 28481 10232 28493 10266
rect 28435 10226 28493 10232
rect 41491 10266 41549 10272
rect 41491 10232 41503 10266
rect 41537 10263 41549 10266
rect 51568 10263 51574 10275
rect 41537 10235 51574 10263
rect 41537 10232 41549 10235
rect 41491 10226 41549 10232
rect 51568 10223 51574 10235
rect 51626 10223 51632 10275
rect 55795 10266 55853 10272
rect 55795 10232 55807 10266
rect 55841 10232 55853 10266
rect 55795 10226 55853 10232
rect 56563 10266 56621 10272
rect 56563 10232 56575 10266
rect 56609 10263 56621 10266
rect 56848 10263 56854 10275
rect 56609 10235 56854 10263
rect 56609 10232 56621 10235
rect 56563 10226 56621 10232
rect 8080 10189 8086 10201
rect 7968 10161 8086 10189
rect 8080 10149 8086 10161
rect 8138 10149 8144 10201
rect 16240 10149 16246 10201
rect 16298 10189 16304 10201
rect 55507 10192 55565 10198
rect 55507 10189 55519 10192
rect 16298 10161 55519 10189
rect 16298 10149 16304 10161
rect 55507 10158 55519 10161
rect 55553 10189 55565 10192
rect 55810 10189 55838 10226
rect 56848 10223 56854 10235
rect 56906 10223 56912 10275
rect 55553 10161 55838 10189
rect 55553 10158 55565 10161
rect 55507 10152 55565 10158
rect 9424 10075 9430 10127
rect 9482 10115 9488 10127
rect 17104 10115 17110 10127
rect 9482 10087 17110 10115
rect 9482 10075 9488 10087
rect 17104 10075 17110 10087
rect 17162 10075 17168 10127
rect 55696 10075 55702 10127
rect 55754 10115 55760 10127
rect 55891 10118 55949 10124
rect 55891 10115 55903 10118
rect 55754 10087 55903 10115
rect 55754 10075 55760 10087
rect 55891 10084 55903 10087
rect 55937 10084 55949 10118
rect 55891 10078 55949 10084
rect 56464 10075 56470 10127
rect 56522 10115 56528 10127
rect 57427 10118 57485 10124
rect 57427 10115 57439 10118
rect 56522 10087 57439 10115
rect 56522 10075 56528 10087
rect 57427 10084 57439 10087
rect 57473 10084 57485 10118
rect 57586 10115 57614 10309
rect 58576 10115 58582 10127
rect 57586 10087 58582 10115
rect 57427 10078 57485 10084
rect 58576 10075 58582 10087
rect 58634 10075 58640 10127
rect 1152 10016 58848 10038
rect 1152 9964 19654 10016
rect 19706 9964 19718 10016
rect 19770 9964 19782 10016
rect 19834 9964 19846 10016
rect 19898 9964 50374 10016
rect 50426 9964 50438 10016
rect 50490 9964 50502 10016
rect 50554 9964 50566 10016
rect 50618 9964 58848 10016
rect 1152 9942 58848 9964
rect 8080 9853 8086 9905
rect 8138 9893 8144 9905
rect 17968 9893 17974 9905
rect 8138 9865 17974 9893
rect 8138 9853 8144 9865
rect 17968 9853 17974 9865
rect 18026 9853 18032 9905
rect 18352 9853 18358 9905
rect 18410 9893 18416 9905
rect 21520 9893 21526 9905
rect 18410 9865 21526 9893
rect 18410 9853 18416 9865
rect 21520 9853 21526 9865
rect 21578 9853 21584 9905
rect 42832 9893 42838 9905
rect 21634 9865 42838 9893
rect 7984 9779 7990 9831
rect 8042 9819 8048 9831
rect 10960 9819 10966 9831
rect 8042 9791 10966 9819
rect 8042 9779 8048 9791
rect 10960 9779 10966 9791
rect 11018 9779 11024 9831
rect 20368 9779 20374 9831
rect 20426 9819 20432 9831
rect 21634 9819 21662 9865
rect 42832 9853 42838 9865
rect 42890 9853 42896 9905
rect 55120 9853 55126 9905
rect 55178 9893 55184 9905
rect 55891 9896 55949 9902
rect 55891 9893 55903 9896
rect 55178 9865 55903 9893
rect 55178 9853 55184 9865
rect 55891 9862 55903 9865
rect 55937 9862 55949 9896
rect 55891 9856 55949 9862
rect 20426 9791 21662 9819
rect 20426 9779 20432 9791
rect 21712 9779 21718 9831
rect 21770 9819 21776 9831
rect 49168 9819 49174 9831
rect 21770 9791 49174 9819
rect 21770 9779 21776 9791
rect 49168 9779 49174 9791
rect 49226 9779 49232 9831
rect 51664 9779 51670 9831
rect 51722 9819 51728 9831
rect 51722 9791 56030 9819
rect 51722 9779 51728 9791
rect 20848 9705 20854 9757
rect 20906 9745 20912 9757
rect 54640 9745 54646 9757
rect 20906 9717 54646 9745
rect 20906 9705 20912 9717
rect 54640 9705 54646 9717
rect 54698 9705 54704 9757
rect 56002 9754 56030 9791
rect 55987 9748 56045 9754
rect 55987 9714 55999 9748
rect 56033 9714 56045 9748
rect 55987 9708 56045 9714
rect 8272 9631 8278 9683
rect 8330 9671 8336 9683
rect 16144 9671 16150 9683
rect 8330 9643 16150 9671
rect 8330 9631 8336 9643
rect 16144 9631 16150 9643
rect 16202 9631 16208 9683
rect 17296 9631 17302 9683
rect 17354 9671 17360 9683
rect 44656 9671 44662 9683
rect 17354 9643 44662 9671
rect 17354 9631 17360 9643
rect 44656 9631 44662 9643
rect 44714 9631 44720 9683
rect 46960 9631 46966 9683
rect 47018 9671 47024 9683
rect 55219 9674 55277 9680
rect 55219 9671 55231 9674
rect 47018 9643 55231 9671
rect 47018 9631 47024 9643
rect 55219 9640 55231 9643
rect 55265 9640 55277 9674
rect 55219 9634 55277 9640
rect 57616 9631 57622 9683
rect 57674 9671 57680 9683
rect 57674 9643 57719 9671
rect 57674 9631 57680 9643
rect 18256 9557 18262 9609
rect 18314 9597 18320 9609
rect 28240 9597 28246 9609
rect 18314 9569 28246 9597
rect 18314 9557 18320 9569
rect 28240 9557 28246 9569
rect 28298 9557 28304 9609
rect 28336 9557 28342 9609
rect 28394 9597 28400 9609
rect 29488 9597 29494 9609
rect 28394 9569 29494 9597
rect 28394 9557 28400 9569
rect 29488 9557 29494 9569
rect 29546 9557 29552 9609
rect 54256 9557 54262 9609
rect 54314 9597 54320 9609
rect 54355 9600 54413 9606
rect 54355 9597 54367 9600
rect 54314 9569 54367 9597
rect 54314 9557 54320 9569
rect 54355 9566 54367 9569
rect 54401 9566 54413 9600
rect 54355 9560 54413 9566
rect 54451 9600 54509 9606
rect 54451 9566 54463 9600
rect 54497 9566 54509 9600
rect 54451 9560 54509 9566
rect 15088 9483 15094 9535
rect 15146 9523 15152 9535
rect 43600 9523 43606 9535
rect 15146 9495 43606 9523
rect 15146 9483 15152 9495
rect 43600 9483 43606 9495
rect 43658 9483 43664 9535
rect 7792 9409 7798 9461
rect 7850 9449 7856 9461
rect 12208 9449 12214 9461
rect 7850 9421 12214 9449
rect 7850 9409 7856 9421
rect 12208 9409 12214 9421
rect 12266 9409 12272 9461
rect 16528 9409 16534 9461
rect 16586 9449 16592 9461
rect 20656 9449 20662 9461
rect 16586 9421 20662 9449
rect 16586 9409 16592 9421
rect 20656 9409 20662 9421
rect 20714 9409 20720 9461
rect 25840 9449 25846 9461
rect 25801 9421 25846 9449
rect 25840 9409 25846 9421
rect 25898 9409 25904 9461
rect 32371 9452 32429 9458
rect 32371 9418 32383 9452
rect 32417 9449 32429 9452
rect 34480 9449 34486 9461
rect 32417 9421 34486 9449
rect 32417 9418 32429 9421
rect 32371 9412 32429 9418
rect 34480 9409 34486 9421
rect 34538 9409 34544 9461
rect 35440 9409 35446 9461
rect 35498 9449 35504 9461
rect 41776 9449 41782 9461
rect 35498 9421 41782 9449
rect 35498 9409 35504 9421
rect 41776 9409 41782 9421
rect 41834 9409 41840 9461
rect 47728 9409 47734 9461
rect 47786 9449 47792 9461
rect 54466 9449 54494 9560
rect 54928 9557 54934 9609
rect 54986 9597 54992 9609
rect 55123 9600 55181 9606
rect 55123 9597 55135 9600
rect 54986 9569 55135 9597
rect 54986 9557 54992 9569
rect 55123 9566 55135 9569
rect 55169 9566 55181 9600
rect 55123 9560 55181 9566
rect 47786 9421 54494 9449
rect 47786 9409 47792 9421
rect 1152 9350 58848 9372
rect 1152 9298 4294 9350
rect 4346 9298 4358 9350
rect 4410 9298 4422 9350
rect 4474 9298 4486 9350
rect 4538 9298 35014 9350
rect 35066 9298 35078 9350
rect 35130 9298 35142 9350
rect 35194 9298 35206 9350
rect 35258 9298 58848 9350
rect 1152 9276 58848 9298
rect 7888 9227 7894 9239
rect 5746 9199 7894 9227
rect 5299 9156 5357 9162
rect 5299 9122 5311 9156
rect 5345 9153 5357 9156
rect 5587 9156 5645 9162
rect 5587 9153 5599 9156
rect 5345 9125 5599 9153
rect 5345 9122 5357 9125
rect 5299 9116 5357 9122
rect 5587 9122 5599 9125
rect 5633 9153 5645 9156
rect 5746 9153 5774 9199
rect 7888 9187 7894 9199
rect 7946 9187 7952 9239
rect 13936 9187 13942 9239
rect 13994 9227 14000 9239
rect 32944 9227 32950 9239
rect 13994 9199 32950 9227
rect 13994 9187 14000 9199
rect 32944 9187 32950 9199
rect 33002 9187 33008 9239
rect 33040 9187 33046 9239
rect 33098 9227 33104 9239
rect 51664 9227 51670 9239
rect 33098 9199 51670 9227
rect 33098 9187 33104 9199
rect 51664 9187 51670 9199
rect 51722 9187 51728 9239
rect 53008 9227 53014 9239
rect 52969 9199 53014 9227
rect 53008 9187 53014 9199
rect 53066 9187 53072 9239
rect 55123 9230 55181 9236
rect 55123 9196 55135 9230
rect 55169 9227 55181 9230
rect 55600 9227 55606 9239
rect 55169 9199 55606 9227
rect 55169 9196 55181 9199
rect 55123 9190 55181 9196
rect 5633 9125 5774 9153
rect 5633 9122 5645 9125
rect 5587 9116 5645 9122
rect 16432 9113 16438 9165
rect 16490 9153 16496 9165
rect 26800 9153 26806 9165
rect 16490 9125 26806 9153
rect 16490 9113 16496 9125
rect 26800 9113 26806 9125
rect 26858 9113 26864 9165
rect 28720 9113 28726 9165
rect 28778 9153 28784 9165
rect 36304 9153 36310 9165
rect 28778 9125 36310 9153
rect 28778 9113 28784 9125
rect 36304 9113 36310 9125
rect 36362 9113 36368 9165
rect 7968 9051 8126 9079
rect 8098 9017 8126 9051
rect 8512 9039 8518 9091
rect 8570 9039 8576 9091
rect 10768 9079 10774 9091
rect 8832 9051 10774 9079
rect 10768 9039 10774 9051
rect 10826 9039 10832 9091
rect 17680 9039 17686 9091
rect 17738 9079 17744 9091
rect 21712 9079 21718 9091
rect 17738 9051 21718 9079
rect 17738 9039 17744 9051
rect 21712 9039 21718 9051
rect 21770 9039 21776 9091
rect 53026 9079 53054 9187
rect 53299 9082 53357 9088
rect 53299 9079 53311 9082
rect 53026 9051 53311 9079
rect 53299 9048 53311 9051
rect 53345 9048 53357 9082
rect 53299 9042 53357 9048
rect 53395 9082 53453 9088
rect 53395 9048 53407 9082
rect 53441 9048 53453 9082
rect 53395 9042 53453 9048
rect 8230 9017 8282 9023
rect 8080 8965 8086 9017
rect 8138 8965 8144 9017
rect 8944 8965 8950 9017
rect 9002 9005 9008 9017
rect 19312 9005 19318 9017
rect 9002 8977 19318 9005
rect 9002 8965 9008 8977
rect 19312 8965 19318 8977
rect 19370 8965 19376 9017
rect 53410 9005 53438 9042
rect 54544 9039 54550 9091
rect 54602 9079 54608 9091
rect 55411 9082 55469 9088
rect 55411 9079 55423 9082
rect 54602 9051 55423 9079
rect 54602 9039 54608 9051
rect 55411 9048 55423 9051
rect 55457 9048 55469 9082
rect 55411 9042 55469 9048
rect 55216 9005 55222 9017
rect 53410 8977 55222 9005
rect 55216 8965 55222 8977
rect 55274 8965 55280 9017
rect 55315 9008 55373 9014
rect 55315 8974 55327 9008
rect 55361 9005 55373 9008
rect 55522 9005 55550 9199
rect 55600 9187 55606 9199
rect 55658 9187 55664 9239
rect 55361 8977 55550 9005
rect 56563 9008 56621 9014
rect 55361 8974 55373 8977
rect 55315 8968 55373 8974
rect 56563 8974 56575 9008
rect 56609 8974 56621 9008
rect 57232 9005 57238 9017
rect 57193 8977 57238 9005
rect 56563 8968 56621 8974
rect 8230 8959 8282 8965
rect 12688 8891 12694 8943
rect 12746 8931 12752 8943
rect 18448 8931 18454 8943
rect 12746 8903 18454 8931
rect 12746 8891 12752 8903
rect 18448 8891 18454 8903
rect 18506 8891 18512 8943
rect 25651 8934 25709 8940
rect 25651 8900 25663 8934
rect 25697 8931 25709 8934
rect 44080 8931 44086 8943
rect 25697 8903 44086 8931
rect 25697 8900 25709 8903
rect 25651 8894 25709 8900
rect 44080 8891 44086 8903
rect 44138 8891 44144 8943
rect 54547 8934 54605 8940
rect 54547 8900 54559 8934
rect 54593 8900 54605 8934
rect 56578 8931 56606 8968
rect 57232 8965 57238 8977
rect 57290 8965 57296 9017
rect 57328 8931 57334 8943
rect 56578 8903 57334 8931
rect 54547 8894 54605 8900
rect 16240 8817 16246 8869
rect 16298 8857 16304 8869
rect 18160 8857 18166 8869
rect 16298 8829 18166 8857
rect 16298 8817 16304 8829
rect 18160 8817 18166 8829
rect 18218 8817 18224 8869
rect 23152 8857 23158 8869
rect 20194 8829 23158 8857
rect 7600 8783 7606 8795
rect 7561 8755 7606 8783
rect 7600 8743 7606 8755
rect 7658 8743 7664 8795
rect 8848 8743 8854 8795
rect 8906 8743 8912 8795
rect 9040 8743 9046 8795
rect 9098 8783 9104 8795
rect 20194 8783 20222 8829
rect 23152 8817 23158 8829
rect 23210 8817 23216 8869
rect 26896 8817 26902 8869
rect 26954 8857 26960 8869
rect 54259 8860 54317 8866
rect 54259 8857 54271 8860
rect 26954 8829 37454 8857
rect 26954 8817 26960 8829
rect 9098 8755 20222 8783
rect 9098 8743 9104 8755
rect 20944 8743 20950 8795
rect 21002 8783 21008 8795
rect 22288 8783 22294 8795
rect 21002 8755 22294 8783
rect 21002 8743 21008 8755
rect 22288 8743 22294 8755
rect 22346 8743 22352 8795
rect 26992 8743 26998 8795
rect 27050 8783 27056 8795
rect 30160 8783 30166 8795
rect 27050 8755 30166 8783
rect 27050 8743 27056 8755
rect 30160 8743 30166 8755
rect 30218 8743 30224 8795
rect 37426 8783 37454 8829
rect 47506 8829 54271 8857
rect 47506 8783 47534 8829
rect 54259 8826 54271 8829
rect 54305 8857 54317 8860
rect 54562 8857 54590 8894
rect 57328 8891 57334 8903
rect 57386 8891 57392 8943
rect 54305 8829 54590 8857
rect 54305 8826 54317 8829
rect 54259 8820 54317 8826
rect 37426 8755 47534 8783
rect 53872 8743 53878 8795
rect 53930 8783 53936 8795
rect 54643 8786 54701 8792
rect 54643 8783 54655 8786
rect 53930 8755 54655 8783
rect 53930 8743 53936 8755
rect 54643 8752 54655 8755
rect 54689 8752 54701 8786
rect 54643 8746 54701 8752
rect 1152 8684 58848 8706
rect 1152 8632 19654 8684
rect 19706 8632 19718 8684
rect 19770 8632 19782 8684
rect 19834 8632 19846 8684
rect 19898 8632 50374 8684
rect 50426 8632 50438 8684
rect 50490 8632 50502 8684
rect 50554 8632 50566 8684
rect 50618 8632 58848 8684
rect 1152 8610 58848 8632
rect 1840 8561 1846 8573
rect 1762 8533 1846 8561
rect 1762 8422 1790 8533
rect 1840 8521 1846 8533
rect 1898 8561 1904 8573
rect 1939 8564 1997 8570
rect 1939 8561 1951 8564
rect 1898 8533 1951 8561
rect 1898 8521 1904 8533
rect 1939 8530 1951 8533
rect 1985 8530 1997 8564
rect 1939 8524 1997 8530
rect 5392 8521 5398 8573
rect 5450 8561 5456 8573
rect 7027 8564 7085 8570
rect 7027 8561 7039 8564
rect 5450 8533 7039 8561
rect 5450 8521 5456 8533
rect 7027 8530 7039 8533
rect 7073 8530 7085 8564
rect 7027 8524 7085 8530
rect 7600 8521 7606 8573
rect 7658 8561 7664 8573
rect 8848 8561 8854 8573
rect 7658 8533 8854 8561
rect 7658 8521 7664 8533
rect 8848 8521 8854 8533
rect 8906 8521 8912 8573
rect 9523 8564 9581 8570
rect 9523 8530 9535 8564
rect 9569 8561 9581 8564
rect 9904 8561 9910 8573
rect 9569 8533 9910 8561
rect 9569 8530 9581 8533
rect 9523 8524 9581 8530
rect 9904 8521 9910 8533
rect 9962 8561 9968 8573
rect 12592 8561 12598 8573
rect 9962 8533 12598 8561
rect 9962 8521 9968 8533
rect 12592 8521 12598 8533
rect 12650 8521 12656 8573
rect 12784 8521 12790 8573
rect 12842 8561 12848 8573
rect 13555 8564 13613 8570
rect 13555 8561 13567 8564
rect 12842 8533 13567 8561
rect 12842 8521 12848 8533
rect 13555 8530 13567 8533
rect 13601 8530 13613 8564
rect 48592 8561 48598 8573
rect 48553 8533 48598 8561
rect 13555 8524 13613 8530
rect 48592 8521 48598 8533
rect 48650 8561 48656 8573
rect 52435 8564 52493 8570
rect 48650 8533 48926 8561
rect 48650 8521 48656 8533
rect 4912 8447 4918 8499
rect 4970 8487 4976 8499
rect 4970 8459 47534 8487
rect 4970 8447 4976 8459
rect 1747 8416 1805 8422
rect 1747 8382 1759 8416
rect 1793 8382 1805 8416
rect 2512 8413 2518 8425
rect 2473 8385 2518 8413
rect 1747 8376 1805 8382
rect 2512 8373 2518 8385
rect 2570 8373 2576 8425
rect 5104 8373 5110 8425
rect 5162 8413 5168 8425
rect 7216 8413 7222 8425
rect 5162 8385 7222 8413
rect 5162 8373 5168 8385
rect 7216 8373 7222 8385
rect 7274 8373 7280 8425
rect 7603 8416 7661 8422
rect 7603 8382 7615 8416
rect 7649 8413 7661 8416
rect 7891 8416 7949 8422
rect 7891 8413 7903 8416
rect 7649 8385 7903 8413
rect 7649 8382 7661 8385
rect 7603 8376 7661 8382
rect 7891 8382 7903 8385
rect 7937 8413 7949 8416
rect 7984 8413 7990 8425
rect 7937 8385 7990 8413
rect 7937 8382 7949 8385
rect 7891 8376 7949 8382
rect 7984 8373 7990 8385
rect 8042 8373 8048 8425
rect 8080 8373 8086 8425
rect 8138 8413 8144 8425
rect 9712 8413 9718 8425
rect 8138 8385 9718 8413
rect 8138 8373 8144 8385
rect 9712 8373 9718 8385
rect 9770 8373 9776 8425
rect 9811 8416 9869 8422
rect 9811 8382 9823 8416
rect 9857 8413 9869 8416
rect 9904 8413 9910 8425
rect 9857 8385 9910 8413
rect 9857 8382 9869 8385
rect 9811 8376 9869 8382
rect 9904 8373 9910 8385
rect 9962 8373 9968 8425
rect 11059 8416 11117 8422
rect 11059 8382 11071 8416
rect 11105 8413 11117 8416
rect 11344 8413 11350 8425
rect 11105 8385 11350 8413
rect 11105 8382 11117 8385
rect 11059 8376 11117 8382
rect 11344 8373 11350 8385
rect 11402 8373 11408 8425
rect 13552 8373 13558 8425
rect 13610 8413 13616 8425
rect 13651 8416 13709 8422
rect 13651 8413 13663 8416
rect 13610 8385 13663 8413
rect 13610 8373 13616 8385
rect 13651 8382 13663 8385
rect 13697 8382 13709 8416
rect 16240 8413 16246 8425
rect 16201 8385 16246 8413
rect 13651 8376 13709 8382
rect 16240 8373 16246 8385
rect 16298 8373 16304 8425
rect 17008 8413 17014 8425
rect 16969 8385 17014 8413
rect 17008 8373 17014 8385
rect 17066 8373 17072 8425
rect 38419 8416 38477 8422
rect 38419 8413 38431 8416
rect 17266 8385 38431 8413
rect 3283 8342 3341 8348
rect 3283 8308 3295 8342
rect 3329 8339 3341 8342
rect 7027 8342 7085 8348
rect 3329 8311 6974 8339
rect 3329 8308 3341 8311
rect 3283 8302 3341 8308
rect 1648 8265 1654 8277
rect 1609 8237 1654 8265
rect 1648 8225 1654 8237
rect 1706 8225 1712 8277
rect 2128 8225 2134 8277
rect 2186 8265 2192 8277
rect 2419 8268 2477 8274
rect 2419 8265 2431 8268
rect 2186 8237 2431 8265
rect 2186 8225 2192 8237
rect 2419 8234 2431 8237
rect 2465 8234 2477 8268
rect 3184 8265 3190 8277
rect 3145 8237 3190 8265
rect 2419 8228 2477 8234
rect 3184 8225 3190 8237
rect 3242 8225 3248 8277
rect 4435 8268 4493 8274
rect 4435 8234 4447 8268
rect 4481 8234 4493 8268
rect 4435 8228 4493 8234
rect 4531 8268 4589 8274
rect 4531 8234 4543 8268
rect 4577 8265 4589 8268
rect 6832 8265 6838 8277
rect 4577 8237 6838 8265
rect 4577 8234 4589 8237
rect 4531 8228 4589 8234
rect 4450 8191 4478 8228
rect 4816 8191 4822 8203
rect 4450 8163 4822 8191
rect 4816 8151 4822 8163
rect 4874 8151 4880 8203
rect 4243 8120 4301 8126
rect 4243 8086 4255 8120
rect 4289 8117 4301 8120
rect 4930 8117 4958 8237
rect 6832 8225 6838 8237
rect 6890 8225 6896 8277
rect 6946 8191 6974 8311
rect 7027 8308 7039 8342
rect 7073 8339 7085 8342
rect 12115 8342 12173 8348
rect 12115 8339 12127 8342
rect 7073 8311 12127 8339
rect 7073 8308 7085 8311
rect 7027 8302 7085 8308
rect 12115 8308 12127 8311
rect 12161 8308 12173 8342
rect 12115 8302 12173 8308
rect 12883 8342 12941 8348
rect 12883 8308 12895 8342
rect 12929 8339 12941 8342
rect 13744 8339 13750 8351
rect 12929 8311 13750 8339
rect 12929 8308 12941 8311
rect 12883 8302 12941 8308
rect 13744 8299 13750 8311
rect 13802 8299 13808 8351
rect 17266 8339 17294 8385
rect 38419 8382 38431 8385
rect 38465 8413 38477 8416
rect 38611 8416 38669 8422
rect 38611 8413 38623 8416
rect 38465 8385 38623 8413
rect 38465 8382 38477 8385
rect 38419 8376 38477 8382
rect 38611 8382 38623 8385
rect 38657 8382 38669 8416
rect 38611 8376 38669 8382
rect 15826 8311 17294 8339
rect 47506 8339 47534 8459
rect 47923 8416 47981 8422
rect 47923 8382 47935 8416
rect 47969 8413 47981 8416
rect 48112 8413 48118 8425
rect 47969 8385 48118 8413
rect 47969 8382 47981 8385
rect 47923 8376 47981 8382
rect 48112 8373 48118 8385
rect 48170 8373 48176 8425
rect 48898 8422 48926 8533
rect 52435 8530 52447 8564
rect 52481 8561 52493 8564
rect 58960 8561 58966 8573
rect 52481 8533 58966 8561
rect 52481 8530 52493 8533
rect 52435 8524 52493 8530
rect 58960 8521 58966 8533
rect 59018 8521 59024 8573
rect 48883 8416 48941 8422
rect 48883 8382 48895 8416
rect 48929 8382 48941 8416
rect 49744 8413 49750 8425
rect 49705 8385 49750 8413
rect 48883 8376 48941 8382
rect 49744 8373 49750 8385
rect 49802 8373 49808 8425
rect 51568 8373 51574 8425
rect 51626 8413 51632 8425
rect 52531 8416 52589 8422
rect 52531 8413 52543 8416
rect 51626 8385 52543 8413
rect 51626 8373 51632 8385
rect 52531 8382 52543 8385
rect 52577 8382 52589 8416
rect 52531 8376 52589 8382
rect 53011 8416 53069 8422
rect 53011 8382 53023 8416
rect 53057 8413 53069 8416
rect 53200 8413 53206 8425
rect 53057 8385 53206 8413
rect 53057 8382 53069 8385
rect 53011 8376 53069 8382
rect 53200 8373 53206 8385
rect 53258 8373 53264 8425
rect 54064 8413 54070 8425
rect 54025 8385 54070 8413
rect 54064 8373 54070 8385
rect 54122 8373 54128 8425
rect 51184 8339 51190 8351
rect 47506 8311 51190 8339
rect 7696 8225 7702 8277
rect 7754 8265 7760 8277
rect 7795 8268 7853 8274
rect 7795 8265 7807 8268
rect 7754 8237 7807 8265
rect 7754 8225 7760 8237
rect 7795 8234 7807 8237
rect 7841 8234 7853 8268
rect 7795 8228 7853 8234
rect 9520 8225 9526 8277
rect 9578 8265 9584 8277
rect 9715 8268 9773 8274
rect 9715 8265 9727 8268
rect 9578 8237 9727 8265
rect 9578 8225 9584 8237
rect 9715 8234 9727 8237
rect 9761 8234 9773 8268
rect 9715 8228 9773 8234
rect 10288 8225 10294 8277
rect 10346 8265 10352 8277
rect 10483 8268 10541 8274
rect 10483 8265 10495 8268
rect 10346 8237 10495 8265
rect 10346 8225 10352 8237
rect 10483 8234 10495 8237
rect 10529 8234 10541 8268
rect 10483 8228 10541 8234
rect 10579 8268 10637 8274
rect 10579 8234 10591 8268
rect 10625 8234 10637 8268
rect 10579 8228 10637 8234
rect 10195 8194 10253 8200
rect 6946 8163 9566 8191
rect 5488 8117 5494 8129
rect 4289 8089 4958 8117
rect 5449 8089 5494 8117
rect 4289 8086 4301 8089
rect 4243 8080 4301 8086
rect 5488 8077 5494 8089
rect 5546 8077 5552 8129
rect 9538 8117 9566 8163
rect 10195 8160 10207 8194
rect 10241 8191 10253 8194
rect 10594 8191 10622 8228
rect 10672 8225 10678 8277
rect 10730 8265 10736 8277
rect 11251 8268 11309 8274
rect 11251 8265 11263 8268
rect 10730 8237 11263 8265
rect 10730 8225 10736 8237
rect 11251 8234 11263 8237
rect 11297 8234 11309 8268
rect 11251 8228 11309 8234
rect 11440 8225 11446 8277
rect 11498 8265 11504 8277
rect 12019 8268 12077 8274
rect 12019 8265 12031 8268
rect 11498 8237 12031 8265
rect 11498 8225 11504 8237
rect 12019 8234 12031 8237
rect 12065 8234 12077 8268
rect 12019 8228 12077 8234
rect 12208 8225 12214 8277
rect 12266 8265 12272 8277
rect 12787 8268 12845 8274
rect 12787 8265 12799 8268
rect 12266 8237 12799 8265
rect 12266 8225 12272 8237
rect 12787 8234 12799 8237
rect 12833 8234 12845 8268
rect 15826 8265 15854 8311
rect 51184 8299 51190 8311
rect 51242 8299 51248 8351
rect 55219 8342 55277 8348
rect 55219 8308 55231 8342
rect 55265 8339 55277 8342
rect 55987 8342 56045 8348
rect 55265 8311 55934 8339
rect 55265 8308 55277 8311
rect 55219 8302 55277 8308
rect 12787 8228 12845 8234
rect 13666 8237 15854 8265
rect 13666 8191 13694 8237
rect 16048 8225 16054 8277
rect 16106 8265 16112 8277
rect 16147 8268 16205 8274
rect 16147 8265 16159 8268
rect 16106 8237 16159 8265
rect 16106 8225 16112 8237
rect 16147 8234 16159 8237
rect 16193 8234 16205 8268
rect 16147 8228 16205 8234
rect 16336 8225 16342 8277
rect 16394 8265 16400 8277
rect 16915 8268 16973 8274
rect 16915 8265 16927 8268
rect 16394 8237 16927 8265
rect 16394 8225 16400 8237
rect 16915 8234 16927 8237
rect 16961 8234 16973 8268
rect 16915 8228 16973 8234
rect 48211 8268 48269 8274
rect 48211 8234 48223 8268
rect 48257 8234 48269 8268
rect 48211 8228 48269 8234
rect 25651 8194 25709 8200
rect 25651 8191 25663 8194
rect 10241 8163 13694 8191
rect 15826 8163 25663 8191
rect 10241 8160 10253 8163
rect 10195 8154 10253 8160
rect 15826 8117 15854 8163
rect 25651 8160 25663 8163
rect 25697 8160 25709 8194
rect 25651 8154 25709 8160
rect 48016 8151 48022 8203
rect 48074 8191 48080 8203
rect 48226 8191 48254 8228
rect 48688 8225 48694 8277
rect 48746 8265 48752 8277
rect 48979 8268 49037 8274
rect 48979 8265 48991 8268
rect 48746 8237 48991 8265
rect 48746 8225 48752 8237
rect 48979 8234 48991 8237
rect 49025 8234 49037 8268
rect 48979 8228 49037 8234
rect 49456 8225 49462 8277
rect 49514 8265 49520 8277
rect 49651 8268 49709 8274
rect 49651 8265 49663 8268
rect 49514 8237 49663 8265
rect 49514 8225 49520 8237
rect 49651 8234 49663 8237
rect 49697 8234 49709 8268
rect 49651 8228 49709 8234
rect 53299 8268 53357 8274
rect 53299 8234 53311 8268
rect 53345 8234 53357 8268
rect 53299 8228 53357 8234
rect 48074 8163 48254 8191
rect 48074 8151 48080 8163
rect 53104 8151 53110 8203
rect 53162 8191 53168 8203
rect 53314 8191 53342 8228
rect 53488 8225 53494 8277
rect 53546 8265 53552 8277
rect 53971 8268 54029 8274
rect 53971 8265 53983 8268
rect 53546 8237 53983 8265
rect 53546 8225 53552 8237
rect 53971 8234 53983 8237
rect 54017 8234 54029 8268
rect 53971 8228 54029 8234
rect 53162 8163 53342 8191
rect 55906 8191 55934 8311
rect 55987 8308 55999 8342
rect 56033 8308 56045 8342
rect 55987 8302 56045 8308
rect 56002 8265 56030 8302
rect 56944 8299 56950 8351
rect 57002 8339 57008 8351
rect 57139 8342 57197 8348
rect 57139 8339 57151 8342
rect 57002 8311 57151 8339
rect 57002 8299 57008 8311
rect 57139 8308 57151 8311
rect 57185 8308 57197 8342
rect 57139 8302 57197 8308
rect 58384 8265 58390 8277
rect 56002 8237 58390 8265
rect 58384 8225 58390 8237
rect 58442 8225 58448 8277
rect 59824 8191 59830 8203
rect 55906 8163 59830 8191
rect 53162 8151 53168 8163
rect 59824 8151 59830 8163
rect 59882 8151 59888 8203
rect 9538 8089 15854 8117
rect 16240 8077 16246 8129
rect 16298 8117 16304 8129
rect 18355 8120 18413 8126
rect 18355 8117 18367 8120
rect 16298 8089 18367 8117
rect 16298 8077 16304 8089
rect 18355 8086 18367 8089
rect 18401 8086 18413 8120
rect 18355 8080 18413 8086
rect 29587 8120 29645 8126
rect 29587 8086 29599 8120
rect 29633 8117 29645 8120
rect 31216 8117 31222 8129
rect 29633 8089 31222 8117
rect 29633 8086 29645 8089
rect 29587 8080 29645 8086
rect 31216 8077 31222 8089
rect 31274 8077 31280 8129
rect 44944 8077 44950 8129
rect 45002 8117 45008 8129
rect 45139 8120 45197 8126
rect 45139 8117 45151 8120
rect 45002 8089 45151 8117
rect 45002 8077 45008 8089
rect 45139 8086 45151 8089
rect 45185 8086 45197 8120
rect 45139 8080 45197 8086
rect 1152 8018 58848 8040
rect 1152 7966 4294 8018
rect 4346 7966 4358 8018
rect 4410 7966 4422 8018
rect 4474 7966 4486 8018
rect 4538 7966 35014 8018
rect 35066 7966 35078 8018
rect 35130 7966 35142 8018
rect 35194 7966 35206 8018
rect 35258 7966 58848 8018
rect 1152 7944 58848 7966
rect 8512 7855 8518 7907
rect 8570 7895 8576 7907
rect 11248 7895 11254 7907
rect 8570 7867 11254 7895
rect 8570 7855 8576 7867
rect 11248 7855 11254 7867
rect 11306 7855 11312 7907
rect 36496 7895 36502 7907
rect 36457 7867 36502 7895
rect 36496 7855 36502 7867
rect 36554 7855 36560 7907
rect 40819 7898 40877 7904
rect 40819 7864 40831 7898
rect 40865 7895 40877 7898
rect 41008 7895 41014 7907
rect 40865 7867 41014 7895
rect 40865 7864 40877 7867
rect 40819 7858 40877 7864
rect 41008 7855 41014 7867
rect 41066 7855 41072 7907
rect 42256 7895 42262 7907
rect 42217 7867 42262 7895
rect 42256 7855 42262 7867
rect 42314 7855 42320 7907
rect 45232 7895 45238 7907
rect 45193 7867 45238 7895
rect 45232 7855 45238 7867
rect 45290 7855 45296 7907
rect 46099 7898 46157 7904
rect 46099 7864 46111 7898
rect 46145 7895 46157 7898
rect 46192 7895 46198 7907
rect 46145 7867 46198 7895
rect 46145 7864 46157 7867
rect 46099 7858 46157 7864
rect 46192 7855 46198 7867
rect 46250 7855 46256 7907
rect 47536 7855 47542 7907
rect 47594 7895 47600 7907
rect 48976 7895 48982 7907
rect 47594 7867 47639 7895
rect 48937 7867 48982 7895
rect 47594 7855 47600 7867
rect 48976 7855 48982 7867
rect 49034 7855 49040 7907
rect 52912 7855 52918 7907
rect 52970 7895 52976 7907
rect 53011 7898 53069 7904
rect 53011 7895 53023 7898
rect 52970 7867 53023 7895
rect 52970 7855 52976 7867
rect 53011 7864 53023 7867
rect 53057 7864 53069 7898
rect 53011 7858 53069 7864
rect 2227 7824 2285 7830
rect 2227 7790 2239 7824
rect 2273 7821 2285 7824
rect 3760 7821 3766 7833
rect 2273 7793 3766 7821
rect 2273 7790 2285 7793
rect 2227 7784 2285 7790
rect 2530 7756 2558 7793
rect 3760 7781 3766 7793
rect 3818 7781 3824 7833
rect 7603 7824 7661 7830
rect 7603 7790 7615 7824
rect 7649 7821 7661 7824
rect 7792 7821 7798 7833
rect 7649 7793 7798 7821
rect 7649 7790 7661 7793
rect 7603 7784 7661 7790
rect 7792 7781 7798 7793
rect 7850 7781 7856 7833
rect 54160 7821 54166 7833
rect 27346 7793 54166 7821
rect 2515 7750 2573 7756
rect 2515 7716 2527 7750
rect 2561 7716 2573 7750
rect 2515 7710 2573 7716
rect 3283 7750 3341 7756
rect 3283 7716 3295 7750
rect 3329 7747 3341 7750
rect 5488 7747 5494 7759
rect 3329 7719 5494 7747
rect 3329 7716 3341 7719
rect 3283 7710 3341 7716
rect 5488 7707 5494 7719
rect 5546 7707 5552 7759
rect 7936 7707 7942 7759
rect 7994 7707 8000 7759
rect 9136 7707 9142 7759
rect 9194 7747 9200 7759
rect 10099 7750 10157 7756
rect 10099 7747 10111 7750
rect 9194 7719 10111 7747
rect 9194 7707 9200 7719
rect 10099 7716 10111 7719
rect 10145 7716 10157 7750
rect 10099 7710 10157 7716
rect 11728 7707 11734 7759
rect 11786 7747 11792 7759
rect 13075 7750 13133 7756
rect 13075 7747 13087 7750
rect 11786 7719 13087 7747
rect 11786 7707 11792 7719
rect 13075 7716 13087 7719
rect 13121 7716 13133 7750
rect 13075 7710 13133 7716
rect 13651 7750 13709 7756
rect 13651 7716 13663 7750
rect 13697 7747 13709 7750
rect 13939 7750 13997 7756
rect 13939 7747 13951 7750
rect 13697 7719 13951 7747
rect 13697 7716 13709 7719
rect 13651 7710 13709 7716
rect 13939 7716 13951 7719
rect 13985 7747 13997 7750
rect 20659 7750 20717 7756
rect 13985 7719 20606 7747
rect 13985 7716 13997 7719
rect 13939 7710 13997 7716
rect 8518 7685 8570 7691
rect 1456 7633 1462 7685
rect 1514 7673 1520 7685
rect 1555 7676 1613 7682
rect 1555 7673 1567 7676
rect 1514 7645 1567 7673
rect 1514 7633 1520 7645
rect 1555 7642 1567 7645
rect 1601 7642 1613 7676
rect 1555 7636 1613 7642
rect 3763 7676 3821 7682
rect 3763 7642 3775 7676
rect 3809 7673 3821 7676
rect 4048 7673 4054 7685
rect 3809 7645 4054 7673
rect 3809 7642 3821 7645
rect 3763 7636 3821 7642
rect 4048 7633 4054 7645
rect 4106 7633 4112 7685
rect 4819 7676 4877 7682
rect 4819 7642 4831 7676
rect 4865 7673 4877 7676
rect 4912 7673 4918 7685
rect 4865 7645 4918 7673
rect 4865 7642 4877 7645
rect 4819 7636 4877 7642
rect 4912 7633 4918 7645
rect 4970 7633 4976 7685
rect 9043 7676 9101 7682
rect 9043 7642 9055 7676
rect 9089 7673 9101 7676
rect 9424 7673 9430 7685
rect 9089 7645 9430 7673
rect 9089 7642 9101 7645
rect 9043 7636 9101 7642
rect 9424 7633 9430 7645
rect 9482 7633 9488 7685
rect 10195 7676 10253 7682
rect 10195 7642 10207 7676
rect 10241 7673 10253 7676
rect 12016 7673 12022 7685
rect 10241 7645 12022 7673
rect 10241 7642 10253 7645
rect 10195 7636 10253 7642
rect 12016 7633 12022 7645
rect 12074 7633 12080 7685
rect 12403 7676 12461 7682
rect 12403 7642 12415 7676
rect 12449 7673 12461 7676
rect 12496 7673 12502 7685
rect 12449 7645 12502 7673
rect 12449 7642 12461 7645
rect 12403 7636 12461 7642
rect 12496 7633 12502 7645
rect 12554 7633 12560 7685
rect 14803 7676 14861 7682
rect 14803 7642 14815 7676
rect 14849 7673 14861 7676
rect 15088 7673 15094 7685
rect 14849 7645 15094 7673
rect 14849 7642 14861 7645
rect 14803 7636 14861 7642
rect 15088 7633 15094 7645
rect 15146 7633 15152 7685
rect 15856 7673 15862 7685
rect 15817 7645 15862 7673
rect 15856 7633 15862 7645
rect 15914 7633 15920 7685
rect 20578 7673 20606 7719
rect 20659 7716 20671 7750
rect 20705 7747 20717 7750
rect 20944 7747 20950 7759
rect 20705 7719 20950 7747
rect 20705 7716 20717 7719
rect 20659 7710 20717 7716
rect 20944 7707 20950 7719
rect 21002 7707 21008 7759
rect 23635 7750 23693 7756
rect 23635 7716 23647 7750
rect 23681 7747 23693 7750
rect 23923 7750 23981 7756
rect 23923 7747 23935 7750
rect 23681 7719 23935 7747
rect 23681 7716 23693 7719
rect 23635 7710 23693 7716
rect 23923 7716 23935 7719
rect 23969 7747 23981 7750
rect 24016 7747 24022 7759
rect 23969 7719 24022 7747
rect 23969 7716 23981 7719
rect 23923 7710 23981 7716
rect 24016 7707 24022 7719
rect 24074 7707 24080 7759
rect 25456 7747 25462 7759
rect 25417 7719 25462 7747
rect 25456 7707 25462 7719
rect 25514 7707 25520 7759
rect 26224 7747 26230 7759
rect 26185 7719 26230 7747
rect 26224 7707 26230 7719
rect 26282 7707 26288 7759
rect 26992 7747 26998 7759
rect 26953 7719 26998 7747
rect 26992 7707 26998 7719
rect 27050 7707 27056 7759
rect 27346 7673 27374 7793
rect 54160 7781 54166 7793
rect 54218 7781 54224 7833
rect 28051 7750 28109 7756
rect 28051 7716 28063 7750
rect 28097 7747 28109 7750
rect 28339 7750 28397 7756
rect 28339 7747 28351 7750
rect 28097 7719 28351 7747
rect 28097 7716 28109 7719
rect 28051 7710 28109 7716
rect 28339 7716 28351 7719
rect 28385 7747 28397 7750
rect 28432 7747 28438 7759
rect 28385 7719 28438 7747
rect 28385 7716 28397 7719
rect 28339 7710 28397 7716
rect 28432 7707 28438 7719
rect 28490 7707 28496 7759
rect 29392 7747 29398 7759
rect 29353 7719 29398 7747
rect 29392 7707 29398 7719
rect 29450 7707 29456 7759
rect 29584 7707 29590 7759
rect 29642 7747 29648 7759
rect 30163 7750 30221 7756
rect 30163 7747 30175 7750
rect 29642 7719 30175 7747
rect 29642 7707 29648 7719
rect 30163 7716 30175 7719
rect 30209 7716 30221 7750
rect 31216 7747 31222 7759
rect 31177 7719 31222 7747
rect 30163 7710 30221 7716
rect 31216 7707 31222 7719
rect 31274 7707 31280 7759
rect 34576 7747 34582 7759
rect 34537 7719 34582 7747
rect 34576 7707 34582 7719
rect 34634 7707 34640 7759
rect 35344 7747 35350 7759
rect 35305 7719 35350 7747
rect 35344 7707 35350 7719
rect 35402 7707 35408 7759
rect 36112 7747 36118 7759
rect 36073 7719 36118 7747
rect 36112 7707 36118 7719
rect 36170 7707 36176 7759
rect 36496 7707 36502 7759
rect 36554 7747 36560 7759
rect 36787 7750 36845 7756
rect 36787 7747 36799 7750
rect 36554 7719 36799 7747
rect 36554 7707 36560 7719
rect 36787 7716 36799 7719
rect 36833 7716 36845 7750
rect 40336 7747 40342 7759
rect 40297 7719 40342 7747
rect 36787 7710 36845 7716
rect 40336 7707 40342 7719
rect 40394 7707 40400 7759
rect 41011 7750 41069 7756
rect 41011 7716 41023 7750
rect 41057 7716 41069 7750
rect 41872 7747 41878 7759
rect 41833 7719 41878 7747
rect 41011 7710 41069 7716
rect 20578 7645 27374 7673
rect 29875 7676 29933 7682
rect 29875 7642 29887 7676
rect 29921 7673 29933 7676
rect 30064 7673 30070 7685
rect 29921 7645 30070 7673
rect 29921 7642 29933 7645
rect 29875 7636 29933 7642
rect 30064 7633 30070 7645
rect 30122 7633 30128 7685
rect 40240 7633 40246 7685
rect 40298 7673 40304 7685
rect 41026 7673 41054 7710
rect 41872 7707 41878 7719
rect 41930 7707 41936 7759
rect 42256 7707 42262 7759
rect 42314 7747 42320 7759
rect 42547 7750 42605 7756
rect 42547 7747 42559 7750
rect 42314 7719 42559 7747
rect 42314 7707 42320 7719
rect 42547 7716 42559 7719
rect 42593 7716 42605 7750
rect 44080 7747 44086 7759
rect 44041 7719 44086 7747
rect 42547 7710 42605 7716
rect 44080 7707 44086 7719
rect 44138 7707 44144 7759
rect 44563 7750 44621 7756
rect 44563 7716 44575 7750
rect 44609 7747 44621 7750
rect 44848 7747 44854 7759
rect 44609 7719 44854 7747
rect 44609 7716 44621 7719
rect 44563 7710 44621 7716
rect 44848 7707 44854 7719
rect 44906 7707 44912 7759
rect 45040 7707 45046 7759
rect 45098 7747 45104 7759
rect 45619 7750 45677 7756
rect 45619 7747 45631 7750
rect 45098 7719 45631 7747
rect 45098 7707 45104 7719
rect 45619 7716 45631 7719
rect 45665 7716 45677 7750
rect 45619 7710 45677 7716
rect 45808 7707 45814 7759
rect 45866 7747 45872 7759
rect 46387 7750 46445 7756
rect 46387 7747 46399 7750
rect 45866 7719 46399 7747
rect 45866 7707 45872 7719
rect 46387 7716 46399 7719
rect 46433 7716 46445 7750
rect 47152 7747 47158 7759
rect 47113 7719 47158 7747
rect 46387 7710 46445 7716
rect 47152 7707 47158 7719
rect 47210 7707 47216 7759
rect 47536 7707 47542 7759
rect 47594 7747 47600 7759
rect 47827 7750 47885 7756
rect 47827 7747 47839 7750
rect 47594 7719 47839 7747
rect 47594 7707 47600 7719
rect 47827 7716 47839 7719
rect 47873 7716 47885 7750
rect 47827 7710 47885 7716
rect 48400 7707 48406 7759
rect 48458 7747 48464 7759
rect 49363 7750 49421 7756
rect 49363 7747 49375 7750
rect 48458 7719 49375 7747
rect 48458 7707 48464 7719
rect 49363 7716 49375 7719
rect 49409 7716 49421 7750
rect 49363 7710 49421 7716
rect 51571 7750 51629 7756
rect 51571 7716 51583 7750
rect 51617 7747 51629 7750
rect 51760 7747 51766 7759
rect 51617 7719 51766 7747
rect 51617 7716 51629 7719
rect 51571 7710 51629 7716
rect 51760 7707 51766 7719
rect 51818 7707 51824 7759
rect 52624 7747 52630 7759
rect 52585 7719 52630 7747
rect 52624 7707 52630 7719
rect 52682 7707 52688 7759
rect 52720 7707 52726 7759
rect 52778 7747 52784 7759
rect 53395 7750 53453 7756
rect 53395 7747 53407 7750
rect 52778 7719 53407 7747
rect 52778 7707 52784 7719
rect 53395 7716 53407 7719
rect 53441 7716 53453 7750
rect 58768 7747 58774 7759
rect 53395 7710 53453 7716
rect 55138 7719 58774 7747
rect 40298 7645 41054 7673
rect 40298 7633 40304 7645
rect 42160 7633 42166 7685
rect 42218 7673 42224 7685
rect 42218 7645 45662 7673
rect 42218 7633 42224 7645
rect 8518 7627 8570 7633
rect 5584 7599 5590 7611
rect 5545 7571 5590 7599
rect 5584 7559 5590 7571
rect 5642 7559 5648 7611
rect 8080 7559 8086 7611
rect 8138 7559 8144 7611
rect 10675 7602 10733 7608
rect 10675 7568 10687 7602
rect 10721 7599 10733 7602
rect 10963 7602 11021 7608
rect 10963 7599 10975 7602
rect 10721 7571 10975 7599
rect 10721 7568 10733 7571
rect 10675 7562 10733 7568
rect 10963 7568 10975 7571
rect 11009 7599 11021 7602
rect 12304 7599 12310 7611
rect 11009 7571 12310 7599
rect 11009 7568 11021 7571
rect 10963 7562 11021 7568
rect 12304 7559 12310 7571
rect 12362 7559 12368 7611
rect 13171 7602 13229 7608
rect 13171 7568 13183 7602
rect 13217 7568 13229 7602
rect 13171 7562 13229 7568
rect 8098 7525 8126 7559
rect 8098 7497 8256 7525
rect 9904 7485 9910 7537
rect 9962 7525 9968 7537
rect 13186 7525 13214 7562
rect 21232 7559 21238 7611
rect 21290 7599 21296 7611
rect 24691 7602 24749 7608
rect 24691 7599 24703 7602
rect 21290 7571 24703 7599
rect 21290 7559 21296 7571
rect 24691 7568 24703 7571
rect 24737 7568 24749 7602
rect 24691 7562 24749 7568
rect 33811 7602 33869 7608
rect 33811 7568 33823 7602
rect 33857 7599 33869 7602
rect 33904 7599 33910 7611
rect 33857 7571 33910 7599
rect 33857 7568 33869 7571
rect 33811 7562 33869 7568
rect 33904 7559 33910 7571
rect 33962 7559 33968 7611
rect 34480 7559 34486 7611
rect 34538 7599 34544 7611
rect 38803 7602 38861 7608
rect 38803 7599 38815 7602
rect 34538 7571 38815 7599
rect 34538 7559 34544 7571
rect 38803 7568 38815 7571
rect 38849 7568 38861 7602
rect 38803 7562 38861 7568
rect 39571 7602 39629 7608
rect 39571 7568 39583 7602
rect 39617 7568 39629 7602
rect 39571 7562 39629 7568
rect 22960 7525 22966 7537
rect 9962 7497 10910 7525
rect 13186 7497 22966 7525
rect 9962 7485 9968 7497
rect 2416 7451 2422 7463
rect 2377 7423 2422 7451
rect 2416 7411 2422 7423
rect 2474 7411 2480 7463
rect 2992 7411 2998 7463
rect 3050 7451 3056 7463
rect 3187 7454 3245 7460
rect 3187 7451 3199 7454
rect 3050 7423 3199 7451
rect 3050 7411 3056 7423
rect 3187 7420 3199 7423
rect 3233 7420 3245 7454
rect 3952 7451 3958 7463
rect 3913 7423 3958 7451
rect 3187 7414 3245 7420
rect 3952 7411 3958 7423
rect 4010 7411 4016 7463
rect 4048 7411 4054 7463
rect 4106 7451 4112 7463
rect 4723 7454 4781 7460
rect 4723 7451 4735 7454
rect 4106 7423 4735 7451
rect 4106 7411 4112 7423
rect 4723 7420 4735 7423
rect 4769 7420 4781 7454
rect 4723 7414 4781 7420
rect 5296 7411 5302 7463
rect 5354 7451 5360 7463
rect 5491 7454 5549 7460
rect 5491 7451 5503 7454
rect 5354 7423 5503 7451
rect 5354 7411 5360 7423
rect 5491 7420 5503 7423
rect 5537 7420 5549 7454
rect 9328 7451 9334 7463
rect 9289 7423 9334 7451
rect 5491 7414 5549 7420
rect 9328 7411 9334 7423
rect 9386 7411 9392 7463
rect 10882 7460 10910 7497
rect 22960 7485 22966 7497
rect 23018 7485 23024 7537
rect 36208 7485 36214 7537
rect 36266 7525 36272 7537
rect 39586 7525 39614 7562
rect 41008 7559 41014 7611
rect 41066 7599 41072 7611
rect 41107 7602 41165 7608
rect 41107 7599 41119 7602
rect 41066 7571 41119 7599
rect 41066 7559 41072 7571
rect 41107 7568 41119 7571
rect 41153 7568 41165 7602
rect 41107 7562 41165 7568
rect 45232 7559 45238 7611
rect 45290 7599 45296 7611
rect 45523 7602 45581 7608
rect 45523 7599 45535 7602
rect 45290 7571 45535 7599
rect 45290 7559 45296 7571
rect 45523 7568 45535 7571
rect 45569 7568 45581 7602
rect 45634 7599 45662 7645
rect 46192 7633 46198 7685
rect 46250 7673 46256 7685
rect 46291 7676 46349 7682
rect 46291 7673 46303 7676
rect 46250 7645 46303 7673
rect 46250 7633 46256 7645
rect 46291 7642 46303 7645
rect 46337 7642 46349 7676
rect 46291 7636 46349 7642
rect 47506 7645 48926 7673
rect 47506 7599 47534 7645
rect 45634 7571 47534 7599
rect 48898 7599 48926 7645
rect 48976 7633 48982 7685
rect 49034 7673 49040 7685
rect 49267 7676 49325 7682
rect 49267 7673 49279 7676
rect 49034 7645 49279 7673
rect 49034 7633 49040 7645
rect 49267 7642 49279 7645
rect 49313 7642 49325 7676
rect 49267 7636 49325 7642
rect 49648 7633 49654 7685
rect 49706 7673 49712 7685
rect 51091 7676 51149 7682
rect 51091 7673 51103 7676
rect 49706 7645 51103 7673
rect 49706 7633 49712 7645
rect 51091 7642 51103 7645
rect 51137 7642 51149 7676
rect 51091 7636 51149 7642
rect 52912 7633 52918 7685
rect 52970 7673 52976 7685
rect 55138 7682 55166 7719
rect 58768 7707 58774 7719
rect 58826 7707 58832 7759
rect 53299 7676 53357 7682
rect 53299 7673 53311 7676
rect 52970 7645 53311 7673
rect 52970 7633 52976 7645
rect 53299 7642 53311 7645
rect 53345 7642 53357 7676
rect 53299 7636 53357 7642
rect 55123 7676 55181 7682
rect 55123 7642 55135 7676
rect 55169 7642 55181 7676
rect 55792 7673 55798 7685
rect 55753 7645 55798 7673
rect 55123 7636 55181 7642
rect 55792 7633 55798 7645
rect 55850 7633 55856 7685
rect 56176 7633 56182 7685
rect 56234 7673 56240 7685
rect 56563 7676 56621 7682
rect 56563 7673 56575 7676
rect 56234 7645 56575 7673
rect 56234 7633 56240 7645
rect 56563 7642 56575 7645
rect 56609 7642 56621 7676
rect 56563 7636 56621 7642
rect 56656 7633 56662 7685
rect 56714 7673 56720 7685
rect 57331 7676 57389 7682
rect 57331 7673 57343 7676
rect 56714 7645 57343 7673
rect 56714 7633 56720 7645
rect 57331 7642 57343 7645
rect 57377 7642 57389 7676
rect 57331 7636 57389 7642
rect 49747 7602 49805 7608
rect 49747 7599 49759 7602
rect 48898 7571 49759 7599
rect 45523 7562 45581 7568
rect 49747 7568 49759 7571
rect 49793 7599 49805 7602
rect 50035 7602 50093 7608
rect 50035 7599 50047 7602
rect 49793 7571 50047 7599
rect 49793 7568 49805 7571
rect 49747 7562 49805 7568
rect 50035 7568 50047 7571
rect 50081 7568 50093 7602
rect 50035 7562 50093 7568
rect 36266 7497 39614 7525
rect 47506 7497 47966 7525
rect 36266 7485 36272 7497
rect 10867 7454 10925 7460
rect 10867 7420 10879 7454
rect 10913 7420 10925 7454
rect 10867 7414 10925 7420
rect 10960 7411 10966 7463
rect 11018 7451 11024 7463
rect 12307 7454 12365 7460
rect 12307 7451 12319 7454
rect 11018 7423 12319 7451
rect 11018 7411 11024 7423
rect 12307 7420 12319 7423
rect 12353 7420 12365 7454
rect 12307 7414 12365 7420
rect 12496 7411 12502 7463
rect 12554 7451 12560 7463
rect 13843 7454 13901 7460
rect 13843 7451 13855 7454
rect 12554 7423 13855 7451
rect 12554 7411 12560 7423
rect 13843 7420 13855 7423
rect 13889 7420 13901 7454
rect 13843 7414 13901 7420
rect 15664 7411 15670 7463
rect 15722 7451 15728 7463
rect 15763 7454 15821 7460
rect 15763 7451 15775 7454
rect 15722 7423 15775 7451
rect 15722 7411 15728 7423
rect 15763 7420 15775 7423
rect 15809 7420 15821 7454
rect 15763 7414 15821 7420
rect 15856 7411 15862 7463
rect 15914 7451 15920 7463
rect 16144 7451 16150 7463
rect 15914 7423 16150 7451
rect 15914 7411 15920 7423
rect 16144 7411 16150 7423
rect 16202 7411 16208 7463
rect 20752 7411 20758 7463
rect 20810 7451 20816 7463
rect 20851 7454 20909 7460
rect 20851 7451 20863 7454
rect 20810 7423 20863 7451
rect 20810 7411 20816 7423
rect 20851 7420 20863 7423
rect 20897 7420 20909 7454
rect 23824 7451 23830 7463
rect 23785 7423 23830 7451
rect 20851 7414 20909 7420
rect 23824 7411 23830 7423
rect 23882 7411 23888 7463
rect 24112 7411 24118 7463
rect 24170 7451 24176 7463
rect 24595 7454 24653 7460
rect 24595 7451 24607 7454
rect 24170 7423 24607 7451
rect 24170 7411 24176 7423
rect 24595 7420 24607 7423
rect 24641 7420 24653 7454
rect 24595 7414 24653 7420
rect 24784 7411 24790 7463
rect 24842 7451 24848 7463
rect 25363 7454 25421 7460
rect 25363 7451 25375 7454
rect 24842 7423 25375 7451
rect 24842 7411 24848 7423
rect 25363 7420 25375 7423
rect 25409 7420 25421 7454
rect 25363 7414 25421 7420
rect 25552 7411 25558 7463
rect 25610 7451 25616 7463
rect 26131 7454 26189 7460
rect 26131 7451 26143 7454
rect 25610 7423 26143 7451
rect 25610 7411 25616 7423
rect 26131 7420 26143 7423
rect 26177 7420 26189 7454
rect 26131 7414 26189 7420
rect 26704 7411 26710 7463
rect 26762 7451 26768 7463
rect 26899 7454 26957 7460
rect 26899 7451 26911 7454
rect 26762 7423 26911 7451
rect 26762 7411 26768 7423
rect 26899 7420 26911 7423
rect 26945 7420 26957 7454
rect 26899 7414 26957 7420
rect 28144 7411 28150 7463
rect 28202 7451 28208 7463
rect 28243 7454 28301 7460
rect 28243 7451 28255 7454
rect 28202 7423 28255 7451
rect 28202 7411 28208 7423
rect 28243 7420 28255 7423
rect 28289 7420 28301 7454
rect 28243 7414 28301 7420
rect 29200 7411 29206 7463
rect 29258 7451 29264 7463
rect 29299 7454 29357 7460
rect 29299 7451 29311 7454
rect 29258 7423 29311 7451
rect 29258 7411 29264 7423
rect 29299 7420 29311 7423
rect 29345 7420 29357 7454
rect 29299 7414 29357 7420
rect 31024 7411 31030 7463
rect 31082 7451 31088 7463
rect 31123 7454 31181 7460
rect 31123 7451 31135 7454
rect 31082 7423 31135 7451
rect 31082 7411 31088 7423
rect 31123 7420 31135 7423
rect 31169 7420 31181 7454
rect 31123 7414 31181 7420
rect 33616 7411 33622 7463
rect 33674 7451 33680 7463
rect 33715 7454 33773 7460
rect 33715 7451 33727 7454
rect 33674 7423 33727 7451
rect 33674 7411 33680 7423
rect 33715 7420 33727 7423
rect 33761 7420 33773 7454
rect 33715 7414 33773 7420
rect 34384 7411 34390 7463
rect 34442 7451 34448 7463
rect 34483 7454 34541 7460
rect 34483 7451 34495 7454
rect 34442 7423 34495 7451
rect 34442 7411 34448 7423
rect 34483 7420 34495 7423
rect 34529 7420 34541 7454
rect 34483 7414 34541 7420
rect 34768 7411 34774 7463
rect 34826 7451 34832 7463
rect 35251 7454 35309 7460
rect 35251 7451 35263 7454
rect 34826 7423 35263 7451
rect 34826 7411 34832 7423
rect 35251 7420 35263 7423
rect 35297 7420 35309 7454
rect 35251 7414 35309 7420
rect 35824 7411 35830 7463
rect 35882 7451 35888 7463
rect 36019 7454 36077 7460
rect 36019 7451 36031 7454
rect 35882 7423 36031 7451
rect 35882 7411 35888 7423
rect 36019 7420 36031 7423
rect 36065 7420 36077 7454
rect 36019 7414 36077 7420
rect 36688 7411 36694 7463
rect 36746 7451 36752 7463
rect 36883 7454 36941 7460
rect 36883 7451 36895 7454
rect 36746 7423 36895 7451
rect 36746 7411 36752 7423
rect 36883 7420 36895 7423
rect 36929 7420 36941 7454
rect 36883 7414 36941 7420
rect 38032 7411 38038 7463
rect 38090 7451 38096 7463
rect 38707 7454 38765 7460
rect 38707 7451 38719 7454
rect 38090 7423 38719 7451
rect 38090 7411 38096 7423
rect 38707 7420 38719 7423
rect 38753 7420 38765 7454
rect 38707 7414 38765 7420
rect 38800 7411 38806 7463
rect 38858 7451 38864 7463
rect 39475 7454 39533 7460
rect 39475 7451 39487 7454
rect 38858 7423 39487 7451
rect 38858 7411 38864 7423
rect 39475 7420 39487 7423
rect 39521 7420 39533 7454
rect 39475 7414 39533 7420
rect 39568 7411 39574 7463
rect 39626 7451 39632 7463
rect 40243 7454 40301 7460
rect 40243 7451 40255 7454
rect 39626 7423 40255 7451
rect 39626 7411 39632 7423
rect 40243 7420 40255 7423
rect 40289 7420 40301 7454
rect 40243 7414 40301 7420
rect 41392 7411 41398 7463
rect 41450 7451 41456 7463
rect 41779 7454 41837 7460
rect 41779 7451 41791 7454
rect 41450 7423 41791 7451
rect 41450 7411 41456 7423
rect 41779 7420 41791 7423
rect 41825 7420 41837 7454
rect 41779 7414 41837 7420
rect 42448 7411 42454 7463
rect 42506 7451 42512 7463
rect 42643 7454 42701 7460
rect 42643 7451 42655 7454
rect 42506 7423 42655 7451
rect 42506 7411 42512 7423
rect 42643 7420 42655 7423
rect 42689 7420 42701 7454
rect 42643 7414 42701 7420
rect 43888 7411 43894 7463
rect 43946 7451 43952 7463
rect 43987 7454 44045 7460
rect 43987 7451 43999 7454
rect 43946 7423 43999 7451
rect 43946 7411 43952 7423
rect 43987 7420 43999 7423
rect 44033 7420 44045 7454
rect 43987 7414 44045 7420
rect 44656 7411 44662 7463
rect 44714 7451 44720 7463
rect 44755 7454 44813 7460
rect 44755 7451 44767 7454
rect 44714 7423 44767 7451
rect 44714 7411 44720 7423
rect 44755 7420 44767 7423
rect 44801 7420 44813 7454
rect 44755 7414 44813 7420
rect 46480 7411 46486 7463
rect 46538 7451 46544 7463
rect 47059 7454 47117 7460
rect 47059 7451 47071 7454
rect 46538 7423 47071 7451
rect 46538 7411 46544 7423
rect 47059 7420 47071 7423
rect 47105 7420 47117 7454
rect 47059 7414 47117 7420
rect 47248 7411 47254 7463
rect 47306 7451 47312 7463
rect 47506 7451 47534 7497
rect 47938 7460 47966 7497
rect 49072 7485 49078 7537
rect 49130 7525 49136 7537
rect 49130 7497 50174 7525
rect 49130 7485 49136 7497
rect 50146 7460 50174 7497
rect 51010 7497 57614 7525
rect 51010 7460 51038 7497
rect 47306 7423 47534 7451
rect 47923 7454 47981 7460
rect 47306 7411 47312 7423
rect 47923 7420 47935 7454
rect 47969 7420 47981 7454
rect 47923 7414 47981 7420
rect 50131 7454 50189 7460
rect 50131 7420 50143 7454
rect 50177 7420 50189 7454
rect 50131 7414 50189 7420
rect 50995 7454 51053 7460
rect 50995 7420 51007 7454
rect 51041 7420 51053 7454
rect 50995 7414 51053 7420
rect 51664 7411 51670 7463
rect 51722 7451 51728 7463
rect 51859 7454 51917 7460
rect 51859 7451 51871 7454
rect 51722 7423 51871 7451
rect 51722 7411 51728 7423
rect 51859 7420 51871 7423
rect 51905 7420 51917 7454
rect 51859 7414 51917 7420
rect 52336 7411 52342 7463
rect 52394 7451 52400 7463
rect 52531 7454 52589 7460
rect 52531 7451 52543 7454
rect 52394 7423 52543 7451
rect 52394 7411 52400 7423
rect 52531 7420 52543 7423
rect 52577 7420 52589 7454
rect 57586 7451 57614 7497
rect 59344 7451 59350 7463
rect 57586 7423 59350 7451
rect 52531 7414 52589 7420
rect 59344 7411 59350 7423
rect 59402 7411 59408 7463
rect 1152 7352 58848 7374
rect 1152 7300 19654 7352
rect 19706 7300 19718 7352
rect 19770 7300 19782 7352
rect 19834 7300 19846 7352
rect 19898 7300 50374 7352
rect 50426 7300 50438 7352
rect 50490 7300 50502 7352
rect 50554 7300 50566 7352
rect 50618 7300 58848 7352
rect 1152 7278 58848 7300
rect 5584 7189 5590 7241
rect 5642 7229 5648 7241
rect 25840 7229 25846 7241
rect 5642 7201 25846 7229
rect 5642 7189 5648 7201
rect 25840 7189 25846 7201
rect 25898 7189 25904 7241
rect 6544 7155 6550 7167
rect 4546 7127 6550 7155
rect 4546 7090 4574 7127
rect 6544 7115 6550 7127
rect 6602 7115 6608 7167
rect 10291 7158 10349 7164
rect 10291 7124 10303 7158
rect 10337 7155 10349 7158
rect 10576 7155 10582 7167
rect 10337 7127 10582 7155
rect 10337 7124 10349 7127
rect 10291 7118 10349 7124
rect 10576 7115 10582 7127
rect 10634 7155 10640 7167
rect 12400 7155 12406 7167
rect 10634 7127 12406 7155
rect 10634 7115 10640 7127
rect 12400 7115 12406 7127
rect 12458 7115 12464 7167
rect 20656 7115 20662 7167
rect 20714 7155 20720 7167
rect 20755 7158 20813 7164
rect 20755 7155 20767 7158
rect 20714 7127 20767 7155
rect 20714 7115 20720 7127
rect 20755 7124 20767 7127
rect 20801 7155 20813 7158
rect 23920 7155 23926 7167
rect 20801 7127 21086 7155
rect 23881 7127 23926 7155
rect 20801 7124 20813 7127
rect 20755 7118 20813 7124
rect 4531 7084 4589 7090
rect 4531 7050 4543 7084
rect 4577 7050 4589 7084
rect 4531 7044 4589 7050
rect 5779 7084 5837 7090
rect 5779 7050 5791 7084
rect 5825 7081 5837 7084
rect 6064 7081 6070 7093
rect 5825 7053 6070 7081
rect 5825 7050 5837 7053
rect 5779 7044 5837 7050
rect 6064 7041 6070 7053
rect 6122 7041 6128 7093
rect 7120 7041 7126 7093
rect 7178 7081 7184 7093
rect 15856 7081 15862 7093
rect 7178 7053 10718 7081
rect 15817 7053 15862 7081
rect 7178 7041 7184 7053
rect 1648 7007 1654 7019
rect 1609 6979 1654 7007
rect 1648 6967 1654 6979
rect 1706 6967 1712 7019
rect 2512 7007 2518 7019
rect 2473 6979 2518 7007
rect 2512 6967 2518 6979
rect 2570 6967 2576 7019
rect 3664 6967 3670 7019
rect 3722 7007 3728 7019
rect 5011 7010 5069 7016
rect 3722 6979 4574 7007
rect 3722 6967 3728 6979
rect 4435 6936 4493 6942
rect 4435 6902 4447 6936
rect 4481 6902 4493 6936
rect 4546 6933 4574 6979
rect 5011 6976 5023 7010
rect 5057 7007 5069 7010
rect 5299 7010 5357 7016
rect 5299 7007 5311 7010
rect 5057 6979 5311 7007
rect 5057 6976 5069 6979
rect 5011 6970 5069 6976
rect 5299 6976 5311 6979
rect 5345 7007 5357 7010
rect 6352 7007 6358 7019
rect 5345 6979 6358 7007
rect 5345 6976 5357 6979
rect 5299 6970 5357 6976
rect 6352 6967 6358 6979
rect 6410 6967 6416 7019
rect 6451 7010 6509 7016
rect 6451 6976 6463 7010
rect 6497 7007 6509 7010
rect 6835 7010 6893 7016
rect 6835 7007 6847 7010
rect 6497 6979 6847 7007
rect 6497 6976 6509 6979
rect 6451 6970 6509 6976
rect 6835 6976 6847 6979
rect 6881 7007 6893 7010
rect 7024 7007 7030 7019
rect 6881 6979 7030 7007
rect 6881 6976 6893 6979
rect 6835 6970 6893 6976
rect 7024 6967 7030 6979
rect 7082 6967 7088 7019
rect 7600 7007 7606 7019
rect 7561 6979 7606 7007
rect 7600 6967 7606 6979
rect 7658 6967 7664 7019
rect 8083 7010 8141 7016
rect 8083 6976 8095 7010
rect 8129 7007 8141 7010
rect 8129 6979 8414 7007
rect 8129 6976 8141 6979
rect 8083 6970 8141 6976
rect 5203 6936 5261 6942
rect 5203 6933 5215 6936
rect 4546 6905 5215 6933
rect 4435 6896 4493 6902
rect 5203 6902 5215 6905
rect 5249 6902 5261 6936
rect 5203 6896 5261 6902
rect 4450 6859 4478 6896
rect 5872 6893 5878 6945
rect 5930 6933 5936 6945
rect 5971 6936 6029 6942
rect 5971 6933 5983 6936
rect 5930 6905 5983 6933
rect 5930 6893 5936 6905
rect 5971 6902 5983 6905
rect 6017 6902 6029 6936
rect 5971 6896 6029 6902
rect 6544 6893 6550 6945
rect 6602 6933 6608 6945
rect 6739 6936 6797 6942
rect 6739 6933 6751 6936
rect 6602 6905 6751 6933
rect 6602 6893 6608 6905
rect 6739 6902 6751 6905
rect 6785 6902 6797 6936
rect 6739 6896 6797 6902
rect 6928 6893 6934 6945
rect 6986 6933 6992 6945
rect 8386 6942 8414 6979
rect 8848 6967 8854 7019
rect 8906 7007 8912 7019
rect 10576 7007 10582 7019
rect 8906 6979 10046 7007
rect 10537 6979 10582 7007
rect 8906 6967 8912 6979
rect 7507 6936 7565 6942
rect 7507 6933 7519 6936
rect 6986 6905 7519 6933
rect 6986 6893 6992 6905
rect 7507 6902 7519 6905
rect 7553 6902 7565 6936
rect 7507 6896 7565 6902
rect 8275 6936 8333 6942
rect 8275 6902 8287 6936
rect 8321 6902 8333 6936
rect 8275 6896 8333 6902
rect 8371 6936 8429 6942
rect 8371 6902 8383 6936
rect 8417 6933 8429 6936
rect 9232 6933 9238 6945
rect 8417 6905 9238 6933
rect 8417 6902 8429 6905
rect 8371 6896 8429 6902
rect 4450 6831 5246 6859
rect 5218 6797 5246 6831
rect 7312 6819 7318 6871
rect 7370 6859 7376 6871
rect 8290 6859 8318 6896
rect 9232 6893 9238 6905
rect 9290 6893 9296 6945
rect 9715 6936 9773 6942
rect 9715 6902 9727 6936
rect 9761 6902 9773 6936
rect 9715 6896 9773 6902
rect 7370 6831 8318 6859
rect 7370 6819 7376 6831
rect 5200 6745 5206 6797
rect 5258 6745 5264 6797
rect 8080 6745 8086 6797
rect 8138 6785 8144 6797
rect 9730 6785 9758 6896
rect 9808 6893 9814 6945
rect 9866 6933 9872 6945
rect 10018 6933 10046 6979
rect 10576 6967 10582 6979
rect 10634 6967 10640 7019
rect 10483 6936 10541 6942
rect 10483 6933 10495 6936
rect 9866 6905 9911 6933
rect 10018 6905 10495 6933
rect 9866 6893 9872 6905
rect 10483 6902 10495 6905
rect 10529 6902 10541 6936
rect 10483 6896 10541 6902
rect 10690 6859 10718 7053
rect 15856 7041 15862 7053
rect 15914 7041 15920 7093
rect 17011 7084 17069 7090
rect 17011 7050 17023 7084
rect 17057 7081 17069 7084
rect 17296 7081 17302 7093
rect 17057 7053 17302 7081
rect 17057 7050 17069 7053
rect 17011 7044 17069 7050
rect 17296 7041 17302 7053
rect 17354 7081 17360 7093
rect 17779 7084 17837 7090
rect 17354 7053 17447 7081
rect 17354 7041 17360 7053
rect 17779 7050 17791 7084
rect 17825 7081 17837 7084
rect 18067 7084 18125 7090
rect 18067 7081 18079 7084
rect 17825 7053 18079 7081
rect 17825 7050 17837 7053
rect 17779 7044 17837 7050
rect 18067 7050 18079 7053
rect 18113 7081 18125 7084
rect 18256 7081 18262 7093
rect 18113 7053 18262 7081
rect 18113 7050 18125 7053
rect 18067 7044 18125 7050
rect 18256 7041 18262 7053
rect 18314 7041 18320 7093
rect 18835 7084 18893 7090
rect 18835 7050 18847 7084
rect 18881 7081 18893 7084
rect 18928 7081 18934 7093
rect 18881 7053 18934 7081
rect 18881 7050 18893 7053
rect 18835 7044 18893 7050
rect 18928 7041 18934 7053
rect 18986 7041 18992 7093
rect 20083 7084 20141 7090
rect 20083 7050 20095 7084
rect 20129 7081 20141 7084
rect 20368 7081 20374 7093
rect 20129 7053 20374 7081
rect 20129 7050 20141 7053
rect 20083 7044 20141 7050
rect 20368 7041 20374 7053
rect 20426 7041 20432 7093
rect 21058 7090 21086 7127
rect 23920 7115 23926 7127
rect 23978 7155 23984 7167
rect 26800 7155 26806 7167
rect 23978 7127 24254 7155
rect 26761 7127 26806 7155
rect 23978 7115 23984 7127
rect 21043 7084 21101 7090
rect 21043 7050 21055 7084
rect 21089 7050 21101 7084
rect 21043 7044 21101 7050
rect 21424 7041 21430 7093
rect 21482 7081 21488 7093
rect 21907 7084 21965 7090
rect 21907 7081 21919 7084
rect 21482 7053 21919 7081
rect 21482 7041 21488 7053
rect 21907 7050 21919 7053
rect 21953 7050 21965 7084
rect 21907 7044 21965 7050
rect 22387 7084 22445 7090
rect 22387 7050 22399 7084
rect 22433 7081 22445 7084
rect 22672 7081 22678 7093
rect 22433 7053 22678 7081
rect 22433 7050 22445 7053
rect 22387 7044 22445 7050
rect 22672 7041 22678 7053
rect 22730 7041 22736 7093
rect 24226 7090 24254 7127
rect 26800 7115 26806 7127
rect 26858 7155 26864 7167
rect 29104 7155 29110 7167
rect 26858 7127 27134 7155
rect 29065 7127 29110 7155
rect 26858 7115 26864 7127
rect 24211 7084 24269 7090
rect 24211 7050 24223 7084
rect 24257 7050 24269 7084
rect 24211 7044 24269 7050
rect 25651 7084 25709 7090
rect 25651 7050 25663 7084
rect 25697 7081 25709 7084
rect 25744 7081 25750 7093
rect 25697 7053 25750 7081
rect 25697 7050 25709 7053
rect 25651 7044 25709 7050
rect 25744 7041 25750 7053
rect 25802 7041 25808 7093
rect 26416 7081 26422 7093
rect 26377 7053 26422 7081
rect 26416 7041 26422 7053
rect 26474 7041 26480 7093
rect 27106 7090 27134 7127
rect 29104 7115 29110 7127
rect 29162 7155 29168 7167
rect 36592 7155 36598 7167
rect 29162 7127 29438 7155
rect 36553 7127 36598 7155
rect 29162 7115 29168 7127
rect 27091 7084 27149 7090
rect 27091 7050 27103 7084
rect 27137 7050 27149 7084
rect 27091 7044 27149 7050
rect 27667 7084 27725 7090
rect 27667 7050 27679 7084
rect 27713 7081 27725 7084
rect 27955 7084 28013 7090
rect 27955 7081 27967 7084
rect 27713 7053 27967 7081
rect 27713 7050 27725 7053
rect 27667 7044 27725 7050
rect 27955 7050 27967 7053
rect 28001 7081 28013 7084
rect 28336 7081 28342 7093
rect 28001 7053 28342 7081
rect 28001 7050 28013 7053
rect 27955 7044 28013 7050
rect 28336 7041 28342 7053
rect 28394 7041 28400 7093
rect 28720 7081 28726 7093
rect 28681 7053 28726 7081
rect 28720 7041 28726 7053
rect 28778 7041 28784 7093
rect 29410 7090 29438 7127
rect 36592 7115 36598 7127
rect 36650 7155 36656 7167
rect 36650 7127 36926 7155
rect 36650 7115 36656 7127
rect 29395 7084 29453 7090
rect 29395 7050 29407 7084
rect 29441 7050 29453 7084
rect 30928 7081 30934 7093
rect 30889 7053 30934 7081
rect 29395 7044 29453 7050
rect 30928 7041 30934 7053
rect 30986 7041 30992 7093
rect 31696 7081 31702 7093
rect 31657 7053 31702 7081
rect 31696 7041 31702 7053
rect 31754 7041 31760 7093
rect 32179 7084 32237 7090
rect 32179 7050 32191 7084
rect 32225 7081 32237 7084
rect 32368 7081 32374 7093
rect 32225 7053 32374 7081
rect 32225 7050 32237 7053
rect 32179 7044 32237 7050
rect 32368 7041 32374 7053
rect 32426 7041 32432 7093
rect 32947 7084 33005 7090
rect 32947 7050 32959 7084
rect 32993 7081 33005 7084
rect 33232 7081 33238 7093
rect 32993 7053 33238 7081
rect 32993 7050 33005 7053
rect 32947 7044 33005 7050
rect 33232 7041 33238 7053
rect 33290 7041 33296 7093
rect 33808 7041 33814 7093
rect 33866 7081 33872 7093
rect 34771 7084 34829 7090
rect 34771 7081 34783 7084
rect 33866 7053 34783 7081
rect 33866 7041 33872 7053
rect 34771 7050 34783 7053
rect 34817 7050 34829 7084
rect 34771 7044 34829 7050
rect 36016 7041 36022 7093
rect 36074 7081 36080 7093
rect 36898 7090 36926 7127
rect 37456 7115 37462 7167
rect 37514 7155 37520 7167
rect 39664 7155 39670 7167
rect 37514 7127 37790 7155
rect 39625 7127 39670 7155
rect 37514 7115 37520 7127
rect 37762 7090 37790 7127
rect 39664 7115 39670 7127
rect 39722 7155 39728 7167
rect 41104 7155 41110 7167
rect 39722 7127 39998 7155
rect 41065 7127 41110 7155
rect 39722 7115 39728 7127
rect 36211 7084 36269 7090
rect 36211 7081 36223 7084
rect 36074 7053 36223 7081
rect 36074 7041 36080 7053
rect 36211 7050 36223 7053
rect 36257 7050 36269 7084
rect 36211 7044 36269 7050
rect 36883 7084 36941 7090
rect 36883 7050 36895 7084
rect 36929 7050 36941 7084
rect 36883 7044 36941 7050
rect 37747 7084 37805 7090
rect 37747 7050 37759 7084
rect 37793 7050 37805 7084
rect 38512 7081 38518 7093
rect 38473 7053 38518 7081
rect 37747 7044 37805 7050
rect 38512 7041 38518 7053
rect 38570 7041 38576 7093
rect 39280 7081 39286 7093
rect 39241 7053 39286 7081
rect 39280 7041 39286 7053
rect 39338 7041 39344 7093
rect 39970 7090 39998 7127
rect 41104 7115 41110 7127
rect 41162 7155 41168 7167
rect 41162 7127 41438 7155
rect 41162 7115 41168 7127
rect 41410 7090 41438 7127
rect 41776 7115 41782 7167
rect 41834 7155 41840 7167
rect 41875 7158 41933 7164
rect 41875 7155 41887 7158
rect 41834 7127 41887 7155
rect 41834 7115 41840 7127
rect 41875 7124 41887 7127
rect 41921 7155 41933 7158
rect 43408 7155 43414 7167
rect 41921 7127 42206 7155
rect 43369 7127 43414 7155
rect 41921 7124 41933 7127
rect 41875 7118 41933 7124
rect 42178 7090 42206 7127
rect 43408 7115 43414 7127
rect 43466 7155 43472 7167
rect 45043 7158 45101 7164
rect 43466 7127 43838 7155
rect 43466 7115 43472 7127
rect 39955 7084 40013 7090
rect 39955 7050 39967 7084
rect 40001 7050 40013 7084
rect 39955 7044 40013 7050
rect 41395 7084 41453 7090
rect 41395 7050 41407 7084
rect 41441 7050 41453 7084
rect 41395 7044 41453 7050
rect 42163 7084 42221 7090
rect 42163 7050 42175 7084
rect 42209 7050 42221 7084
rect 42163 7044 42221 7050
rect 42739 7084 42797 7090
rect 42739 7050 42751 7084
rect 42785 7081 42797 7084
rect 42928 7081 42934 7093
rect 42785 7053 42934 7081
rect 42785 7050 42797 7053
rect 42739 7044 42797 7050
rect 42928 7041 42934 7053
rect 42986 7041 42992 7093
rect 43810 7090 43838 7127
rect 45043 7124 45055 7158
rect 45089 7155 45101 7158
rect 45136 7155 45142 7167
rect 45089 7127 45142 7155
rect 45089 7124 45101 7127
rect 45043 7118 45101 7124
rect 45136 7115 45142 7127
rect 45194 7155 45200 7167
rect 48787 7158 48845 7164
rect 45194 7127 45278 7155
rect 45194 7115 45200 7127
rect 45250 7090 45278 7127
rect 48787 7124 48799 7158
rect 48833 7155 48845 7158
rect 48880 7155 48886 7167
rect 48833 7127 48886 7155
rect 48833 7124 48845 7127
rect 48787 7118 48845 7124
rect 48880 7115 48886 7127
rect 48938 7155 48944 7167
rect 48938 7127 49022 7155
rect 48938 7115 48944 7127
rect 43795 7084 43853 7090
rect 43795 7050 43807 7084
rect 43841 7050 43853 7084
rect 43795 7044 43853 7050
rect 45235 7084 45293 7090
rect 45235 7050 45247 7084
rect 45281 7050 45293 7084
rect 45235 7044 45293 7050
rect 46483 7084 46541 7090
rect 46483 7050 46495 7084
rect 46529 7081 46541 7084
rect 46672 7081 46678 7093
rect 46529 7053 46678 7081
rect 46529 7050 46541 7053
rect 46483 7044 46541 7050
rect 46672 7041 46678 7053
rect 46730 7041 46736 7093
rect 47539 7084 47597 7090
rect 47539 7050 47551 7084
rect 47585 7081 47597 7084
rect 47632 7081 47638 7093
rect 47585 7053 47638 7081
rect 47585 7050 47597 7053
rect 47539 7044 47597 7050
rect 47632 7041 47638 7053
rect 47690 7041 47696 7093
rect 48304 7081 48310 7093
rect 48265 7053 48310 7081
rect 48304 7041 48310 7053
rect 48362 7041 48368 7093
rect 48994 7090 49022 7127
rect 49840 7115 49846 7167
rect 49898 7155 49904 7167
rect 52435 7158 52493 7164
rect 52435 7155 52447 7158
rect 49898 7127 52447 7155
rect 49898 7115 49904 7127
rect 52435 7124 52447 7127
rect 52481 7155 52493 7158
rect 52481 7127 52766 7155
rect 52481 7124 52493 7127
rect 52435 7118 52493 7124
rect 48979 7084 49037 7090
rect 48979 7050 48991 7084
rect 49025 7050 49037 7084
rect 48979 7044 49037 7050
rect 50035 7084 50093 7090
rect 50035 7050 50047 7084
rect 50081 7081 50093 7084
rect 50224 7081 50230 7093
rect 50081 7053 50230 7081
rect 50081 7050 50093 7053
rect 50035 7044 50093 7050
rect 50224 7041 50230 7053
rect 50282 7041 50288 7093
rect 52048 7081 52054 7093
rect 52009 7053 52054 7081
rect 52048 7041 52054 7053
rect 52106 7041 52112 7093
rect 52738 7090 52766 7127
rect 52723 7084 52781 7090
rect 52723 7050 52735 7084
rect 52769 7050 52781 7084
rect 52723 7044 52781 7050
rect 11248 7007 11254 7019
rect 11209 6979 11254 7007
rect 11248 6967 11254 6979
rect 11306 6967 11312 7019
rect 12688 7007 12694 7019
rect 12649 6979 12694 7007
rect 12688 6967 12694 6979
rect 12746 6967 12752 7019
rect 15091 7010 15149 7016
rect 15091 6976 15103 7010
rect 15137 7007 15149 7010
rect 23443 7010 23501 7016
rect 15137 6979 22718 7007
rect 15137 6976 15149 6979
rect 15091 6970 15149 6976
rect 12304 6893 12310 6945
rect 12362 6933 12368 6945
rect 12880 6933 12886 6945
rect 12362 6905 12886 6933
rect 12362 6893 12368 6905
rect 12880 6893 12886 6905
rect 12938 6893 12944 6945
rect 13456 6893 13462 6945
rect 13514 6933 13520 6945
rect 13555 6936 13613 6942
rect 13555 6933 13567 6936
rect 13514 6905 13567 6933
rect 13514 6893 13520 6905
rect 13555 6902 13567 6905
rect 13601 6902 13613 6936
rect 13555 6896 13613 6902
rect 13651 6936 13709 6942
rect 13651 6902 13663 6936
rect 13697 6933 13709 6936
rect 13744 6933 13750 6945
rect 13697 6905 13750 6933
rect 13697 6902 13709 6905
rect 13651 6896 13709 6902
rect 13744 6893 13750 6905
rect 13802 6893 13808 6945
rect 14608 6893 14614 6945
rect 14666 6933 14672 6945
rect 14995 6936 15053 6942
rect 14995 6933 15007 6936
rect 14666 6905 15007 6933
rect 14666 6893 14672 6905
rect 14995 6902 15007 6905
rect 15041 6902 15053 6936
rect 14995 6896 15053 6902
rect 15376 6893 15382 6945
rect 15434 6933 15440 6945
rect 15763 6936 15821 6942
rect 15763 6933 15775 6936
rect 15434 6905 15775 6933
rect 15434 6893 15440 6905
rect 15763 6902 15775 6905
rect 15809 6902 15821 6936
rect 15763 6896 15821 6902
rect 17104 6893 17110 6945
rect 17162 6933 17168 6945
rect 17203 6936 17261 6942
rect 17203 6933 17215 6936
rect 17162 6905 17215 6933
rect 17162 6893 17168 6905
rect 17203 6902 17215 6905
rect 17249 6902 17261 6936
rect 17203 6896 17261 6902
rect 17872 6893 17878 6945
rect 17930 6933 17936 6945
rect 17971 6936 18029 6942
rect 17971 6933 17983 6936
rect 17930 6905 17983 6933
rect 17930 6893 17936 6905
rect 17971 6902 17983 6905
rect 18017 6902 18029 6936
rect 17971 6896 18029 6902
rect 18544 6893 18550 6945
rect 18602 6933 18608 6945
rect 18739 6936 18797 6942
rect 18739 6933 18751 6936
rect 18602 6905 18751 6933
rect 18602 6893 18608 6905
rect 18739 6902 18751 6905
rect 18785 6902 18797 6936
rect 18739 6896 18797 6902
rect 20275 6936 20333 6942
rect 20275 6902 20287 6936
rect 20321 6933 20333 6936
rect 20368 6933 20374 6945
rect 20321 6905 20374 6933
rect 20321 6902 20333 6905
rect 20275 6896 20333 6902
rect 20368 6893 20374 6905
rect 20426 6893 20432 6945
rect 20944 6893 20950 6945
rect 21002 6933 21008 6945
rect 21139 6936 21197 6942
rect 21139 6933 21151 6936
rect 21002 6905 21151 6933
rect 21002 6893 21008 6905
rect 21139 6902 21151 6905
rect 21185 6902 21197 6936
rect 21139 6896 21197 6902
rect 21232 6893 21238 6945
rect 21290 6933 21296 6945
rect 21811 6936 21869 6942
rect 21811 6933 21823 6936
rect 21290 6905 21823 6933
rect 21290 6893 21296 6905
rect 21811 6902 21823 6905
rect 21857 6902 21869 6936
rect 21811 6896 21869 6902
rect 22000 6893 22006 6945
rect 22058 6933 22064 6945
rect 22579 6936 22637 6942
rect 22579 6933 22591 6936
rect 22058 6905 22591 6933
rect 22058 6893 22064 6905
rect 22579 6902 22591 6905
rect 22625 6902 22637 6936
rect 22579 6896 22637 6902
rect 10690 6831 15854 6859
rect 8138 6757 9758 6785
rect 15826 6785 15854 6831
rect 16240 6785 16246 6797
rect 15826 6757 16246 6785
rect 8138 6745 8144 6757
rect 16240 6745 16246 6757
rect 16298 6745 16304 6797
rect 22690 6785 22718 6979
rect 23443 6976 23455 7010
rect 23489 7007 23501 7010
rect 25168 7007 25174 7019
rect 23489 6979 25174 7007
rect 23489 6976 23501 6979
rect 23443 6970 23501 6976
rect 25168 6967 25174 6979
rect 25226 6967 25232 7019
rect 25936 6967 25942 7019
rect 25994 7007 26000 7019
rect 25994 6979 27230 7007
rect 25994 6967 26000 6979
rect 23344 6933 23350 6945
rect 23305 6905 23350 6933
rect 23344 6893 23350 6905
rect 23402 6893 23408 6945
rect 23920 6893 23926 6945
rect 23978 6933 23984 6945
rect 24115 6936 24173 6942
rect 24115 6933 24127 6936
rect 23978 6905 24127 6933
rect 23978 6893 23984 6905
rect 24115 6902 24127 6905
rect 24161 6902 24173 6936
rect 24115 6896 24173 6902
rect 24592 6893 24598 6945
rect 24650 6933 24656 6945
rect 27202 6942 27230 6979
rect 31408 6967 31414 7019
rect 31466 7007 31472 7019
rect 31466 6979 32510 7007
rect 31466 6967 31472 6979
rect 25555 6936 25613 6942
rect 25555 6933 25567 6936
rect 24650 6905 25567 6933
rect 24650 6893 24656 6905
rect 25555 6902 25567 6905
rect 25601 6902 25613 6936
rect 25555 6896 25613 6902
rect 26323 6936 26381 6942
rect 26323 6902 26335 6936
rect 26369 6902 26381 6936
rect 26323 6896 26381 6902
rect 27187 6936 27245 6942
rect 27187 6902 27199 6936
rect 27233 6902 27245 6936
rect 27859 6936 27917 6942
rect 27859 6933 27871 6936
rect 27187 6896 27245 6902
rect 27346 6905 27871 6933
rect 25168 6819 25174 6871
rect 25226 6859 25232 6871
rect 26338 6859 26366 6896
rect 25226 6831 26366 6859
rect 25226 6819 25232 6831
rect 26992 6819 26998 6871
rect 27050 6859 27056 6871
rect 27346 6859 27374 6905
rect 27859 6902 27871 6905
rect 27905 6902 27917 6936
rect 27859 6896 27917 6902
rect 28627 6936 28685 6942
rect 28627 6902 28639 6936
rect 28673 6902 28685 6936
rect 29488 6933 29494 6945
rect 29449 6905 29494 6933
rect 28627 6896 28685 6902
rect 27050 6831 27374 6859
rect 27050 6819 27056 6831
rect 27760 6819 27766 6871
rect 27818 6859 27824 6871
rect 28642 6859 28670 6896
rect 29488 6893 29494 6905
rect 29546 6893 29552 6945
rect 29968 6893 29974 6945
rect 30026 6933 30032 6945
rect 32482 6942 32510 6979
rect 32560 6967 32566 7019
rect 32618 7007 32624 7019
rect 34003 7010 34061 7016
rect 34003 7007 34015 7010
rect 32618 6979 34015 7007
rect 32618 6967 32624 6979
rect 34003 6976 34015 6979
rect 34049 6976 34061 7010
rect 34003 6970 34061 6976
rect 38530 6979 40094 7007
rect 38530 6945 38558 6979
rect 30835 6936 30893 6942
rect 30835 6933 30847 6936
rect 30026 6905 30847 6933
rect 30026 6893 30032 6905
rect 30835 6902 30847 6905
rect 30881 6902 30893 6936
rect 30835 6896 30893 6902
rect 31603 6936 31661 6942
rect 31603 6902 31615 6936
rect 31649 6902 31661 6936
rect 31603 6896 31661 6902
rect 32467 6936 32525 6942
rect 32467 6902 32479 6936
rect 32513 6902 32525 6936
rect 32467 6896 32525 6902
rect 33139 6936 33197 6942
rect 33139 6902 33151 6936
rect 33185 6902 33197 6936
rect 33139 6896 33197 6902
rect 33907 6936 33965 6942
rect 33907 6902 33919 6936
rect 33953 6902 33965 6936
rect 34675 6936 34733 6942
rect 34675 6933 34687 6936
rect 33907 6896 33965 6902
rect 34018 6905 34687 6933
rect 27818 6831 28670 6859
rect 27818 6819 27824 6831
rect 30736 6819 30742 6871
rect 30794 6859 30800 6871
rect 31618 6859 31646 6896
rect 30794 6831 31646 6859
rect 30794 6819 30800 6831
rect 32176 6819 32182 6871
rect 32234 6859 32240 6871
rect 33154 6859 33182 6896
rect 32234 6831 33182 6859
rect 32234 6819 32240 6831
rect 26608 6785 26614 6797
rect 22690 6757 26614 6785
rect 26608 6745 26614 6757
rect 26666 6745 26672 6797
rect 32944 6745 32950 6797
rect 33002 6785 33008 6797
rect 33922 6785 33950 6896
rect 34018 6871 34046 6905
rect 34675 6902 34687 6905
rect 34721 6902 34733 6936
rect 34675 6896 34733 6902
rect 35536 6893 35542 6945
rect 35594 6933 35600 6945
rect 36115 6936 36173 6942
rect 36115 6933 36127 6936
rect 35594 6905 36127 6933
rect 35594 6893 35600 6905
rect 36115 6902 36127 6905
rect 36161 6902 36173 6936
rect 36115 6896 36173 6902
rect 36400 6893 36406 6945
rect 36458 6933 36464 6945
rect 36979 6936 37037 6942
rect 36979 6933 36991 6936
rect 36458 6905 36991 6933
rect 36458 6893 36464 6905
rect 36979 6902 36991 6905
rect 37025 6902 37037 6936
rect 36979 6896 37037 6902
rect 37072 6893 37078 6945
rect 37130 6933 37136 6945
rect 37651 6936 37709 6942
rect 37651 6933 37663 6936
rect 37130 6905 37663 6933
rect 37130 6893 37136 6905
rect 37651 6902 37663 6905
rect 37697 6902 37709 6936
rect 37651 6896 37709 6902
rect 38419 6936 38477 6942
rect 38419 6902 38431 6936
rect 38465 6902 38477 6936
rect 38419 6896 38477 6902
rect 34000 6819 34006 6871
rect 34058 6819 34064 6871
rect 37360 6819 37366 6871
rect 37418 6859 37424 6871
rect 38434 6859 38462 6896
rect 38512 6893 38518 6945
rect 38570 6893 38576 6945
rect 40066 6942 40094 6979
rect 41200 6967 41206 7019
rect 41258 7007 41264 7019
rect 44275 7010 44333 7016
rect 41258 6979 43070 7007
rect 41258 6967 41264 6979
rect 43042 6942 43070 6979
rect 44275 6976 44287 7010
rect 44321 7007 44333 7010
rect 44563 7010 44621 7016
rect 44563 7007 44575 7010
rect 44321 6979 44575 7007
rect 44321 6976 44333 6979
rect 44275 6970 44333 6976
rect 44563 6976 44575 6979
rect 44609 7007 44621 7010
rect 47824 7007 47830 7019
rect 44609 6979 47830 7007
rect 44609 6976 44621 6979
rect 44563 6970 44621 6976
rect 47824 6967 47830 6979
rect 47882 6967 47888 7019
rect 54067 7010 54125 7016
rect 54067 6976 54079 7010
rect 54113 6976 54125 7010
rect 54736 7007 54742 7019
rect 54697 6979 54742 7007
rect 54067 6970 54125 6976
rect 39187 6936 39245 6942
rect 39187 6902 39199 6936
rect 39233 6902 39245 6936
rect 39187 6896 39245 6902
rect 40051 6936 40109 6942
rect 40051 6902 40063 6936
rect 40097 6902 40109 6936
rect 41491 6936 41549 6942
rect 41491 6933 41503 6936
rect 40051 6896 40109 6902
rect 40162 6905 41503 6933
rect 37418 6831 38462 6859
rect 37418 6819 37424 6831
rect 33002 6757 33950 6785
rect 33002 6745 33008 6757
rect 37648 6745 37654 6797
rect 37706 6785 37712 6797
rect 39202 6785 39230 6896
rect 39856 6819 39862 6871
rect 39914 6859 39920 6871
rect 40162 6859 40190 6905
rect 41491 6902 41503 6905
rect 41537 6902 41549 6936
rect 41491 6896 41549 6902
rect 42259 6936 42317 6942
rect 42259 6902 42271 6936
rect 42305 6902 42317 6936
rect 42259 6896 42317 6902
rect 43027 6936 43085 6942
rect 43027 6902 43039 6936
rect 43073 6902 43085 6936
rect 43027 6896 43085 6902
rect 43699 6936 43757 6942
rect 43699 6902 43711 6936
rect 43745 6902 43757 6936
rect 43699 6896 43757 6902
rect 44467 6936 44525 6942
rect 44467 6902 44479 6936
rect 44513 6902 44525 6936
rect 44467 6896 44525 6902
rect 45331 6936 45389 6942
rect 45331 6902 45343 6936
rect 45377 6902 45389 6936
rect 45331 6896 45389 6902
rect 39914 6831 40190 6859
rect 39914 6819 39920 6831
rect 41296 6819 41302 6871
rect 41354 6859 41360 6871
rect 42274 6859 42302 6896
rect 41354 6831 42302 6859
rect 41354 6819 41360 6831
rect 42832 6819 42838 6871
rect 42890 6859 42896 6871
rect 43714 6859 43742 6896
rect 42890 6831 43742 6859
rect 42890 6819 42896 6831
rect 37706 6757 39230 6785
rect 37706 6745 37712 6757
rect 43600 6745 43606 6797
rect 43658 6785 43664 6797
rect 44482 6785 44510 6896
rect 44560 6819 44566 6871
rect 44618 6859 44624 6871
rect 45346 6859 45374 6896
rect 45424 6893 45430 6945
rect 45482 6933 45488 6945
rect 46771 6936 46829 6942
rect 46771 6933 46783 6936
rect 45482 6905 46783 6933
rect 45482 6893 45488 6905
rect 46771 6902 46783 6905
rect 46817 6902 46829 6936
rect 46771 6896 46829 6902
rect 47056 6893 47062 6945
rect 47114 6933 47120 6945
rect 47443 6936 47501 6942
rect 47443 6933 47455 6936
rect 47114 6905 47455 6933
rect 47114 6893 47120 6905
rect 47443 6902 47455 6905
rect 47489 6902 47501 6936
rect 47443 6896 47501 6902
rect 48211 6936 48269 6942
rect 48211 6902 48223 6936
rect 48257 6902 48269 6936
rect 48211 6896 48269 6902
rect 44618 6831 45374 6859
rect 44618 6819 44624 6831
rect 46864 6819 46870 6871
rect 46922 6859 46928 6871
rect 48226 6859 48254 6896
rect 48880 6893 48886 6945
rect 48938 6933 48944 6945
rect 49075 6936 49133 6942
rect 49075 6933 49087 6936
rect 48938 6905 49087 6933
rect 48938 6893 48944 6905
rect 49075 6902 49087 6905
rect 49121 6902 49133 6936
rect 49075 6896 49133 6902
rect 50128 6893 50134 6945
rect 50186 6933 50192 6945
rect 50323 6936 50381 6942
rect 50323 6933 50335 6936
rect 50186 6905 50335 6933
rect 50186 6893 50192 6905
rect 50323 6902 50335 6905
rect 50369 6902 50381 6936
rect 50323 6896 50381 6902
rect 51376 6893 51382 6945
rect 51434 6933 51440 6945
rect 51955 6936 52013 6942
rect 51955 6933 51967 6936
rect 51434 6905 51967 6933
rect 51434 6893 51440 6905
rect 51955 6902 51967 6905
rect 52001 6902 52013 6936
rect 52816 6933 52822 6945
rect 52777 6905 52822 6933
rect 51955 6896 52013 6902
rect 52816 6893 52822 6905
rect 52874 6893 52880 6945
rect 54082 6933 54110 6970
rect 54736 6967 54742 6979
rect 54794 6967 54800 7019
rect 55408 6967 55414 7019
rect 55466 7007 55472 7019
rect 55507 7010 55565 7016
rect 55507 7007 55519 7010
rect 55466 6979 55519 7007
rect 55466 6967 55472 6979
rect 55507 6976 55519 6979
rect 55553 6976 55565 7010
rect 55507 6970 55565 6976
rect 57811 7010 57869 7016
rect 57811 6976 57823 7010
rect 57857 7007 57869 7010
rect 58480 7007 58486 7019
rect 57857 6979 58486 7007
rect 57857 6976 57869 6979
rect 57811 6970 57869 6976
rect 58480 6967 58486 6979
rect 58538 6967 58544 7019
rect 56368 6933 56374 6945
rect 54082 6905 56374 6933
rect 56368 6893 56374 6905
rect 56426 6893 56432 6945
rect 46922 6831 48254 6859
rect 46922 6819 46928 6831
rect 43658 6757 44510 6785
rect 43658 6745 43664 6757
rect 1152 6686 58848 6708
rect 1152 6634 4294 6686
rect 4346 6634 4358 6686
rect 4410 6634 4422 6686
rect 4474 6634 4486 6686
rect 4538 6634 35014 6686
rect 35066 6634 35078 6686
rect 35130 6634 35142 6686
rect 35194 6634 35206 6686
rect 35258 6634 58848 6686
rect 1152 6612 58848 6634
rect 5392 6563 5398 6575
rect 5353 6535 5398 6563
rect 5392 6523 5398 6535
rect 5450 6563 5456 6575
rect 5450 6535 5726 6563
rect 5450 6523 5456 6535
rect 5698 6424 5726 6535
rect 7906 6535 8270 6563
rect 7603 6492 7661 6498
rect 7603 6458 7615 6492
rect 7649 6489 7661 6492
rect 7906 6489 7934 6535
rect 7649 6461 7934 6489
rect 8242 6489 8270 6535
rect 8464 6523 8470 6575
rect 8522 6563 8528 6575
rect 9328 6563 9334 6575
rect 8522 6535 9334 6563
rect 8522 6523 8528 6535
rect 9328 6523 9334 6535
rect 9386 6523 9392 6575
rect 15952 6563 15958 6575
rect 15913 6535 15958 6563
rect 15952 6523 15958 6535
rect 16010 6563 16016 6575
rect 30256 6563 30262 6575
rect 16010 6535 16286 6563
rect 30217 6535 30262 6563
rect 16010 6523 16016 6535
rect 9040 6489 9046 6501
rect 8242 6461 9046 6489
rect 7649 6458 7661 6461
rect 7603 6452 7661 6458
rect 9040 6449 9046 6461
rect 9098 6449 9104 6501
rect 13651 6492 13709 6498
rect 13651 6458 13663 6492
rect 13697 6489 13709 6492
rect 13697 6461 13982 6489
rect 13697 6458 13709 6461
rect 13651 6452 13709 6458
rect 13954 6427 13982 6461
rect 5683 6418 5741 6424
rect 5683 6384 5695 6418
rect 5729 6384 5741 6418
rect 7120 6415 7126 6427
rect 7081 6387 7126 6415
rect 5683 6378 5741 6384
rect 7120 6375 7126 6387
rect 7178 6375 7184 6427
rect 7216 6375 7222 6427
rect 7274 6415 7280 6427
rect 8368 6415 8374 6427
rect 7274 6387 7968 6415
rect 8256 6387 8374 6415
rect 7274 6375 7280 6387
rect 8368 6375 8374 6387
rect 8426 6375 8432 6427
rect 13072 6375 13078 6427
rect 13130 6415 13136 6427
rect 13843 6418 13901 6424
rect 13843 6415 13855 6418
rect 13130 6387 13855 6415
rect 13130 6375 13136 6387
rect 13843 6384 13855 6387
rect 13889 6384 13901 6418
rect 13843 6378 13901 6384
rect 13936 6375 13942 6427
rect 13994 6415 14000 6427
rect 15472 6415 15478 6427
rect 13994 6387 14039 6415
rect 15433 6387 15478 6415
rect 13994 6375 14000 6387
rect 15472 6375 15478 6387
rect 15530 6375 15536 6427
rect 16258 6424 16286 6535
rect 30256 6523 30262 6535
rect 30314 6563 30320 6575
rect 31792 6563 31798 6575
rect 30314 6535 30590 6563
rect 31753 6535 31798 6563
rect 30314 6523 30320 6535
rect 16243 6418 16301 6424
rect 16243 6384 16255 6418
rect 16289 6384 16301 6418
rect 16243 6378 16301 6384
rect 17395 6418 17453 6424
rect 17395 6384 17407 6418
rect 17441 6415 17453 6418
rect 17680 6415 17686 6427
rect 17441 6387 17686 6415
rect 17441 6384 17453 6387
rect 17395 6378 17453 6384
rect 17680 6375 17686 6387
rect 17738 6375 17744 6427
rect 18448 6415 18454 6427
rect 18409 6387 18454 6415
rect 18448 6375 18454 6387
rect 18506 6375 18512 6427
rect 18931 6418 18989 6424
rect 18931 6384 18943 6418
rect 18977 6415 18989 6418
rect 19120 6415 19126 6427
rect 18977 6387 19126 6415
rect 18977 6384 18989 6387
rect 18931 6378 18989 6384
rect 19120 6375 19126 6387
rect 19178 6375 19184 6427
rect 19699 6418 19757 6424
rect 19699 6384 19711 6418
rect 19745 6415 19757 6418
rect 19984 6415 19990 6427
rect 19745 6387 19990 6415
rect 19745 6384 19757 6387
rect 19699 6378 19757 6384
rect 19984 6375 19990 6387
rect 20042 6375 20048 6427
rect 20755 6418 20813 6424
rect 20755 6384 20767 6418
rect 20801 6415 20813 6418
rect 20848 6415 20854 6427
rect 20801 6387 20854 6415
rect 20801 6384 20813 6387
rect 20755 6378 20813 6384
rect 20848 6375 20854 6387
rect 20906 6375 20912 6427
rect 21520 6415 21526 6427
rect 21481 6387 21526 6415
rect 21520 6375 21526 6387
rect 21578 6375 21584 6427
rect 23728 6415 23734 6427
rect 23689 6387 23734 6415
rect 23728 6375 23734 6387
rect 23786 6375 23792 6427
rect 24211 6418 24269 6424
rect 24211 6384 24223 6418
rect 24257 6415 24269 6418
rect 24496 6415 24502 6427
rect 24257 6387 24502 6415
rect 24257 6384 24269 6387
rect 24211 6378 24269 6384
rect 24496 6375 24502 6387
rect 24554 6375 24560 6427
rect 28240 6415 28246 6427
rect 28201 6387 28246 6415
rect 28240 6375 28246 6387
rect 28298 6375 28304 6427
rect 29008 6415 29014 6427
rect 28969 6387 29014 6415
rect 29008 6375 29014 6387
rect 29066 6375 29072 6427
rect 30562 6424 30590 6535
rect 31792 6523 31798 6535
rect 31850 6563 31856 6575
rect 34771 6566 34829 6572
rect 31850 6535 32222 6563
rect 31850 6523 31856 6535
rect 30547 6418 30605 6424
rect 30547 6384 30559 6418
rect 30593 6384 30605 6418
rect 30547 6378 30605 6384
rect 30640 6375 30646 6427
rect 30698 6415 30704 6427
rect 32194 6424 32222 6535
rect 34771 6532 34783 6566
rect 34817 6563 34829 6566
rect 34864 6563 34870 6575
rect 34817 6535 34870 6563
rect 34817 6532 34829 6535
rect 34771 6526 34829 6532
rect 34864 6523 34870 6535
rect 34922 6563 34928 6575
rect 36880 6563 36886 6575
rect 34922 6535 35006 6563
rect 36841 6535 36886 6563
rect 34922 6523 34928 6535
rect 32083 6418 32141 6424
rect 32083 6415 32095 6418
rect 30698 6387 32095 6415
rect 30698 6375 30704 6387
rect 32083 6384 32095 6387
rect 32129 6384 32141 6418
rect 32083 6378 32141 6384
rect 32179 6418 32237 6424
rect 32179 6384 32191 6418
rect 32225 6384 32237 6418
rect 33520 6415 33526 6427
rect 33481 6387 33526 6415
rect 32179 6378 32237 6384
rect 33520 6375 33526 6387
rect 33578 6375 33584 6427
rect 34003 6418 34061 6424
rect 34003 6384 34015 6418
rect 34049 6415 34061 6418
rect 34192 6415 34198 6427
rect 34049 6387 34198 6415
rect 34049 6384 34061 6387
rect 34003 6378 34061 6384
rect 34192 6375 34198 6387
rect 34250 6375 34256 6427
rect 34978 6424 35006 6535
rect 36880 6523 36886 6535
rect 36938 6563 36944 6575
rect 51280 6563 51286 6575
rect 36938 6535 37310 6563
rect 51241 6535 51286 6563
rect 36938 6523 36944 6535
rect 37282 6424 37310 6535
rect 51280 6523 51286 6535
rect 51338 6563 51344 6575
rect 51338 6535 51614 6563
rect 51338 6523 51344 6535
rect 39859 6492 39917 6498
rect 39859 6458 39871 6492
rect 39905 6489 39917 6492
rect 47728 6489 47734 6501
rect 39905 6461 47734 6489
rect 39905 6458 39917 6461
rect 39859 6452 39917 6458
rect 47728 6449 47734 6461
rect 47786 6449 47792 6501
rect 34963 6418 35021 6424
rect 34963 6384 34975 6418
rect 35009 6384 35021 6418
rect 34963 6378 35021 6384
rect 37267 6418 37325 6424
rect 37267 6384 37279 6418
rect 37313 6384 37325 6418
rect 37267 6378 37325 6384
rect 42547 6418 42605 6424
rect 42547 6384 42559 6418
rect 42593 6415 42605 6418
rect 42736 6415 42742 6427
rect 42593 6387 42742 6415
rect 42593 6384 42605 6387
rect 42547 6378 42605 6384
rect 42736 6375 42742 6387
rect 42794 6375 42800 6427
rect 44752 6375 44758 6427
rect 44810 6415 44816 6427
rect 44851 6418 44909 6424
rect 44851 6415 44863 6418
rect 44810 6387 44863 6415
rect 44810 6375 44816 6387
rect 44851 6384 44863 6387
rect 44897 6384 44909 6418
rect 50896 6415 50902 6427
rect 50857 6387 50902 6415
rect 44851 6378 44909 6384
rect 50896 6375 50902 6387
rect 50954 6375 50960 6427
rect 51586 6424 51614 6535
rect 51571 6418 51629 6424
rect 51571 6384 51583 6418
rect 51617 6384 51629 6418
rect 52432 6415 52438 6427
rect 52393 6387 52438 6415
rect 51571 6378 51629 6384
rect 52432 6375 52438 6387
rect 52490 6375 52496 6427
rect 56848 6415 56854 6427
rect 53314 6387 56854 6415
rect 1552 6341 1558 6353
rect 1513 6313 1558 6341
rect 1552 6301 1558 6313
rect 1610 6301 1616 6353
rect 2032 6301 2038 6353
rect 2090 6341 2096 6353
rect 2323 6344 2381 6350
rect 2323 6341 2335 6344
rect 2090 6313 2335 6341
rect 2090 6301 2096 6313
rect 2323 6310 2335 6313
rect 2369 6310 2381 6344
rect 3184 6341 3190 6353
rect 3145 6313 3190 6341
rect 2323 6304 2381 6310
rect 3184 6301 3190 6313
rect 3242 6301 3248 6353
rect 3856 6301 3862 6353
rect 3914 6341 3920 6353
rect 3955 6344 4013 6350
rect 3955 6341 3967 6344
rect 3914 6313 3967 6341
rect 3914 6301 3920 6313
rect 3955 6310 3967 6313
rect 4001 6310 4013 6344
rect 3955 6304 4013 6310
rect 4624 6301 4630 6353
rect 4682 6341 4688 6353
rect 4723 6344 4781 6350
rect 4723 6341 4735 6344
rect 4682 6313 4735 6341
rect 4682 6301 4688 6313
rect 4723 6310 4735 6313
rect 4769 6310 4781 6344
rect 9424 6341 9430 6353
rect 9385 6313 9430 6341
rect 4723 6304 4781 6310
rect 9424 6301 9430 6313
rect 9482 6301 9488 6353
rect 10096 6301 10102 6353
rect 10154 6341 10160 6353
rect 10195 6344 10253 6350
rect 10195 6341 10207 6344
rect 10154 6313 10207 6341
rect 10154 6301 10160 6313
rect 10195 6310 10207 6313
rect 10241 6310 10253 6344
rect 10195 6304 10253 6310
rect 10864 6301 10870 6353
rect 10922 6341 10928 6353
rect 10963 6344 11021 6350
rect 10963 6341 10975 6344
rect 10922 6313 10975 6341
rect 10922 6301 10928 6313
rect 10963 6310 10975 6313
rect 11009 6310 11021 6344
rect 10963 6304 11021 6310
rect 11632 6301 11638 6353
rect 11690 6341 11696 6353
rect 12211 6344 12269 6350
rect 12211 6341 12223 6344
rect 11690 6313 12223 6341
rect 11690 6301 11696 6313
rect 12211 6310 12223 6313
rect 12257 6310 12269 6344
rect 12211 6304 12269 6310
rect 12400 6301 12406 6353
rect 12458 6341 12464 6353
rect 12979 6344 13037 6350
rect 12979 6341 12991 6344
rect 12458 6313 12991 6341
rect 12458 6301 12464 6313
rect 12979 6310 12991 6313
rect 13025 6310 13037 6344
rect 12979 6304 13037 6310
rect 18736 6301 18742 6353
rect 18794 6341 18800 6353
rect 22963 6344 23021 6350
rect 22963 6341 22975 6344
rect 18794 6313 22975 6341
rect 18794 6301 18800 6313
rect 22963 6310 22975 6313
rect 23009 6310 23021 6344
rect 25648 6341 25654 6353
rect 25609 6313 25654 6341
rect 22963 6304 23021 6310
rect 25648 6301 25654 6313
rect 25706 6301 25712 6353
rect 26800 6341 26806 6353
rect 26761 6313 26806 6341
rect 26800 6301 26806 6313
rect 26858 6301 26864 6353
rect 29680 6341 29686 6353
rect 29641 6313 29686 6341
rect 29680 6301 29686 6313
rect 29738 6301 29744 6353
rect 31216 6341 31222 6353
rect 31177 6313 31222 6341
rect 31216 6301 31222 6313
rect 31274 6301 31280 6353
rect 36304 6341 36310 6353
rect 36265 6313 36310 6341
rect 36304 6301 36310 6313
rect 36362 6301 36368 6353
rect 38896 6341 38902 6353
rect 38857 6313 38902 6341
rect 38896 6301 38902 6313
rect 38954 6301 38960 6353
rect 40336 6341 40342 6353
rect 40297 6313 40342 6341
rect 40336 6301 40342 6313
rect 40394 6301 40400 6353
rect 41872 6341 41878 6353
rect 41833 6313 41878 6341
rect 41872 6301 41878 6313
rect 41930 6301 41936 6353
rect 45520 6341 45526 6353
rect 45481 6313 45526 6341
rect 45520 6301 45526 6313
rect 45578 6301 45584 6353
rect 46960 6341 46966 6353
rect 46921 6313 46966 6341
rect 46960 6301 46966 6313
rect 47018 6301 47024 6353
rect 47728 6341 47734 6353
rect 47689 6313 47734 6341
rect 47728 6301 47734 6313
rect 47786 6301 47792 6353
rect 48784 6301 48790 6353
rect 48842 6341 48848 6353
rect 49171 6344 49229 6350
rect 49171 6341 49183 6344
rect 48842 6313 49183 6341
rect 48842 6301 48848 6313
rect 49171 6310 49183 6313
rect 49217 6310 49229 6344
rect 49171 6304 49229 6310
rect 49552 6301 49558 6353
rect 49610 6341 49616 6353
rect 53314 6350 53342 6387
rect 56848 6375 56854 6387
rect 56906 6375 56912 6427
rect 49939 6344 49997 6350
rect 49939 6341 49951 6344
rect 49610 6313 49951 6341
rect 49610 6301 49616 6313
rect 49939 6310 49951 6313
rect 49985 6310 49997 6344
rect 49939 6304 49997 6310
rect 53299 6344 53357 6350
rect 53299 6310 53311 6344
rect 53345 6310 53357 6344
rect 53299 6304 53357 6310
rect 53968 6301 53974 6353
rect 54026 6341 54032 6353
rect 54451 6344 54509 6350
rect 54451 6341 54463 6344
rect 54026 6313 54463 6341
rect 54026 6301 54032 6313
rect 54451 6310 54463 6313
rect 54497 6310 54509 6344
rect 54451 6304 54509 6310
rect 55219 6344 55277 6350
rect 55219 6310 55231 6344
rect 55265 6310 55277 6344
rect 55219 6304 55277 6310
rect 55987 6344 56045 6350
rect 55987 6310 55999 6344
rect 56033 6310 56045 6344
rect 55987 6304 56045 6310
rect 57043 6344 57101 6350
rect 57043 6310 57055 6344
rect 57089 6310 57101 6344
rect 57043 6304 57101 6310
rect 57811 6344 57869 6350
rect 57811 6310 57823 6344
rect 57857 6341 57869 6344
rect 58096 6341 58102 6353
rect 57857 6313 58102 6341
rect 57857 6310 57869 6313
rect 57811 6304 57869 6310
rect 14707 6270 14765 6276
rect 14707 6236 14719 6270
rect 14753 6267 14765 6270
rect 15760 6267 15766 6279
rect 14753 6239 15766 6267
rect 14753 6236 14765 6239
rect 14707 6230 14765 6236
rect 15760 6227 15766 6239
rect 15818 6227 15824 6279
rect 41299 6270 41357 6276
rect 41299 6236 41311 6270
rect 41345 6267 41357 6270
rect 43792 6267 43798 6279
rect 41345 6239 43798 6267
rect 41345 6236 41357 6239
rect 41299 6230 41357 6236
rect 43792 6227 43798 6239
rect 43850 6227 43856 6279
rect 44080 6267 44086 6279
rect 44041 6239 44086 6267
rect 44080 6227 44086 6239
rect 44138 6227 44144 6279
rect 54352 6227 54358 6279
rect 54410 6267 54416 6279
rect 55234 6267 55262 6304
rect 54410 6239 55262 6267
rect 54410 6227 54416 6239
rect 14224 6153 14230 6205
rect 14282 6193 14288 6205
rect 14282 6165 15422 6193
rect 14282 6153 14288 6165
rect 5488 6079 5494 6131
rect 5546 6119 5552 6131
rect 5587 6122 5645 6128
rect 5587 6119 5599 6122
rect 5546 6091 5599 6119
rect 5546 6079 5552 6091
rect 5587 6088 5599 6091
rect 5633 6088 5645 6122
rect 5587 6082 5645 6088
rect 6256 6079 6262 6131
rect 6314 6119 6320 6131
rect 7027 6122 7085 6128
rect 7027 6119 7039 6122
rect 6314 6091 7039 6119
rect 6314 6079 6320 6091
rect 7027 6088 7039 6091
rect 7073 6088 7085 6122
rect 7027 6082 7085 6088
rect 14512 6079 14518 6131
rect 14570 6119 14576 6131
rect 15394 6128 15422 6165
rect 18928 6153 18934 6205
rect 18986 6193 18992 6205
rect 18986 6165 19934 6193
rect 18986 6153 18992 6165
rect 14611 6122 14669 6128
rect 14611 6119 14623 6122
rect 14570 6091 14623 6119
rect 14570 6079 14576 6091
rect 14611 6088 14623 6091
rect 14657 6088 14669 6122
rect 14611 6082 14669 6088
rect 15379 6122 15437 6128
rect 15379 6088 15391 6122
rect 15425 6088 15437 6122
rect 15379 6082 15437 6088
rect 16147 6122 16205 6128
rect 16147 6088 16159 6122
rect 16193 6119 16205 6122
rect 16528 6119 16534 6131
rect 16193 6091 16534 6119
rect 16193 6088 16205 6091
rect 16147 6082 16205 6088
rect 16528 6079 16534 6091
rect 16586 6079 16592 6131
rect 17584 6119 17590 6131
rect 17545 6091 17590 6119
rect 17584 6079 17590 6091
rect 17642 6079 17648 6131
rect 18256 6079 18262 6131
rect 18314 6119 18320 6131
rect 18355 6122 18413 6128
rect 18355 6119 18367 6122
rect 18314 6091 18367 6119
rect 18314 6079 18320 6091
rect 18355 6088 18367 6091
rect 18401 6088 18413 6122
rect 18355 6082 18413 6088
rect 19219 6122 19277 6128
rect 19219 6088 19231 6122
rect 19265 6119 19277 6122
rect 19312 6119 19318 6131
rect 19265 6091 19318 6119
rect 19265 6088 19277 6091
rect 19219 6082 19277 6088
rect 19312 6079 19318 6091
rect 19370 6079 19376 6131
rect 19906 6128 19934 6165
rect 20080 6153 20086 6205
rect 20138 6193 20144 6205
rect 20138 6165 21470 6193
rect 20138 6153 20144 6165
rect 19891 6122 19949 6128
rect 19891 6088 19903 6122
rect 19937 6088 19949 6122
rect 20656 6119 20662 6131
rect 20617 6091 20662 6119
rect 19891 6082 19949 6088
rect 20656 6079 20662 6091
rect 20714 6079 20720 6131
rect 21442 6128 21470 6165
rect 22288 6153 22294 6205
rect 22346 6193 22352 6205
rect 22346 6165 23678 6193
rect 22346 6153 22352 6165
rect 21427 6122 21485 6128
rect 21427 6088 21439 6122
rect 21473 6088 21485 6122
rect 21427 6082 21485 6088
rect 21520 6079 21526 6131
rect 21578 6119 21584 6131
rect 23650 6128 23678 6165
rect 31792 6153 31798 6205
rect 31850 6193 31856 6205
rect 31850 6165 33470 6193
rect 31850 6153 31856 6165
rect 22867 6122 22925 6128
rect 22867 6119 22879 6122
rect 21578 6091 22879 6119
rect 21578 6079 21584 6091
rect 22867 6088 22879 6091
rect 22913 6088 22925 6122
rect 22867 6082 22925 6088
rect 23635 6122 23693 6128
rect 23635 6088 23647 6122
rect 23681 6088 23693 6122
rect 23635 6082 23693 6088
rect 24016 6079 24022 6131
rect 24074 6119 24080 6131
rect 24403 6122 24461 6128
rect 24403 6119 24415 6122
rect 24074 6091 24415 6119
rect 24074 6079 24080 6091
rect 24403 6088 24415 6091
rect 24449 6088 24461 6122
rect 24403 6082 24461 6088
rect 26320 6079 26326 6131
rect 26378 6119 26384 6131
rect 28147 6122 28205 6128
rect 28147 6119 28159 6122
rect 26378 6091 28159 6119
rect 26378 6079 26384 6091
rect 28147 6088 28159 6091
rect 28193 6088 28205 6122
rect 28147 6082 28205 6088
rect 28915 6122 28973 6128
rect 28915 6088 28927 6122
rect 28961 6119 28973 6122
rect 29008 6119 29014 6131
rect 28961 6091 29014 6119
rect 28961 6088 28973 6091
rect 28915 6082 28973 6088
rect 29008 6079 29014 6091
rect 29066 6079 29072 6131
rect 29776 6079 29782 6131
rect 29834 6119 29840 6131
rect 33442 6128 33470 6165
rect 33712 6153 33718 6205
rect 33770 6193 33776 6205
rect 33770 6165 35102 6193
rect 33770 6153 33776 6165
rect 30643 6122 30701 6128
rect 30643 6119 30655 6122
rect 29834 6091 30655 6119
rect 29834 6079 29840 6091
rect 30643 6088 30655 6091
rect 30689 6088 30701 6122
rect 30643 6082 30701 6088
rect 33427 6122 33485 6128
rect 33427 6088 33439 6122
rect 33473 6088 33485 6122
rect 34288 6119 34294 6131
rect 34249 6091 34294 6119
rect 33427 6082 33485 6088
rect 34288 6079 34294 6091
rect 34346 6079 34352 6131
rect 35074 6128 35102 6165
rect 40624 6153 40630 6205
rect 40682 6193 40688 6205
rect 40682 6165 41342 6193
rect 40682 6153 40688 6165
rect 35059 6122 35117 6128
rect 35059 6088 35071 6122
rect 35105 6088 35117 6122
rect 35059 6082 35117 6088
rect 37171 6122 37229 6128
rect 37171 6088 37183 6122
rect 37217 6119 37229 6122
rect 37264 6119 37270 6131
rect 37217 6091 37270 6119
rect 37217 6088 37229 6091
rect 37171 6082 37229 6088
rect 37264 6079 37270 6091
rect 37322 6079 37328 6131
rect 39184 6079 39190 6131
rect 39242 6119 39248 6131
rect 41203 6122 41261 6128
rect 41203 6119 41215 6122
rect 39242 6091 41215 6119
rect 39242 6079 39248 6091
rect 41203 6088 41215 6091
rect 41249 6088 41261 6122
rect 41314 6119 41342 6165
rect 42160 6153 42166 6205
rect 42218 6193 42224 6205
rect 42218 6165 44030 6193
rect 42218 6153 42224 6165
rect 44002 6128 44030 6165
rect 51568 6153 51574 6205
rect 51626 6193 51632 6205
rect 51626 6165 52382 6193
rect 51626 6153 51632 6165
rect 42835 6122 42893 6128
rect 42835 6119 42847 6122
rect 41314 6091 42847 6119
rect 41203 6082 41261 6088
rect 42835 6088 42847 6091
rect 42881 6088 42893 6122
rect 42835 6082 42893 6088
rect 43987 6122 44045 6128
rect 43987 6088 43999 6122
rect 44033 6088 44045 6122
rect 43987 6082 44045 6088
rect 44176 6079 44182 6131
rect 44234 6119 44240 6131
rect 44755 6122 44813 6128
rect 44755 6119 44767 6122
rect 44234 6091 44767 6119
rect 44234 6079 44240 6091
rect 44755 6088 44767 6091
rect 44801 6088 44813 6122
rect 44755 6082 44813 6088
rect 49744 6079 49750 6131
rect 49802 6119 49808 6131
rect 50803 6122 50861 6128
rect 50803 6119 50815 6122
rect 49802 6091 50815 6119
rect 49802 6079 49808 6091
rect 50803 6088 50815 6091
rect 50849 6088 50861 6122
rect 50803 6082 50861 6088
rect 51088 6079 51094 6131
rect 51146 6119 51152 6131
rect 52354 6128 52382 6165
rect 55024 6153 55030 6205
rect 55082 6193 55088 6205
rect 56002 6193 56030 6304
rect 57058 6267 57086 6304
rect 58096 6301 58102 6313
rect 58154 6301 58160 6353
rect 58864 6267 58870 6279
rect 57058 6239 58870 6267
rect 58864 6227 58870 6239
rect 58922 6227 58928 6279
rect 55082 6165 56030 6193
rect 55082 6153 55088 6165
rect 51667 6122 51725 6128
rect 51667 6119 51679 6122
rect 51146 6091 51679 6119
rect 51146 6079 51152 6091
rect 51667 6088 51679 6091
rect 51713 6088 51725 6122
rect 51667 6082 51725 6088
rect 52339 6122 52397 6128
rect 52339 6088 52351 6122
rect 52385 6088 52397 6122
rect 52339 6082 52397 6088
rect 1152 6020 58848 6042
rect 1152 5968 19654 6020
rect 19706 5968 19718 6020
rect 19770 5968 19782 6020
rect 19834 5968 19846 6020
rect 19898 5968 50374 6020
rect 50426 5968 50438 6020
rect 50490 5968 50502 6020
rect 50554 5968 50566 6020
rect 50618 5968 58848 6020
rect 1152 5946 58848 5968
rect 3568 5857 3574 5909
rect 3626 5897 3632 5909
rect 7792 5897 7798 5909
rect 3626 5869 7798 5897
rect 3626 5857 3632 5869
rect 7792 5857 7798 5869
rect 7850 5857 7856 5909
rect 44080 5857 44086 5909
rect 44138 5897 44144 5909
rect 44138 5869 47534 5897
rect 44138 5857 44144 5869
rect 47506 5823 47534 5869
rect 49264 5857 49270 5909
rect 49322 5897 49328 5909
rect 49648 5897 49654 5909
rect 49322 5869 49654 5897
rect 49322 5857 49328 5869
rect 49648 5857 49654 5869
rect 49706 5857 49712 5909
rect 47506 5795 55454 5823
rect 7024 5709 7030 5761
rect 7082 5749 7088 5761
rect 44944 5749 44950 5761
rect 7082 5721 44950 5749
rect 7082 5709 7088 5721
rect 44944 5709 44950 5721
rect 45002 5709 45008 5761
rect 55426 5758 55454 5795
rect 55411 5752 55469 5758
rect 55411 5718 55423 5752
rect 55457 5718 55469 5752
rect 55411 5712 55469 5718
rect 1072 5635 1078 5687
rect 1130 5675 1136 5687
rect 1555 5678 1613 5684
rect 1555 5675 1567 5678
rect 1130 5647 1567 5675
rect 1130 5635 1136 5647
rect 1555 5644 1567 5647
rect 1601 5644 1613 5678
rect 1555 5638 1613 5644
rect 2896 5635 2902 5687
rect 2954 5675 2960 5687
rect 4435 5678 4493 5684
rect 2954 5647 2999 5675
rect 2954 5635 2960 5647
rect 4435 5644 4447 5678
rect 4481 5675 4493 5678
rect 4912 5675 4918 5687
rect 4481 5647 4918 5675
rect 4481 5644 4493 5647
rect 4435 5638 4493 5644
rect 4912 5635 4918 5647
rect 4970 5635 4976 5687
rect 5104 5675 5110 5687
rect 5065 5647 5110 5675
rect 5104 5635 5110 5647
rect 5162 5635 5168 5687
rect 5776 5635 5782 5687
rect 5834 5675 5840 5687
rect 6832 5675 6838 5687
rect 5834 5647 6014 5675
rect 6793 5647 6838 5675
rect 5834 5635 5840 5647
rect 5986 5610 6014 5647
rect 6832 5635 6838 5647
rect 6890 5635 6896 5687
rect 7216 5635 7222 5687
rect 7274 5675 7280 5687
rect 7603 5678 7661 5684
rect 7603 5675 7615 5678
rect 7274 5647 7615 5675
rect 7274 5635 7280 5647
rect 7603 5644 7615 5647
rect 7649 5644 7661 5678
rect 7603 5638 7661 5644
rect 7987 5678 8045 5684
rect 7987 5644 7999 5678
rect 8033 5675 8045 5678
rect 8371 5678 8429 5684
rect 8371 5675 8383 5678
rect 8033 5647 8383 5675
rect 8033 5644 8045 5647
rect 7987 5638 8045 5644
rect 8371 5644 8383 5647
rect 8417 5644 8429 5678
rect 8371 5638 8429 5644
rect 8752 5635 8758 5687
rect 8810 5675 8816 5687
rect 9619 5678 9677 5684
rect 9619 5675 9631 5678
rect 8810 5647 9631 5675
rect 8810 5635 8816 5647
rect 9619 5644 9631 5647
rect 9665 5644 9677 5678
rect 9619 5638 9677 5644
rect 10192 5635 10198 5687
rect 10250 5675 10256 5687
rect 10387 5678 10445 5684
rect 10387 5675 10399 5678
rect 10250 5647 10399 5675
rect 10250 5635 10256 5647
rect 10387 5644 10399 5647
rect 10433 5644 10445 5678
rect 10387 5638 10445 5644
rect 10480 5635 10486 5687
rect 10538 5675 10544 5687
rect 11155 5678 11213 5684
rect 11155 5675 11167 5678
rect 10538 5647 11167 5675
rect 10538 5635 10544 5647
rect 11155 5644 11167 5647
rect 11201 5644 11213 5678
rect 12592 5675 12598 5687
rect 12553 5647 12598 5675
rect 11155 5638 11213 5644
rect 12592 5635 12598 5647
rect 12650 5635 12656 5687
rect 13360 5675 13366 5687
rect 13321 5647 13366 5675
rect 13360 5635 13366 5647
rect 13418 5635 13424 5687
rect 14992 5675 14998 5687
rect 14953 5647 14998 5675
rect 14992 5635 14998 5647
rect 15050 5635 15056 5687
rect 15856 5675 15862 5687
rect 15817 5647 15862 5675
rect 15856 5635 15862 5647
rect 15914 5635 15920 5687
rect 16144 5635 16150 5687
rect 16202 5675 16208 5687
rect 16531 5678 16589 5684
rect 16531 5675 16543 5678
rect 16202 5647 16543 5675
rect 16202 5635 16208 5647
rect 16531 5644 16543 5647
rect 16577 5644 16589 5678
rect 16531 5638 16589 5644
rect 17296 5635 17302 5687
rect 17354 5675 17360 5687
rect 18736 5675 18742 5687
rect 17354 5647 17399 5675
rect 18697 5647 18742 5675
rect 17354 5635 17360 5647
rect 18736 5635 18742 5647
rect 18794 5635 18800 5687
rect 20176 5675 20182 5687
rect 20137 5647 20182 5675
rect 20176 5635 20182 5647
rect 20234 5635 20240 5687
rect 20560 5635 20566 5687
rect 20618 5675 20624 5687
rect 20947 5678 21005 5684
rect 20947 5675 20959 5678
rect 20618 5647 20959 5675
rect 20618 5635 20624 5647
rect 20947 5644 20959 5647
rect 20993 5644 21005 5678
rect 20947 5638 21005 5644
rect 21619 5678 21677 5684
rect 21619 5644 21631 5678
rect 21665 5675 21677 5678
rect 21715 5678 21773 5684
rect 21715 5675 21727 5678
rect 21665 5647 21727 5675
rect 21665 5644 21677 5647
rect 21619 5638 21677 5644
rect 21715 5644 21727 5647
rect 21761 5644 21773 5678
rect 21715 5638 21773 5644
rect 21808 5635 21814 5687
rect 21866 5675 21872 5687
rect 22483 5678 22541 5684
rect 22483 5675 22495 5678
rect 21866 5647 22495 5675
rect 21866 5635 21872 5647
rect 22483 5644 22495 5647
rect 22529 5644 22541 5678
rect 22483 5638 22541 5644
rect 23056 5635 23062 5687
rect 23114 5675 23120 5687
rect 23251 5678 23309 5684
rect 23251 5675 23263 5678
rect 23114 5647 23263 5675
rect 23114 5635 23120 5647
rect 23251 5644 23263 5647
rect 23297 5644 23309 5678
rect 23251 5638 23309 5644
rect 23440 5635 23446 5687
rect 23498 5675 23504 5687
rect 24019 5678 24077 5684
rect 24019 5675 24031 5678
rect 23498 5647 24031 5675
rect 23498 5635 23504 5647
rect 24019 5644 24031 5647
rect 24065 5644 24077 5678
rect 24019 5638 24077 5644
rect 24592 5635 24598 5687
rect 24650 5675 24656 5687
rect 25459 5678 25517 5684
rect 25459 5675 25471 5678
rect 24650 5647 25471 5675
rect 24650 5635 24656 5647
rect 25459 5644 25471 5647
rect 25505 5644 25517 5678
rect 26224 5675 26230 5687
rect 26185 5647 26230 5675
rect 25459 5638 25517 5644
rect 26224 5635 26230 5647
rect 26282 5635 26288 5687
rect 26611 5678 26669 5684
rect 26611 5644 26623 5678
rect 26657 5675 26669 5678
rect 26995 5678 27053 5684
rect 26995 5675 27007 5678
rect 26657 5647 27007 5675
rect 26657 5644 26669 5647
rect 26611 5638 26669 5644
rect 26995 5644 27007 5647
rect 27041 5644 27053 5678
rect 26995 5638 27053 5644
rect 27376 5635 27382 5687
rect 27434 5675 27440 5687
rect 27763 5678 27821 5684
rect 27763 5675 27775 5678
rect 27434 5647 27775 5675
rect 27434 5635 27440 5647
rect 27763 5644 27775 5647
rect 27809 5644 27821 5678
rect 27763 5638 27821 5644
rect 27856 5635 27862 5687
rect 27914 5675 27920 5687
rect 28531 5678 28589 5684
rect 28531 5675 28543 5678
rect 27914 5647 28543 5675
rect 27914 5635 27920 5647
rect 28531 5644 28543 5647
rect 28577 5644 28589 5678
rect 28531 5638 28589 5644
rect 28816 5635 28822 5687
rect 28874 5675 28880 5687
rect 29299 5678 29357 5684
rect 29299 5675 29311 5678
rect 28874 5647 29311 5675
rect 28874 5635 28880 5647
rect 29299 5644 29311 5647
rect 29345 5644 29357 5678
rect 29299 5638 29357 5644
rect 30256 5635 30262 5687
rect 30314 5675 30320 5687
rect 30739 5678 30797 5684
rect 30739 5675 30751 5678
rect 30314 5647 30751 5675
rect 30314 5635 30320 5647
rect 30739 5644 30751 5647
rect 30785 5644 30797 5678
rect 30739 5638 30797 5644
rect 30832 5635 30838 5687
rect 30890 5675 30896 5687
rect 31507 5678 31565 5684
rect 31507 5675 31519 5678
rect 30890 5647 31519 5675
rect 30890 5635 30896 5647
rect 31507 5644 31519 5647
rect 31553 5644 31565 5678
rect 31507 5638 31565 5644
rect 31696 5635 31702 5687
rect 31754 5675 31760 5687
rect 32275 5678 32333 5684
rect 32275 5675 32287 5678
rect 31754 5647 32287 5675
rect 31754 5635 31760 5647
rect 32275 5644 32287 5647
rect 32321 5644 32333 5678
rect 33136 5675 33142 5687
rect 33097 5647 33142 5675
rect 32275 5638 32333 5644
rect 33136 5635 33142 5647
rect 33194 5635 33200 5687
rect 33232 5635 33238 5687
rect 33290 5675 33296 5687
rect 33811 5678 33869 5684
rect 33811 5675 33823 5678
rect 33290 5647 33823 5675
rect 33290 5635 33296 5647
rect 33811 5644 33823 5647
rect 33857 5644 33869 5678
rect 34672 5675 34678 5687
rect 34633 5647 34678 5675
rect 33811 5638 33869 5644
rect 34672 5635 34678 5647
rect 34730 5635 34736 5687
rect 36016 5675 36022 5687
rect 35977 5647 36022 5675
rect 36016 5635 36022 5647
rect 36074 5635 36080 5687
rect 36208 5635 36214 5687
rect 36266 5675 36272 5687
rect 36787 5678 36845 5684
rect 36787 5675 36799 5678
rect 36266 5647 36799 5675
rect 36266 5635 36272 5647
rect 36787 5644 36799 5647
rect 36833 5644 36845 5678
rect 37552 5675 37558 5687
rect 37513 5647 37558 5675
rect 36787 5638 36845 5644
rect 37552 5635 37558 5647
rect 37610 5635 37616 5687
rect 37939 5678 37997 5684
rect 37939 5644 37951 5678
rect 37985 5675 37997 5678
rect 38323 5678 38381 5684
rect 38323 5675 38335 5678
rect 37985 5647 38335 5675
rect 37985 5644 37997 5647
rect 37939 5638 37997 5644
rect 38323 5644 38335 5647
rect 38369 5644 38381 5678
rect 39088 5675 39094 5687
rect 39049 5647 39094 5675
rect 38323 5638 38381 5644
rect 39088 5635 39094 5647
rect 39146 5635 39152 5687
rect 39280 5635 39286 5687
rect 39338 5675 39344 5687
rect 39859 5678 39917 5684
rect 39859 5675 39871 5678
rect 39338 5647 39871 5675
rect 39338 5635 39344 5647
rect 39859 5644 39871 5647
rect 39905 5644 39917 5678
rect 39859 5638 39917 5644
rect 40720 5635 40726 5687
rect 40778 5675 40784 5687
rect 41299 5678 41357 5684
rect 41299 5675 41311 5678
rect 40778 5647 41311 5675
rect 40778 5635 40784 5647
rect 41299 5644 41311 5647
rect 41345 5644 41357 5678
rect 41299 5638 41357 5644
rect 41776 5635 41782 5687
rect 41834 5675 41840 5687
rect 42067 5678 42125 5684
rect 42067 5675 42079 5678
rect 41834 5647 42079 5675
rect 41834 5635 41840 5647
rect 42067 5644 42079 5647
rect 42113 5644 42125 5678
rect 42067 5638 42125 5644
rect 42256 5635 42262 5687
rect 42314 5675 42320 5687
rect 42835 5678 42893 5684
rect 42835 5675 42847 5678
rect 42314 5647 42847 5675
rect 42314 5635 42320 5647
rect 42835 5644 42847 5647
rect 42881 5644 42893 5678
rect 42835 5638 42893 5644
rect 43216 5635 43222 5687
rect 43274 5675 43280 5687
rect 43603 5678 43661 5684
rect 43603 5675 43615 5678
rect 43274 5647 43615 5675
rect 43274 5635 43280 5647
rect 43603 5644 43615 5647
rect 43649 5644 43661 5678
rect 43603 5638 43661 5644
rect 43696 5635 43702 5687
rect 43754 5675 43760 5687
rect 44371 5678 44429 5684
rect 44371 5675 44383 5678
rect 43754 5647 44383 5675
rect 43754 5635 43760 5647
rect 44371 5644 44383 5647
rect 44417 5644 44429 5678
rect 45136 5675 45142 5687
rect 45097 5647 45142 5675
rect 44371 5638 44429 5644
rect 45136 5635 45142 5647
rect 45194 5635 45200 5687
rect 46096 5635 46102 5687
rect 46154 5675 46160 5687
rect 46579 5678 46637 5684
rect 46579 5675 46591 5678
rect 46154 5647 46591 5675
rect 46154 5635 46160 5647
rect 46579 5644 46591 5647
rect 46625 5644 46637 5678
rect 46579 5638 46637 5644
rect 46672 5635 46678 5687
rect 46730 5675 46736 5687
rect 47347 5678 47405 5684
rect 47347 5675 47359 5678
rect 46730 5647 47359 5675
rect 46730 5635 46736 5647
rect 47347 5644 47359 5647
rect 47393 5644 47405 5678
rect 47347 5638 47405 5644
rect 47536 5635 47542 5687
rect 47594 5675 47600 5687
rect 48115 5678 48173 5684
rect 48115 5675 48127 5678
rect 47594 5647 48127 5675
rect 47594 5635 47600 5647
rect 48115 5644 48127 5647
rect 48161 5644 48173 5678
rect 48976 5675 48982 5687
rect 48937 5647 48982 5675
rect 48115 5638 48173 5644
rect 48976 5635 48982 5647
rect 49034 5635 49040 5687
rect 49648 5675 49654 5687
rect 49609 5647 49654 5675
rect 49648 5635 49654 5647
rect 49706 5635 49712 5687
rect 50515 5678 50573 5684
rect 50515 5644 50527 5678
rect 50561 5675 50573 5678
rect 50704 5675 50710 5687
rect 50561 5647 50710 5675
rect 50561 5644 50573 5647
rect 50515 5638 50573 5644
rect 50704 5635 50710 5647
rect 50762 5635 50768 5687
rect 52144 5675 52150 5687
rect 52105 5647 52150 5675
rect 52144 5635 52150 5647
rect 52202 5635 52208 5687
rect 52528 5635 52534 5687
rect 52586 5675 52592 5687
rect 52915 5678 52973 5684
rect 52915 5675 52927 5678
rect 52586 5647 52927 5675
rect 52586 5635 52592 5647
rect 52915 5644 52927 5647
rect 52961 5644 52973 5678
rect 53680 5675 53686 5687
rect 53641 5647 53686 5675
rect 52915 5638 52973 5644
rect 53680 5635 53686 5647
rect 53738 5635 53744 5687
rect 54451 5678 54509 5684
rect 54451 5644 54463 5678
rect 54497 5644 54509 5678
rect 54451 5638 54509 5644
rect 55987 5678 56045 5684
rect 55987 5644 55999 5678
rect 56033 5644 56045 5678
rect 57424 5675 57430 5687
rect 57385 5647 57430 5675
rect 55987 5638 56045 5644
rect 5971 5604 6029 5610
rect 5971 5570 5983 5604
rect 6017 5570 6029 5604
rect 5971 5564 6029 5570
rect 6067 5604 6125 5610
rect 6067 5570 6079 5604
rect 6113 5601 6125 5604
rect 46288 5601 46294 5613
rect 6113 5573 46294 5601
rect 6113 5570 6125 5573
rect 6067 5564 6125 5570
rect 5779 5530 5837 5536
rect 5779 5496 5791 5530
rect 5825 5527 5837 5530
rect 6082 5527 6110 5564
rect 46288 5561 46294 5573
rect 46346 5561 46352 5613
rect 53584 5561 53590 5613
rect 53642 5601 53648 5613
rect 54466 5601 54494 5638
rect 53642 5573 54494 5601
rect 56002 5601 56030 5638
rect 57424 5635 57430 5647
rect 57482 5635 57488 5687
rect 59632 5601 59638 5613
rect 56002 5573 59638 5601
rect 53642 5561 53648 5573
rect 59632 5561 59638 5573
rect 59690 5561 59696 5613
rect 5825 5499 6110 5527
rect 5825 5496 5837 5499
rect 5779 5490 5837 5496
rect 7600 5487 7606 5539
rect 7658 5527 7664 5539
rect 7987 5530 8045 5536
rect 7987 5527 7999 5530
rect 7658 5499 7999 5527
rect 7658 5487 7664 5499
rect 7987 5496 7999 5499
rect 8033 5496 8045 5530
rect 7987 5490 8045 5496
rect 21619 5530 21677 5536
rect 21619 5496 21631 5530
rect 21665 5527 21677 5530
rect 21712 5527 21718 5539
rect 21665 5499 21718 5527
rect 21665 5496 21677 5499
rect 21619 5490 21677 5496
rect 21712 5487 21718 5499
rect 21770 5487 21776 5539
rect 26032 5487 26038 5539
rect 26090 5527 26096 5539
rect 26611 5530 26669 5536
rect 26611 5527 26623 5530
rect 26090 5499 26623 5527
rect 26090 5487 26096 5499
rect 26611 5496 26623 5499
rect 26657 5496 26669 5530
rect 26611 5490 26669 5496
rect 37456 5487 37462 5539
rect 37514 5527 37520 5539
rect 37939 5530 37997 5536
rect 37939 5527 37951 5530
rect 37514 5499 37951 5527
rect 37514 5487 37520 5499
rect 37939 5496 37951 5499
rect 37985 5496 37997 5530
rect 37939 5490 37997 5496
rect 3760 5413 3766 5465
rect 3818 5453 3824 5465
rect 8368 5453 8374 5465
rect 3818 5425 8374 5453
rect 3818 5413 3824 5425
rect 8368 5413 8374 5425
rect 8426 5413 8432 5465
rect 1152 5354 58848 5376
rect 1152 5302 4294 5354
rect 4346 5302 4358 5354
rect 4410 5302 4422 5354
rect 4474 5302 4486 5354
rect 4538 5302 35014 5354
rect 35066 5302 35078 5354
rect 35130 5302 35142 5354
rect 35194 5302 35206 5354
rect 35258 5302 58848 5354
rect 1152 5280 58848 5302
rect 5008 5191 5014 5243
rect 5066 5231 5072 5243
rect 7507 5234 7565 5240
rect 7507 5231 7519 5234
rect 5066 5203 7519 5231
rect 5066 5191 5072 5203
rect 7507 5200 7519 5203
rect 7553 5231 7565 5234
rect 7699 5234 7757 5240
rect 7699 5231 7711 5234
rect 7553 5203 7711 5231
rect 7553 5200 7565 5203
rect 7507 5194 7565 5200
rect 7699 5200 7711 5203
rect 7745 5200 7757 5234
rect 7699 5194 7757 5200
rect 8467 5234 8525 5240
rect 8467 5200 8479 5234
rect 8513 5231 8525 5234
rect 8513 5203 8654 5231
rect 8513 5200 8525 5203
rect 8467 5194 8525 5200
rect 8626 5143 8654 5203
rect 304 4969 310 5021
rect 362 5009 368 5021
rect 1555 5012 1613 5018
rect 1555 5009 1567 5012
rect 362 4981 1567 5009
rect 362 4969 368 4981
rect 1555 4978 1567 4981
rect 1601 4978 1613 5012
rect 1555 4972 1613 4978
rect 1840 4969 1846 5021
rect 1898 5009 1904 5021
rect 2323 5012 2381 5018
rect 2323 5009 2335 5012
rect 1898 4981 2335 5009
rect 1898 4969 1904 4981
rect 2323 4978 2335 4981
rect 2369 4978 2381 5012
rect 3088 5009 3094 5021
rect 3049 4981 3094 5009
rect 2323 4972 2381 4978
rect 3088 4969 3094 4981
rect 3146 4969 3152 5021
rect 4144 5009 4150 5021
rect 4105 4981 4150 5009
rect 4144 4969 4150 4981
rect 4202 4969 4208 5021
rect 5392 5009 5398 5021
rect 5353 4981 5398 5009
rect 5392 4969 5398 4981
rect 5450 4969 5456 5021
rect 6064 4969 6070 5021
rect 6122 5009 6128 5021
rect 6931 5012 6989 5018
rect 6931 5009 6943 5012
rect 6122 4981 6943 5009
rect 6122 4969 6128 4981
rect 6931 4978 6943 4981
rect 6977 4978 6989 5012
rect 9232 5009 9238 5021
rect 9193 4981 9238 5009
rect 6931 4972 6989 4978
rect 9232 4969 9238 4981
rect 9290 4969 9296 5021
rect 10000 5009 10006 5021
rect 9961 4981 10006 5009
rect 10000 4969 10006 4981
rect 10058 4969 10064 5021
rect 10576 4969 10582 5021
rect 10634 5009 10640 5021
rect 10771 5012 10829 5018
rect 10771 5009 10783 5012
rect 10634 4981 10783 5009
rect 10634 4969 10640 4981
rect 10771 4978 10783 4981
rect 10817 4978 10829 5012
rect 10771 4972 10829 4978
rect 11824 4969 11830 5021
rect 11882 5009 11888 5021
rect 12211 5012 12269 5018
rect 12211 5009 12223 5012
rect 11882 4981 12223 5009
rect 11882 4969 11888 4981
rect 12211 4978 12223 4981
rect 12257 4978 12269 5012
rect 12976 5009 12982 5021
rect 12937 4981 12982 5009
rect 12211 4972 12269 4978
rect 12976 4969 12982 4981
rect 13034 4969 13040 5021
rect 13936 5009 13942 5021
rect 13897 4981 13942 5009
rect 13936 4969 13942 4981
rect 13994 4969 14000 5021
rect 14416 4969 14422 5021
rect 14474 5009 14480 5021
rect 14707 5012 14765 5018
rect 14707 5009 14719 5012
rect 14474 4981 14719 5009
rect 14474 4969 14480 4981
rect 14707 4978 14719 4981
rect 14753 4978 14765 5012
rect 14707 4972 14765 4978
rect 14800 4969 14806 5021
rect 14858 5009 14864 5021
rect 15475 5012 15533 5018
rect 15475 5009 15487 5012
rect 14858 4981 15487 5009
rect 14858 4969 14864 4981
rect 15475 4978 15487 4981
rect 15521 4978 15533 5012
rect 15475 4972 15533 4978
rect 16339 5012 16397 5018
rect 16339 4978 16351 5012
rect 16385 5009 16397 5012
rect 16432 5009 16438 5021
rect 16385 4981 16438 5009
rect 16385 4978 16397 4981
rect 16339 4972 16397 4978
rect 16432 4969 16438 4981
rect 16490 4969 16496 5021
rect 17488 5009 17494 5021
rect 17449 4981 17494 5009
rect 17488 4969 17494 4981
rect 17546 4969 17552 5021
rect 17968 4969 17974 5021
rect 18026 5009 18032 5021
rect 18259 5012 18317 5018
rect 18259 5009 18271 5012
rect 18026 4981 18271 5009
rect 18026 4969 18032 4981
rect 18259 4978 18271 4981
rect 18305 4978 18317 5012
rect 19024 5009 19030 5021
rect 18985 4981 19030 5009
rect 18259 4972 18317 4978
rect 19024 4969 19030 4981
rect 19082 4969 19088 5021
rect 19120 4969 19126 5021
rect 19178 5009 19184 5021
rect 19795 5012 19853 5018
rect 19795 5009 19807 5012
rect 19178 4981 19807 5009
rect 19178 4969 19184 4981
rect 19795 4978 19807 4981
rect 19841 4978 19853 5012
rect 19795 4972 19853 4978
rect 20464 4969 20470 5021
rect 20522 5009 20528 5021
rect 20563 5012 20621 5018
rect 20563 5009 20575 5012
rect 20522 4981 20575 5009
rect 20522 4969 20528 4981
rect 20563 4978 20575 4981
rect 20609 4978 20621 5012
rect 20563 4972 20621 4978
rect 21232 4969 21238 5021
rect 21290 5009 21296 5021
rect 21331 5012 21389 5018
rect 21331 5009 21343 5012
rect 21290 4981 21343 5009
rect 21290 4969 21296 4981
rect 21331 4978 21343 4981
rect 21377 4978 21389 5012
rect 22768 5009 22774 5021
rect 22729 4981 22774 5009
rect 21331 4972 21389 4978
rect 22768 4969 22774 4981
rect 22826 4969 22832 5021
rect 23536 5009 23542 5021
rect 23497 4981 23542 5009
rect 23536 4969 23542 4981
rect 23594 4969 23600 5021
rect 24307 5012 24365 5018
rect 24307 4978 24319 5012
rect 24353 4978 24365 5012
rect 25072 5009 25078 5021
rect 25033 4981 25078 5009
rect 24307 4972 24365 4978
rect 7942 4947 7994 4953
rect 23152 4895 23158 4947
rect 23210 4935 23216 4947
rect 24322 4935 24350 4972
rect 25072 4969 25078 4981
rect 25130 4969 25136 5021
rect 25840 5009 25846 5021
rect 25801 4981 25846 5009
rect 25840 4969 25846 4981
rect 25898 4969 25904 5021
rect 26608 5009 26614 5021
rect 26569 4981 26614 5009
rect 26608 4969 26614 4981
rect 26666 4969 26672 5021
rect 28048 5009 28054 5021
rect 28009 4981 28054 5009
rect 28048 4969 28054 4981
rect 28106 4969 28112 5021
rect 28912 5009 28918 5021
rect 28873 4981 28918 5009
rect 28912 4969 28918 4981
rect 28970 4969 28976 5021
rect 29296 4969 29302 5021
rect 29354 5009 29360 5021
rect 29587 5012 29645 5018
rect 29587 5009 29599 5012
rect 29354 4981 29599 5009
rect 29354 4969 29360 4981
rect 29587 4978 29599 4981
rect 29633 4978 29645 5012
rect 30352 5009 30358 5021
rect 30313 4981 30358 5009
rect 29587 4972 29645 4978
rect 30352 4969 30358 4981
rect 30410 4969 30416 5021
rect 31120 5009 31126 5021
rect 31081 4981 31126 5009
rect 31120 4969 31126 4981
rect 31178 4969 31184 5021
rect 31888 5009 31894 5021
rect 31849 4981 31894 5009
rect 31888 4969 31894 4981
rect 31946 4969 31952 5021
rect 33328 5009 33334 5021
rect 33289 4981 33334 5009
rect 33328 4969 33334 4981
rect 33386 4969 33392 5021
rect 34096 5009 34102 5021
rect 34057 4981 34102 5009
rect 34096 4969 34102 4981
rect 34154 4969 34160 5021
rect 34864 5009 34870 5021
rect 34825 4981 34870 5009
rect 34864 4969 34870 4981
rect 34922 4969 34928 5021
rect 35635 5012 35693 5018
rect 35635 4978 35647 5012
rect 35681 4978 35693 5012
rect 35635 4972 35693 4978
rect 23210 4907 24350 4935
rect 23210 4895 23216 4907
rect 34576 4895 34582 4947
rect 34634 4935 34640 4947
rect 35650 4935 35678 4972
rect 36112 4969 36118 5021
rect 36170 5009 36176 5021
rect 36403 5012 36461 5018
rect 36403 5009 36415 5012
rect 36170 4981 36415 5009
rect 36170 4969 36176 4981
rect 36403 4978 36415 4981
rect 36449 4978 36461 5012
rect 36403 4972 36461 4978
rect 36880 4969 36886 5021
rect 36938 5009 36944 5021
rect 37171 5012 37229 5018
rect 37171 5009 37183 5012
rect 36938 4981 37183 5009
rect 36938 4969 36944 4981
rect 37171 4978 37183 4981
rect 37217 4978 37229 5012
rect 38608 5009 38614 5021
rect 38569 4981 38614 5009
rect 37171 4972 37229 4978
rect 38608 4969 38614 4981
rect 38666 4969 38672 5021
rect 39376 5009 39382 5021
rect 39337 4981 39382 5009
rect 39376 4969 39382 4981
rect 39434 4969 39440 5021
rect 40144 5009 40150 5021
rect 40105 4981 40150 5009
rect 40144 4969 40150 4981
rect 40202 4969 40208 5021
rect 40912 5009 40918 5021
rect 40873 4981 40918 5009
rect 40912 4969 40918 4981
rect 40970 4969 40976 5021
rect 41680 5009 41686 5021
rect 41641 4981 41686 5009
rect 41680 4969 41686 4981
rect 41738 4969 41744 5021
rect 42064 4969 42070 5021
rect 42122 5009 42128 5021
rect 42451 5012 42509 5018
rect 42451 5009 42463 5012
rect 42122 4981 42463 5009
rect 42122 4969 42128 4981
rect 42451 4978 42463 4981
rect 42497 4978 42509 5012
rect 42451 4972 42509 4978
rect 43312 4969 43318 5021
rect 43370 5009 43376 5021
rect 43891 5012 43949 5018
rect 43891 5009 43903 5012
rect 43370 4981 43903 5009
rect 43370 4969 43376 4981
rect 43891 4978 43903 4981
rect 43937 4978 43949 5012
rect 44752 5009 44758 5021
rect 44713 4981 44758 5009
rect 43891 4972 43949 4978
rect 44752 4969 44758 4981
rect 44810 4969 44816 5021
rect 45424 5009 45430 5021
rect 45385 4981 45430 5009
rect 45424 4969 45430 4981
rect 45482 4969 45488 5021
rect 46192 5009 46198 5021
rect 46153 4981 46198 5009
rect 46192 4969 46198 4981
rect 46250 4969 46256 5021
rect 46288 4969 46294 5021
rect 46346 5009 46352 5021
rect 46963 5012 47021 5018
rect 46963 5009 46975 5012
rect 46346 4981 46975 5009
rect 46346 4969 46352 4981
rect 46963 4978 46975 4981
rect 47009 4978 47021 5012
rect 46963 4972 47021 4978
rect 47632 4969 47638 5021
rect 47690 5009 47696 5021
rect 47731 5012 47789 5018
rect 47731 5009 47743 5012
rect 47690 4981 47743 5009
rect 47690 4969 47696 4981
rect 47731 4978 47743 4981
rect 47777 4978 47789 5012
rect 49360 5009 49366 5021
rect 49321 4981 49366 5009
rect 47731 4972 47789 4978
rect 49360 4969 49366 4981
rect 49418 4969 49424 5021
rect 50416 5009 50422 5021
rect 50377 4981 50422 5009
rect 50416 4969 50422 4981
rect 50474 4969 50480 5021
rect 50896 4969 50902 5021
rect 50954 5009 50960 5021
rect 51091 5012 51149 5018
rect 51091 5009 51103 5012
rect 50954 4981 51103 5009
rect 50954 4969 50960 4981
rect 51091 4978 51103 4981
rect 51137 4978 51149 5012
rect 51856 5009 51862 5021
rect 51817 4981 51862 5009
rect 51091 4972 51149 4978
rect 51856 4969 51862 4981
rect 51914 4969 51920 5021
rect 52240 4969 52246 5021
rect 52298 5009 52304 5021
rect 52627 5012 52685 5018
rect 52627 5009 52639 5012
rect 52298 4981 52639 5009
rect 52298 4969 52304 4981
rect 52627 4978 52639 4981
rect 52673 4978 52685 5012
rect 52627 4972 52685 4978
rect 53296 4969 53302 5021
rect 53354 5009 53360 5021
rect 54451 5012 54509 5018
rect 54451 5009 54463 5012
rect 53354 4981 54463 5009
rect 53354 4969 53360 4981
rect 54451 4978 54463 4981
rect 54497 4978 54509 5012
rect 54451 4972 54509 4978
rect 55603 5012 55661 5018
rect 55603 4978 55615 5012
rect 55649 4978 55661 5012
rect 55603 4972 55661 4978
rect 56371 5012 56429 5018
rect 56371 4978 56383 5012
rect 56417 4978 56429 5012
rect 57040 5009 57046 5021
rect 57001 4981 57046 5009
rect 56371 4972 56429 4978
rect 34634 4907 35678 4935
rect 34634 4895 34640 4907
rect 7942 4889 7994 4895
rect 8368 4861 8374 4873
rect 8256 4833 8374 4861
rect 8368 4821 8374 4833
rect 8426 4821 8432 4873
rect 55618 4861 55646 4972
rect 56386 4935 56414 4972
rect 57040 4969 57046 4981
rect 57098 4969 57104 5021
rect 57808 4935 57814 4947
rect 56386 4907 57814 4935
rect 57808 4895 57814 4907
rect 57866 4895 57872 4947
rect 59248 4861 59254 4873
rect 55618 4833 59254 4861
rect 59248 4821 59254 4833
rect 59306 4821 59312 4873
rect 1152 4688 58848 4710
rect 1152 4636 19654 4688
rect 19706 4636 19718 4688
rect 19770 4636 19782 4688
rect 19834 4636 19846 4688
rect 19898 4636 50374 4688
rect 50426 4636 50438 4688
rect 50490 4636 50502 4688
rect 50554 4636 50566 4688
rect 50618 4636 58848 4688
rect 1152 4614 58848 4636
rect 7888 4525 7894 4577
rect 7946 4565 7952 4577
rect 9232 4565 9238 4577
rect 7946 4537 9238 4565
rect 7946 4525 7952 4537
rect 9232 4525 9238 4537
rect 9290 4525 9296 4577
rect 11152 4525 11158 4577
rect 11210 4565 11216 4577
rect 15763 4568 15821 4574
rect 15763 4565 15775 4568
rect 11210 4537 15775 4565
rect 11210 4525 11216 4537
rect 15763 4534 15775 4537
rect 15809 4534 15821 4568
rect 15763 4528 15821 4534
rect 12112 4451 12118 4503
rect 12170 4491 12176 4503
rect 16531 4494 16589 4500
rect 16531 4491 16543 4494
rect 12170 4463 16543 4491
rect 12170 4451 12176 4463
rect 16531 4460 16543 4463
rect 16577 4460 16589 4494
rect 16531 4454 16589 4460
rect 33904 4451 33910 4503
rect 33962 4491 33968 4503
rect 35344 4491 35350 4503
rect 33962 4463 35350 4491
rect 33962 4451 33968 4463
rect 35344 4451 35350 4463
rect 35402 4451 35408 4503
rect 784 4377 790 4429
rect 842 4417 848 4429
rect 842 4389 2366 4417
rect 842 4377 848 4389
rect 1168 4303 1174 4355
rect 1226 4343 1232 4355
rect 2338 4352 2366 4389
rect 11056 4377 11062 4429
rect 11114 4417 11120 4429
rect 15088 4417 15094 4429
rect 11114 4389 15094 4417
rect 11114 4377 11120 4389
rect 15088 4377 15094 4389
rect 15146 4377 15152 4429
rect 1555 4346 1613 4352
rect 1555 4343 1567 4346
rect 1226 4315 1567 4343
rect 1226 4303 1232 4315
rect 1555 4312 1567 4315
rect 1601 4312 1613 4346
rect 1555 4306 1613 4312
rect 2323 4346 2381 4352
rect 2323 4312 2335 4346
rect 2369 4312 2381 4346
rect 3091 4346 3149 4352
rect 3091 4343 3103 4346
rect 2323 4306 2381 4312
rect 2866 4315 3103 4343
rect 1360 4229 1366 4281
rect 1418 4269 1424 4281
rect 2866 4269 2894 4315
rect 3091 4312 3103 4315
rect 3137 4312 3149 4346
rect 3091 4306 3149 4312
rect 4339 4346 4397 4352
rect 4339 4312 4351 4346
rect 4385 4312 4397 4346
rect 4339 4306 4397 4312
rect 1418 4241 2894 4269
rect 1418 4229 1424 4241
rect 3760 4229 3766 4281
rect 3818 4269 3824 4281
rect 4354 4269 4382 4306
rect 4720 4303 4726 4355
rect 4778 4343 4784 4355
rect 5107 4346 5165 4352
rect 5107 4343 5119 4346
rect 4778 4315 5119 4343
rect 4778 4303 4784 4315
rect 5107 4312 5119 4315
rect 5153 4312 5165 4346
rect 5875 4346 5933 4352
rect 5875 4343 5887 4346
rect 5107 4306 5165 4312
rect 5602 4315 5887 4343
rect 3818 4241 4382 4269
rect 3818 4229 3824 4241
rect 5008 4229 5014 4281
rect 5066 4269 5072 4281
rect 5602 4269 5630 4315
rect 5875 4312 5887 4315
rect 5921 4312 5933 4346
rect 5875 4306 5933 4312
rect 6643 4346 6701 4352
rect 6643 4312 6655 4346
rect 6689 4312 6701 4346
rect 7408 4343 7414 4355
rect 7369 4315 7414 4343
rect 6643 4306 6701 4312
rect 5066 4241 5630 4269
rect 5066 4229 5072 4241
rect 5680 4229 5686 4281
rect 5738 4269 5744 4281
rect 6658 4269 6686 4306
rect 7408 4303 7414 4315
rect 7466 4303 7472 4355
rect 8179 4346 8237 4352
rect 8179 4312 8191 4346
rect 8225 4312 8237 4346
rect 9616 4343 9622 4355
rect 9577 4315 9622 4343
rect 8179 4306 8237 4312
rect 5738 4241 6686 4269
rect 5738 4229 5744 4241
rect 3472 4155 3478 4207
rect 3530 4195 3536 4207
rect 4912 4195 4918 4207
rect 3530 4167 4918 4195
rect 3530 4155 3536 4167
rect 4912 4155 4918 4167
rect 4970 4155 4976 4207
rect 6448 4155 6454 4207
rect 6506 4195 6512 4207
rect 8194 4195 8222 4306
rect 9616 4303 9622 4315
rect 9674 4303 9680 4355
rect 10384 4343 10390 4355
rect 10345 4315 10390 4343
rect 10384 4303 10390 4315
rect 10442 4303 10448 4355
rect 10768 4303 10774 4355
rect 10826 4343 10832 4355
rect 11155 4346 11213 4352
rect 11155 4343 11167 4346
rect 10826 4315 11167 4343
rect 10826 4303 10832 4315
rect 11155 4312 11167 4315
rect 11201 4312 11213 4346
rect 11923 4346 11981 4352
rect 11923 4343 11935 4346
rect 11155 4306 11213 4312
rect 11266 4315 11935 4343
rect 9808 4229 9814 4281
rect 9866 4269 9872 4281
rect 10192 4269 10198 4281
rect 9866 4241 10198 4269
rect 9866 4229 9872 4241
rect 10192 4229 10198 4241
rect 10250 4229 10256 4281
rect 6506 4167 8222 4195
rect 6506 4155 6512 4167
rect 11152 4155 11158 4207
rect 11210 4195 11216 4207
rect 11266 4195 11294 4315
rect 11923 4312 11935 4315
rect 11969 4312 11981 4346
rect 11923 4306 11981 4312
rect 12691 4346 12749 4352
rect 12691 4312 12703 4346
rect 12737 4312 12749 4346
rect 13552 4343 13558 4355
rect 13513 4315 13558 4343
rect 12691 4306 12749 4312
rect 11440 4229 11446 4281
rect 11498 4269 11504 4281
rect 12706 4269 12734 4306
rect 13552 4303 13558 4315
rect 13610 4303 13616 4355
rect 15472 4343 15478 4355
rect 15433 4315 15478 4343
rect 15472 4303 15478 4315
rect 15530 4303 15536 4355
rect 15952 4303 15958 4355
rect 16010 4343 16016 4355
rect 16243 4346 16301 4352
rect 16243 4343 16255 4346
rect 16010 4315 16255 4343
rect 16010 4303 16016 4315
rect 16243 4312 16255 4315
rect 16289 4312 16301 4346
rect 16243 4306 16301 4312
rect 17011 4346 17069 4352
rect 17011 4312 17023 4346
rect 17057 4312 17069 4346
rect 17779 4346 17837 4352
rect 17779 4343 17791 4346
rect 17011 4306 17069 4312
rect 17266 4315 17791 4343
rect 11498 4241 12734 4269
rect 11498 4229 11504 4241
rect 14896 4229 14902 4281
rect 14954 4269 14960 4281
rect 16528 4269 16534 4281
rect 14954 4241 16534 4269
rect 14954 4229 14960 4241
rect 16528 4229 16534 4241
rect 16586 4229 16592 4281
rect 11210 4167 11294 4195
rect 11210 4155 11216 4167
rect 16240 4155 16246 4207
rect 16298 4195 16304 4207
rect 17026 4195 17054 4306
rect 17266 4269 17294 4315
rect 17779 4312 17791 4315
rect 17825 4312 17837 4346
rect 17779 4306 17837 4312
rect 18547 4346 18605 4352
rect 18547 4312 18559 4346
rect 18593 4312 18605 4346
rect 20272 4343 20278 4355
rect 20233 4315 20278 4343
rect 18547 4306 18605 4312
rect 16298 4167 17054 4195
rect 17122 4241 17294 4269
rect 16298 4155 16304 4167
rect 16912 4081 16918 4133
rect 16970 4121 16976 4133
rect 17122 4121 17150 4241
rect 17680 4229 17686 4281
rect 17738 4269 17744 4281
rect 18562 4269 18590 4306
rect 20272 4303 20278 4315
rect 20330 4303 20336 4355
rect 21040 4343 21046 4355
rect 21001 4315 21046 4343
rect 21040 4303 21046 4315
rect 21098 4303 21104 4355
rect 21808 4343 21814 4355
rect 21769 4315 21814 4343
rect 21808 4303 21814 4315
rect 21866 4303 21872 4355
rect 23248 4343 23254 4355
rect 23209 4315 23254 4343
rect 23248 4303 23254 4315
rect 23306 4303 23312 4355
rect 24019 4346 24077 4352
rect 24019 4312 24031 4346
rect 24065 4312 24077 4346
rect 25456 4343 25462 4355
rect 25417 4315 25462 4343
rect 24019 4306 24077 4312
rect 17738 4241 18590 4269
rect 17738 4229 17744 4241
rect 22000 4229 22006 4281
rect 22058 4269 22064 4281
rect 24034 4269 24062 4306
rect 25456 4303 25462 4315
rect 25514 4303 25520 4355
rect 26128 4303 26134 4355
rect 26186 4343 26192 4355
rect 26227 4346 26285 4352
rect 26227 4343 26239 4346
rect 26186 4315 26239 4343
rect 26186 4303 26192 4315
rect 26227 4312 26239 4315
rect 26273 4312 26285 4346
rect 26227 4306 26285 4312
rect 26512 4303 26518 4355
rect 26570 4343 26576 4355
rect 26995 4346 27053 4352
rect 26995 4343 27007 4346
rect 26570 4315 27007 4343
rect 26570 4303 26576 4315
rect 26995 4312 27007 4315
rect 27041 4312 27053 4346
rect 28336 4343 28342 4355
rect 28297 4315 28342 4343
rect 26995 4306 27053 4312
rect 28336 4303 28342 4315
rect 28394 4303 28400 4355
rect 29104 4343 29110 4355
rect 29065 4315 29110 4343
rect 29104 4303 29110 4315
rect 29162 4303 29168 4355
rect 30928 4343 30934 4355
rect 30889 4315 30934 4343
rect 30928 4303 30934 4315
rect 30986 4303 30992 4355
rect 31696 4343 31702 4355
rect 31657 4315 31702 4343
rect 31696 4303 31702 4315
rect 31754 4303 31760 4355
rect 32752 4343 32758 4355
rect 32713 4315 32758 4343
rect 32752 4303 32758 4315
rect 32810 4303 32816 4355
rect 33904 4343 33910 4355
rect 33865 4315 33910 4343
rect 33904 4303 33910 4315
rect 33962 4303 33968 4355
rect 34576 4303 34582 4355
rect 34634 4343 34640 4355
rect 34675 4346 34733 4352
rect 34675 4343 34687 4346
rect 34634 4315 34687 4343
rect 34634 4303 34640 4315
rect 34675 4312 34687 4315
rect 34721 4312 34733 4346
rect 36019 4346 36077 4352
rect 36019 4343 36031 4346
rect 34675 4306 34733 4312
rect 34786 4315 36031 4343
rect 22058 4241 24062 4269
rect 22058 4229 22064 4241
rect 34192 4229 34198 4281
rect 34250 4269 34256 4281
rect 34786 4269 34814 4315
rect 36019 4312 36031 4315
rect 36065 4312 36077 4346
rect 36784 4343 36790 4355
rect 36745 4315 36790 4343
rect 36019 4306 36077 4312
rect 36784 4303 36790 4315
rect 36842 4303 36848 4355
rect 37555 4346 37613 4352
rect 37555 4343 37567 4346
rect 37426 4315 37567 4343
rect 34250 4241 34814 4269
rect 34250 4229 34256 4241
rect 37168 4229 37174 4281
rect 37226 4269 37232 4281
rect 37426 4269 37454 4315
rect 37555 4312 37567 4315
rect 37601 4312 37613 4346
rect 38992 4343 38998 4355
rect 38953 4315 38998 4343
rect 37555 4306 37613 4312
rect 38992 4303 38998 4315
rect 39050 4303 39056 4355
rect 39760 4343 39766 4355
rect 39721 4315 39766 4343
rect 39760 4303 39766 4315
rect 39818 4303 39824 4355
rect 41968 4343 41974 4355
rect 41929 4315 41974 4343
rect 41968 4303 41974 4315
rect 42026 4303 42032 4355
rect 42352 4303 42358 4355
rect 42410 4343 42416 4355
rect 42739 4346 42797 4352
rect 42739 4343 42751 4346
rect 42410 4315 42751 4343
rect 42410 4303 42416 4315
rect 42739 4312 42751 4315
rect 42785 4312 42797 4346
rect 42739 4306 42797 4312
rect 43408 4303 43414 4355
rect 43466 4343 43472 4355
rect 43507 4346 43565 4352
rect 43507 4343 43519 4346
rect 43466 4315 43519 4343
rect 43466 4303 43472 4315
rect 43507 4312 43519 4315
rect 43553 4312 43565 4346
rect 44944 4343 44950 4355
rect 44905 4315 44950 4343
rect 43507 4306 43565 4312
rect 44944 4303 44950 4315
rect 45002 4303 45008 4355
rect 46768 4343 46774 4355
rect 46729 4315 46774 4343
rect 46768 4303 46774 4315
rect 46826 4303 46832 4355
rect 47539 4346 47597 4352
rect 47539 4312 47551 4346
rect 47585 4312 47597 4346
rect 47539 4306 47597 4312
rect 37226 4241 37454 4269
rect 37226 4229 37232 4241
rect 43792 4229 43798 4281
rect 43850 4269 43856 4281
rect 44467 4272 44525 4278
rect 44467 4269 44479 4272
rect 43850 4241 44479 4269
rect 43850 4229 43856 4241
rect 44467 4238 44479 4241
rect 44513 4238 44525 4272
rect 44467 4232 44525 4238
rect 47440 4229 47446 4281
rect 47498 4269 47504 4281
rect 47554 4269 47582 4306
rect 47824 4303 47830 4355
rect 47882 4343 47888 4355
rect 48307 4346 48365 4352
rect 48307 4343 48319 4346
rect 47882 4315 48319 4343
rect 47882 4303 47888 4315
rect 48307 4312 48319 4315
rect 48353 4312 48365 4346
rect 48307 4306 48365 4312
rect 49075 4346 49133 4352
rect 49075 4312 49087 4346
rect 49121 4312 49133 4346
rect 49840 4343 49846 4355
rect 49801 4315 49846 4343
rect 49075 4306 49133 4312
rect 47498 4241 47582 4269
rect 47498 4229 47504 4241
rect 48592 4229 48598 4281
rect 48650 4269 48656 4281
rect 49090 4269 49118 4306
rect 49840 4303 49846 4315
rect 49898 4303 49904 4355
rect 50611 4346 50669 4352
rect 50611 4312 50623 4346
rect 50657 4312 50669 4346
rect 50611 4306 50669 4312
rect 51859 4346 51917 4352
rect 51859 4312 51871 4346
rect 51905 4312 51917 4346
rect 52624 4343 52630 4355
rect 52585 4315 52630 4343
rect 51859 4306 51917 4312
rect 48650 4241 49118 4269
rect 48650 4229 48656 4241
rect 49936 4229 49942 4281
rect 49994 4269 50000 4281
rect 50626 4269 50654 4306
rect 49994 4241 50654 4269
rect 49994 4229 50000 4241
rect 50992 4229 50998 4281
rect 51050 4269 51056 4281
rect 51874 4269 51902 4306
rect 52624 4303 52630 4315
rect 52682 4303 52688 4355
rect 53395 4346 53453 4352
rect 53395 4312 53407 4346
rect 53441 4312 53453 4346
rect 53395 4306 53453 4312
rect 51050 4241 51902 4269
rect 51050 4229 51056 4241
rect 53008 4229 53014 4281
rect 53066 4269 53072 4281
rect 53410 4269 53438 4306
rect 54064 4303 54070 4355
rect 54122 4343 54128 4355
rect 54163 4346 54221 4352
rect 54163 4343 54175 4346
rect 54122 4315 54175 4343
rect 54122 4303 54128 4315
rect 54163 4312 54175 4315
rect 54209 4312 54221 4346
rect 55600 4343 55606 4355
rect 55561 4315 55606 4343
rect 54163 4306 54221 4312
rect 55600 4303 55606 4315
rect 55658 4303 55664 4355
rect 56656 4303 56662 4355
rect 56714 4343 56720 4355
rect 57139 4346 57197 4352
rect 57139 4343 57151 4346
rect 56714 4315 57151 4343
rect 56714 4303 56720 4315
rect 57139 4312 57151 4315
rect 57185 4312 57197 4346
rect 57139 4306 57197 4312
rect 53066 4241 53438 4269
rect 53066 4229 53072 4241
rect 57328 4229 57334 4281
rect 57386 4269 57392 4281
rect 59152 4269 59158 4281
rect 57386 4241 59158 4269
rect 57386 4229 57392 4241
rect 59152 4229 59158 4241
rect 59210 4229 59216 4281
rect 27472 4155 27478 4207
rect 27530 4195 27536 4207
rect 29008 4195 29014 4207
rect 27530 4167 29014 4195
rect 27530 4155 27536 4167
rect 29008 4155 29014 4167
rect 29066 4155 29072 4207
rect 38512 4155 38518 4207
rect 38570 4195 38576 4207
rect 40144 4195 40150 4207
rect 38570 4167 40150 4195
rect 38570 4155 38576 4167
rect 40144 4155 40150 4167
rect 40202 4155 40208 4207
rect 55216 4155 55222 4207
rect 55274 4195 55280 4207
rect 57904 4195 57910 4207
rect 55274 4167 57910 4195
rect 55274 4155 55280 4167
rect 57904 4155 57910 4167
rect 57962 4155 57968 4207
rect 16970 4093 17150 4121
rect 16970 4081 16976 4093
rect 17200 4081 17206 4133
rect 17258 4121 17264 4133
rect 41491 4124 41549 4130
rect 41491 4121 41503 4124
rect 17258 4093 41503 4121
rect 17258 4081 17264 4093
rect 41491 4090 41503 4093
rect 41537 4090 41549 4124
rect 41491 4084 41549 4090
rect 1152 4022 58848 4044
rect 1152 3970 4294 4022
rect 4346 3970 4358 4022
rect 4410 3970 4422 4022
rect 4474 3970 4486 4022
rect 4538 3970 35014 4022
rect 35066 3970 35078 4022
rect 35130 3970 35142 4022
rect 35194 3970 35206 4022
rect 35258 3970 58848 4022
rect 1152 3948 58848 3970
rect 1936 3859 1942 3911
rect 1994 3899 2000 3911
rect 2992 3899 2998 3911
rect 1994 3871 2998 3899
rect 1994 3859 2000 3871
rect 2992 3859 2998 3871
rect 3050 3859 3056 3911
rect 9040 3859 9046 3911
rect 9098 3899 9104 3911
rect 10576 3899 10582 3911
rect 9098 3871 10582 3899
rect 9098 3859 9104 3871
rect 10576 3859 10582 3871
rect 10634 3859 10640 3911
rect 12304 3859 12310 3911
rect 12362 3899 12368 3911
rect 12403 3902 12461 3908
rect 12403 3899 12415 3902
rect 12362 3871 12415 3899
rect 12362 3859 12368 3871
rect 12403 3868 12415 3871
rect 12449 3868 12461 3902
rect 12403 3862 12461 3868
rect 13168 3859 13174 3911
rect 13226 3899 13232 3911
rect 13939 3902 13997 3908
rect 13939 3899 13951 3902
rect 13226 3871 13951 3899
rect 13226 3859 13232 3871
rect 13939 3868 13951 3871
rect 13985 3868 13997 3902
rect 13939 3862 13997 3868
rect 14128 3859 14134 3911
rect 14186 3899 14192 3911
rect 15475 3902 15533 3908
rect 15475 3899 15487 3902
rect 14186 3871 15487 3899
rect 14186 3859 14192 3871
rect 15475 3868 15487 3871
rect 15521 3868 15533 3902
rect 15475 3862 15533 3868
rect 15760 3859 15766 3911
rect 15818 3899 15824 3911
rect 17200 3899 17206 3911
rect 15818 3871 17206 3899
rect 15818 3859 15824 3871
rect 17200 3859 17206 3871
rect 17258 3859 17264 3911
rect 17776 3859 17782 3911
rect 17834 3899 17840 3911
rect 18547 3902 18605 3908
rect 18547 3899 18559 3902
rect 17834 3871 18559 3899
rect 17834 3859 17840 3871
rect 18547 3868 18559 3871
rect 18593 3868 18605 3902
rect 18547 3862 18605 3868
rect 21328 3859 21334 3911
rect 21386 3899 21392 3911
rect 22768 3899 22774 3911
rect 21386 3871 22774 3899
rect 21386 3859 21392 3871
rect 22768 3859 22774 3871
rect 22826 3859 22832 3911
rect 28528 3859 28534 3911
rect 28586 3899 28592 3911
rect 29488 3899 29494 3911
rect 28586 3871 29494 3899
rect 28586 3859 28592 3871
rect 29488 3859 29494 3871
rect 29546 3859 29552 3911
rect 32560 3859 32566 3911
rect 32618 3899 32624 3911
rect 34288 3899 34294 3911
rect 32618 3871 34294 3899
rect 32618 3859 32624 3871
rect 34288 3859 34294 3871
rect 34346 3859 34352 3911
rect 38704 3899 38710 3911
rect 37426 3871 38710 3899
rect 496 3785 502 3837
rect 554 3825 560 3837
rect 1648 3825 1654 3837
rect 554 3797 1654 3825
rect 554 3785 560 3797
rect 1648 3785 1654 3797
rect 1706 3785 1712 3837
rect 2320 3785 2326 3837
rect 2378 3825 2384 3837
rect 3088 3825 3094 3837
rect 2378 3797 3094 3825
rect 2378 3785 2384 3797
rect 3088 3785 3094 3797
rect 3146 3785 3152 3837
rect 8272 3785 8278 3837
rect 8330 3825 8336 3837
rect 10000 3825 10006 3837
rect 8330 3797 10006 3825
rect 8330 3785 8336 3797
rect 10000 3785 10006 3797
rect 10058 3785 10064 3837
rect 16528 3785 16534 3837
rect 16586 3825 16592 3837
rect 17296 3825 17302 3837
rect 16586 3797 17302 3825
rect 16586 3785 16592 3797
rect 17296 3785 17302 3797
rect 17354 3785 17360 3837
rect 19408 3785 19414 3837
rect 19466 3825 19472 3837
rect 20656 3825 20662 3837
rect 19466 3797 20662 3825
rect 19466 3785 19472 3797
rect 20656 3785 20662 3797
rect 20714 3785 20720 3837
rect 24208 3785 24214 3837
rect 24266 3825 24272 3837
rect 25840 3825 25846 3837
rect 24266 3797 25846 3825
rect 24266 3785 24272 3797
rect 25840 3785 25846 3797
rect 25898 3785 25904 3837
rect 26416 3785 26422 3837
rect 26474 3825 26480 3837
rect 28048 3825 28054 3837
rect 26474 3797 28054 3825
rect 26474 3785 26480 3797
rect 28048 3785 28054 3797
rect 28106 3785 28112 3837
rect 29008 3785 29014 3837
rect 29066 3825 29072 3837
rect 30352 3825 30358 3837
rect 29066 3797 30358 3825
rect 29066 3785 29072 3797
rect 30352 3785 30358 3797
rect 30410 3785 30416 3837
rect 33424 3785 33430 3837
rect 33482 3825 33488 3837
rect 34864 3825 34870 3837
rect 33482 3797 34870 3825
rect 33482 3785 33488 3797
rect 34864 3785 34870 3797
rect 34922 3785 34928 3837
rect 976 3711 982 3763
rect 1034 3751 1040 3763
rect 2416 3751 2422 3763
rect 1034 3723 2422 3751
rect 1034 3711 1040 3723
rect 2416 3711 2422 3723
rect 2474 3711 2480 3763
rect 2992 3711 2998 3763
rect 3050 3751 3056 3763
rect 3280 3751 3286 3763
rect 3050 3723 3286 3751
rect 3050 3711 3056 3723
rect 3280 3711 3286 3723
rect 3338 3711 3344 3763
rect 3376 3711 3382 3763
rect 3434 3751 3440 3763
rect 3434 3723 4670 3751
rect 3434 3711 3440 3723
rect 592 3637 598 3689
rect 650 3677 656 3689
rect 1456 3677 1462 3689
rect 650 3649 1462 3677
rect 650 3637 656 3649
rect 1456 3637 1462 3649
rect 1514 3637 1520 3689
rect 1555 3680 1613 3686
rect 1555 3646 1567 3680
rect 1601 3646 1613 3680
rect 1555 3640 1613 3646
rect 112 3563 118 3615
rect 170 3603 176 3615
rect 1570 3603 1598 3640
rect 1648 3637 1654 3689
rect 1706 3677 1712 3689
rect 2323 3680 2381 3686
rect 2323 3677 2335 3680
rect 1706 3649 2335 3677
rect 1706 3637 1712 3649
rect 2323 3646 2335 3649
rect 2369 3646 2381 3680
rect 2323 3640 2381 3646
rect 2704 3637 2710 3689
rect 2762 3677 2768 3689
rect 3091 3680 3149 3686
rect 3091 3677 3103 3680
rect 2762 3649 3103 3677
rect 2762 3637 2768 3649
rect 3091 3646 3103 3649
rect 3137 3646 3149 3680
rect 3091 3640 3149 3646
rect 3568 3637 3574 3689
rect 3626 3677 3632 3689
rect 4642 3686 4670 3723
rect 8752 3711 8758 3763
rect 8810 3751 8816 3763
rect 37426 3751 37454 3871
rect 38704 3859 38710 3871
rect 38762 3859 38768 3911
rect 40048 3859 40054 3911
rect 40106 3899 40112 3911
rect 41680 3899 41686 3911
rect 40106 3871 41686 3899
rect 40106 3859 40112 3871
rect 41680 3859 41686 3871
rect 41738 3859 41744 3911
rect 37840 3785 37846 3837
rect 37898 3825 37904 3837
rect 39376 3825 39382 3837
rect 37898 3797 39382 3825
rect 37898 3785 37904 3797
rect 39376 3785 39382 3797
rect 39434 3785 39440 3837
rect 49168 3785 49174 3837
rect 49226 3825 49232 3837
rect 50704 3825 50710 3837
rect 49226 3797 50710 3825
rect 49226 3785 49232 3797
rect 50704 3785 50710 3797
rect 50762 3785 50768 3837
rect 8810 3723 37454 3751
rect 8810 3711 8816 3723
rect 44560 3711 44566 3763
rect 44618 3751 44624 3763
rect 44618 3723 45470 3751
rect 44618 3711 44624 3723
rect 3859 3680 3917 3686
rect 3859 3677 3871 3680
rect 3626 3649 3871 3677
rect 3626 3637 3632 3649
rect 3859 3646 3871 3649
rect 3905 3646 3917 3680
rect 3859 3640 3917 3646
rect 4627 3680 4685 3686
rect 4627 3646 4639 3680
rect 4673 3646 4685 3680
rect 5584 3677 5590 3689
rect 5545 3649 5590 3677
rect 4627 3640 4685 3646
rect 5584 3637 5590 3649
rect 5642 3637 5648 3689
rect 6352 3637 6358 3689
rect 6410 3677 6416 3689
rect 6931 3680 6989 3686
rect 6931 3677 6943 3680
rect 6410 3649 6943 3677
rect 6410 3637 6416 3649
rect 6931 3646 6943 3649
rect 6977 3646 6989 3680
rect 6931 3640 6989 3646
rect 7024 3637 7030 3689
rect 7082 3677 7088 3689
rect 7699 3680 7757 3686
rect 7699 3677 7711 3680
rect 7082 3649 7711 3677
rect 7082 3637 7088 3649
rect 7699 3646 7711 3649
rect 7745 3646 7757 3680
rect 7699 3640 7757 3646
rect 7792 3637 7798 3689
rect 7850 3677 7856 3689
rect 8467 3680 8525 3686
rect 8467 3677 8479 3680
rect 7850 3649 8479 3677
rect 7850 3637 7856 3649
rect 8467 3646 8479 3649
rect 8513 3646 8525 3680
rect 8467 3640 8525 3646
rect 8560 3637 8566 3689
rect 8618 3677 8624 3689
rect 9235 3680 9293 3686
rect 9235 3677 9247 3680
rect 8618 3649 9247 3677
rect 8618 3637 8624 3649
rect 9235 3646 9247 3649
rect 9281 3646 9293 3680
rect 9235 3640 9293 3646
rect 9328 3637 9334 3689
rect 9386 3677 9392 3689
rect 10003 3680 10061 3686
rect 10003 3677 10015 3680
rect 9386 3649 10015 3677
rect 9386 3637 9392 3649
rect 10003 3646 10015 3649
rect 10049 3646 10061 3680
rect 10003 3640 10061 3646
rect 10771 3680 10829 3686
rect 10771 3646 10783 3680
rect 10817 3646 10829 3680
rect 10771 3640 10829 3646
rect 12979 3680 13037 3686
rect 12979 3646 12991 3680
rect 13025 3677 13037 3680
rect 13168 3677 13174 3689
rect 13025 3649 13174 3677
rect 13025 3646 13037 3649
rect 12979 3640 13037 3646
rect 5200 3603 5206 3615
rect 170 3575 1598 3603
rect 2866 3575 5206 3603
rect 170 3563 176 3575
rect 1456 3489 1462 3541
rect 1514 3529 1520 3541
rect 2128 3529 2134 3541
rect 1514 3501 2134 3529
rect 1514 3489 1520 3501
rect 2128 3489 2134 3501
rect 2186 3489 2192 3541
rect 2416 3415 2422 3467
rect 2474 3455 2480 3467
rect 2866 3455 2894 3575
rect 5200 3563 5206 3575
rect 5258 3563 5264 3615
rect 10000 3489 10006 3541
rect 10058 3529 10064 3541
rect 10786 3529 10814 3640
rect 13168 3637 13174 3649
rect 13226 3637 13232 3689
rect 13648 3677 13654 3689
rect 13609 3649 13654 3677
rect 13648 3637 13654 3649
rect 13706 3637 13712 3689
rect 14128 3637 14134 3689
rect 14186 3677 14192 3689
rect 14419 3680 14477 3686
rect 14419 3677 14431 3680
rect 14186 3649 14431 3677
rect 14186 3637 14192 3649
rect 14419 3646 14431 3649
rect 14465 3646 14477 3680
rect 14419 3640 14477 3646
rect 14800 3637 14806 3689
rect 14858 3677 14864 3689
rect 15187 3680 15245 3686
rect 15187 3677 15199 3680
rect 14858 3649 15199 3677
rect 14858 3637 14864 3649
rect 15187 3646 15199 3649
rect 15233 3646 15245 3680
rect 15187 3640 15245 3646
rect 15280 3637 15286 3689
rect 15338 3677 15344 3689
rect 15955 3680 16013 3686
rect 15955 3677 15967 3680
rect 15338 3649 15967 3677
rect 15338 3637 15344 3649
rect 15955 3646 15967 3649
rect 16001 3646 16013 3680
rect 15955 3640 16013 3646
rect 17392 3637 17398 3689
rect 17450 3677 17456 3689
rect 17491 3680 17549 3686
rect 17491 3677 17503 3680
rect 17450 3649 17503 3677
rect 17450 3637 17456 3649
rect 17491 3646 17503 3649
rect 17537 3646 17549 3680
rect 17491 3640 17549 3646
rect 18160 3637 18166 3689
rect 18218 3677 18224 3689
rect 18259 3680 18317 3686
rect 18259 3677 18271 3680
rect 18218 3649 18271 3677
rect 18218 3637 18224 3649
rect 18259 3646 18271 3649
rect 18305 3646 18317 3680
rect 18259 3640 18317 3646
rect 18448 3637 18454 3689
rect 18506 3677 18512 3689
rect 19027 3680 19085 3686
rect 19027 3677 19039 3680
rect 18506 3649 19039 3677
rect 18506 3637 18512 3649
rect 19027 3646 19039 3649
rect 19073 3646 19085 3680
rect 19027 3640 19085 3646
rect 19216 3637 19222 3689
rect 19274 3677 19280 3689
rect 19795 3680 19853 3686
rect 19795 3677 19807 3680
rect 19274 3649 19807 3677
rect 19274 3637 19280 3649
rect 19795 3646 19807 3649
rect 19841 3646 19853 3680
rect 19795 3640 19853 3646
rect 19984 3637 19990 3689
rect 20042 3677 20048 3689
rect 20563 3680 20621 3686
rect 20563 3677 20575 3680
rect 20042 3649 20575 3677
rect 20042 3637 20048 3649
rect 20563 3646 20575 3649
rect 20609 3646 20621 3680
rect 20563 3640 20621 3646
rect 20656 3637 20662 3689
rect 20714 3677 20720 3689
rect 21331 3680 21389 3686
rect 21331 3677 21343 3680
rect 20714 3649 21343 3677
rect 20714 3637 20720 3649
rect 21331 3646 21343 3649
rect 21377 3646 21389 3680
rect 21331 3640 21389 3646
rect 22096 3637 22102 3689
rect 22154 3677 22160 3689
rect 22771 3680 22829 3686
rect 22771 3677 22783 3680
rect 22154 3649 22783 3677
rect 22154 3637 22160 3649
rect 22771 3646 22783 3649
rect 22817 3646 22829 3680
rect 22771 3640 22829 3646
rect 22864 3637 22870 3689
rect 22922 3677 22928 3689
rect 23539 3680 23597 3686
rect 23539 3677 23551 3680
rect 22922 3649 23551 3677
rect 22922 3637 22928 3649
rect 23539 3646 23551 3649
rect 23585 3646 23597 3680
rect 23539 3640 23597 3646
rect 23632 3637 23638 3689
rect 23690 3677 23696 3689
rect 24307 3680 24365 3686
rect 24307 3677 24319 3680
rect 23690 3649 24319 3677
rect 23690 3637 23696 3649
rect 24307 3646 24319 3649
rect 24353 3646 24365 3680
rect 24307 3640 24365 3646
rect 24400 3637 24406 3689
rect 24458 3677 24464 3689
rect 25075 3680 25133 3686
rect 25075 3677 25087 3680
rect 24458 3649 25087 3677
rect 24458 3637 24464 3649
rect 25075 3646 25087 3649
rect 25121 3646 25133 3680
rect 25075 3640 25133 3646
rect 25843 3680 25901 3686
rect 25843 3646 25855 3680
rect 25889 3646 25901 3680
rect 25843 3640 25901 3646
rect 26611 3680 26669 3686
rect 26611 3646 26623 3680
rect 26657 3646 26669 3680
rect 26611 3640 26669 3646
rect 24688 3563 24694 3615
rect 24746 3603 24752 3615
rect 25858 3603 25886 3640
rect 24746 3575 25886 3603
rect 24746 3563 24752 3575
rect 10058 3501 10814 3529
rect 10058 3489 10064 3501
rect 17296 3489 17302 3541
rect 17354 3529 17360 3541
rect 17488 3529 17494 3541
rect 17354 3501 17494 3529
rect 17354 3489 17360 3501
rect 17488 3489 17494 3501
rect 17546 3489 17552 3541
rect 22576 3489 22582 3541
rect 22634 3529 22640 3541
rect 23344 3529 23350 3541
rect 22634 3501 23350 3529
rect 22634 3489 22640 3501
rect 23344 3489 23350 3501
rect 23402 3489 23408 3541
rect 25840 3489 25846 3541
rect 25898 3529 25904 3541
rect 26626 3529 26654 3640
rect 27280 3637 27286 3689
rect 27338 3677 27344 3689
rect 28051 3680 28109 3686
rect 28051 3677 28063 3680
rect 27338 3649 28063 3677
rect 27338 3637 27344 3649
rect 28051 3646 28063 3649
rect 28097 3646 28109 3680
rect 28051 3640 28109 3646
rect 28819 3680 28877 3686
rect 28819 3646 28831 3680
rect 28865 3646 28877 3680
rect 28819 3640 28877 3646
rect 29683 3680 29741 3686
rect 29683 3646 29695 3680
rect 29729 3646 29741 3680
rect 29683 3640 29741 3646
rect 25898 3501 26654 3529
rect 25898 3489 25904 3501
rect 28048 3489 28054 3541
rect 28106 3529 28112 3541
rect 28834 3529 28862 3640
rect 28106 3501 28862 3529
rect 28106 3489 28112 3501
rect 2474 3427 2894 3455
rect 2474 3415 2480 3427
rect 3280 3415 3286 3467
rect 3338 3455 3344 3467
rect 3952 3455 3958 3467
rect 3338 3427 3958 3455
rect 3338 3415 3344 3427
rect 3952 3415 3958 3427
rect 4010 3415 4016 3467
rect 12016 3415 12022 3467
rect 12074 3455 12080 3467
rect 13360 3455 13366 3467
rect 12074 3427 13366 3455
rect 12074 3415 12080 3427
rect 13360 3415 13366 3427
rect 13418 3415 13424 3467
rect 22960 3415 22966 3467
rect 23018 3455 23024 3467
rect 24016 3455 24022 3467
rect 23018 3427 24022 3455
rect 23018 3415 23024 3427
rect 24016 3415 24022 3427
rect 24074 3415 24080 3467
rect 28720 3415 28726 3467
rect 28778 3455 28784 3467
rect 29698 3455 29726 3640
rect 29872 3637 29878 3689
rect 29930 3677 29936 3689
rect 30355 3680 30413 3686
rect 30355 3677 30367 3680
rect 29930 3649 30367 3677
rect 29930 3637 29936 3649
rect 30355 3646 30367 3649
rect 30401 3646 30413 3680
rect 30355 3640 30413 3646
rect 30448 3637 30454 3689
rect 30506 3677 30512 3689
rect 31123 3680 31181 3686
rect 31123 3677 31135 3680
rect 30506 3649 31135 3677
rect 30506 3637 30512 3649
rect 31123 3646 31135 3649
rect 31169 3646 31181 3680
rect 31123 3640 31181 3646
rect 31312 3637 31318 3689
rect 31370 3677 31376 3689
rect 31891 3680 31949 3686
rect 31891 3677 31903 3680
rect 31370 3649 31903 3677
rect 31370 3637 31376 3649
rect 31891 3646 31903 3649
rect 31937 3646 31949 3680
rect 31891 3640 31949 3646
rect 32464 3637 32470 3689
rect 32522 3677 32528 3689
rect 33331 3680 33389 3686
rect 33331 3677 33343 3680
rect 32522 3649 33343 3677
rect 32522 3637 32528 3649
rect 33331 3646 33343 3649
rect 33377 3646 33389 3680
rect 33331 3640 33389 3646
rect 33520 3637 33526 3689
rect 33578 3677 33584 3689
rect 34099 3680 34157 3686
rect 34099 3677 34111 3680
rect 33578 3649 34111 3677
rect 33578 3637 33584 3649
rect 34099 3646 34111 3649
rect 34145 3646 34157 3680
rect 34099 3640 34157 3646
rect 34288 3637 34294 3689
rect 34346 3677 34352 3689
rect 34867 3680 34925 3686
rect 34867 3677 34879 3680
rect 34346 3649 34879 3677
rect 34346 3637 34352 3649
rect 34867 3646 34879 3649
rect 34913 3646 34925 3680
rect 34867 3640 34925 3646
rect 34960 3637 34966 3689
rect 35018 3677 35024 3689
rect 35635 3680 35693 3686
rect 35635 3677 35647 3680
rect 35018 3649 35647 3677
rect 35018 3637 35024 3649
rect 35635 3646 35647 3649
rect 35681 3646 35693 3680
rect 35635 3640 35693 3646
rect 35728 3637 35734 3689
rect 35786 3677 35792 3689
rect 36403 3680 36461 3686
rect 36403 3677 36415 3680
rect 35786 3649 36415 3677
rect 35786 3637 35792 3649
rect 36403 3646 36415 3649
rect 36449 3646 36461 3680
rect 36403 3640 36461 3646
rect 36496 3637 36502 3689
rect 36554 3677 36560 3689
rect 37171 3680 37229 3686
rect 37171 3677 37183 3680
rect 36554 3649 37183 3677
rect 36554 3637 36560 3649
rect 37171 3646 37183 3649
rect 37217 3646 37229 3680
rect 37171 3640 37229 3646
rect 37936 3637 37942 3689
rect 37994 3677 38000 3689
rect 38611 3680 38669 3686
rect 38611 3677 38623 3680
rect 37994 3649 38623 3677
rect 37994 3637 38000 3649
rect 38611 3646 38623 3649
rect 38657 3646 38669 3680
rect 38611 3640 38669 3646
rect 38704 3637 38710 3689
rect 38762 3677 38768 3689
rect 39379 3680 39437 3686
rect 39379 3677 39391 3680
rect 38762 3649 39391 3677
rect 38762 3637 38768 3649
rect 39379 3646 39391 3649
rect 39425 3646 39437 3680
rect 39379 3640 39437 3646
rect 40147 3680 40205 3686
rect 40147 3646 40159 3680
rect 40193 3646 40205 3680
rect 40147 3640 40205 3646
rect 40915 3680 40973 3686
rect 40915 3646 40927 3680
rect 40961 3646 40973 3680
rect 40915 3640 40973 3646
rect 40162 3603 40190 3640
rect 39394 3575 40190 3603
rect 39394 3541 39422 3575
rect 39376 3489 39382 3541
rect 39434 3489 39440 3541
rect 40144 3489 40150 3541
rect 40202 3529 40208 3541
rect 40930 3529 40958 3640
rect 41008 3637 41014 3689
rect 41066 3677 41072 3689
rect 41683 3680 41741 3686
rect 41683 3677 41695 3680
rect 41066 3649 41695 3677
rect 41066 3637 41072 3649
rect 41683 3646 41695 3649
rect 41729 3646 41741 3680
rect 41683 3640 41741 3646
rect 42451 3680 42509 3686
rect 42451 3646 42463 3680
rect 42497 3646 42509 3680
rect 42451 3640 42509 3646
rect 41584 3563 41590 3615
rect 41642 3603 41648 3615
rect 42466 3603 42494 3640
rect 42736 3637 42742 3689
rect 42794 3677 42800 3689
rect 45442 3686 45470 3723
rect 55888 3711 55894 3763
rect 55946 3751 55952 3763
rect 55946 3723 56798 3751
rect 55946 3711 55952 3723
rect 43891 3680 43949 3686
rect 43891 3677 43903 3680
rect 42794 3649 43903 3677
rect 42794 3637 42800 3649
rect 43891 3646 43903 3649
rect 43937 3646 43949 3680
rect 43891 3640 43949 3646
rect 44659 3680 44717 3686
rect 44659 3646 44671 3680
rect 44705 3646 44717 3680
rect 44659 3640 44717 3646
rect 45427 3680 45485 3686
rect 45427 3646 45439 3680
rect 45473 3646 45485 3680
rect 45427 3640 45485 3646
rect 46195 3680 46253 3686
rect 46195 3646 46207 3680
rect 46241 3646 46253 3680
rect 46195 3640 46253 3646
rect 46963 3680 47021 3686
rect 46963 3646 46975 3680
rect 47009 3646 47021 3680
rect 46963 3640 47021 3646
rect 41642 3575 42494 3603
rect 41642 3563 41648 3575
rect 43792 3563 43798 3615
rect 43850 3603 43856 3615
rect 44674 3603 44702 3640
rect 43850 3575 44702 3603
rect 43850 3563 43856 3575
rect 45232 3563 45238 3615
rect 45290 3603 45296 3615
rect 46210 3603 46238 3640
rect 45290 3575 46238 3603
rect 45290 3563 45296 3575
rect 40202 3501 40958 3529
rect 40202 3489 40208 3501
rect 41200 3489 41206 3541
rect 41258 3529 41264 3541
rect 41680 3529 41686 3541
rect 41258 3501 41686 3529
rect 41258 3489 41264 3501
rect 41680 3489 41686 3501
rect 41738 3489 41744 3541
rect 46000 3489 46006 3541
rect 46058 3529 46064 3541
rect 46978 3529 47006 3640
rect 47152 3637 47158 3689
rect 47210 3677 47216 3689
rect 47731 3680 47789 3686
rect 47731 3677 47743 3680
rect 47210 3649 47743 3677
rect 47210 3637 47216 3649
rect 47731 3646 47743 3649
rect 47777 3646 47789 3680
rect 47731 3640 47789 3646
rect 48208 3637 48214 3689
rect 48266 3677 48272 3689
rect 49171 3680 49229 3686
rect 49171 3677 49183 3680
rect 48266 3649 49183 3677
rect 48266 3637 48272 3649
rect 49171 3646 49183 3649
rect 49217 3646 49229 3680
rect 49171 3640 49229 3646
rect 50515 3680 50573 3686
rect 50515 3646 50527 3680
rect 50561 3677 50573 3680
rect 50704 3677 50710 3689
rect 50561 3649 50710 3677
rect 50561 3646 50573 3649
rect 50515 3640 50573 3646
rect 50704 3637 50710 3649
rect 50762 3637 50768 3689
rect 50800 3637 50806 3689
rect 50858 3677 50864 3689
rect 51187 3680 51245 3686
rect 51187 3677 51199 3680
rect 50858 3649 51199 3677
rect 50858 3637 50864 3649
rect 51187 3646 51199 3649
rect 51233 3646 51245 3680
rect 51187 3640 51245 3646
rect 51280 3637 51286 3689
rect 51338 3677 51344 3689
rect 51955 3680 52013 3686
rect 51955 3677 51967 3680
rect 51338 3649 51967 3677
rect 51338 3637 51344 3649
rect 51955 3646 51967 3649
rect 52001 3646 52013 3680
rect 51955 3640 52013 3646
rect 52048 3637 52054 3689
rect 52106 3677 52112 3689
rect 52723 3680 52781 3686
rect 52723 3677 52735 3680
rect 52106 3649 52735 3677
rect 52106 3637 52112 3649
rect 52723 3646 52735 3649
rect 52769 3646 52781 3680
rect 52723 3640 52781 3646
rect 53392 3637 53398 3689
rect 53450 3677 53456 3689
rect 56770 3686 56798 3723
rect 54451 3680 54509 3686
rect 54451 3677 54463 3680
rect 53450 3649 54463 3677
rect 53450 3637 53456 3649
rect 54451 3646 54463 3649
rect 54497 3646 54509 3680
rect 54451 3640 54509 3646
rect 55219 3680 55277 3686
rect 55219 3646 55231 3680
rect 55265 3646 55277 3680
rect 55219 3640 55277 3646
rect 55987 3680 56045 3686
rect 55987 3646 55999 3680
rect 56033 3646 56045 3680
rect 55987 3640 56045 3646
rect 56755 3680 56813 3686
rect 56755 3646 56767 3680
rect 56801 3646 56813 3680
rect 56755 3640 56813 3646
rect 57523 3680 57581 3686
rect 57523 3646 57535 3680
rect 57569 3646 57581 3680
rect 57523 3640 57581 3646
rect 46058 3501 47006 3529
rect 46058 3489 46064 3501
rect 52048 3489 52054 3541
rect 52106 3529 52112 3541
rect 52816 3529 52822 3541
rect 52106 3501 52822 3529
rect 52106 3489 52112 3501
rect 52816 3489 52822 3501
rect 52874 3489 52880 3541
rect 54448 3489 54454 3541
rect 54506 3529 54512 3541
rect 55234 3529 55262 3640
rect 54506 3501 55262 3529
rect 54506 3489 54512 3501
rect 28778 3427 29726 3455
rect 28778 3415 28784 3427
rect 33040 3415 33046 3467
rect 33098 3455 33104 3467
rect 33808 3455 33814 3467
rect 33098 3427 33814 3455
rect 33098 3415 33104 3427
rect 33808 3415 33814 3427
rect 33866 3415 33872 3467
rect 43504 3415 43510 3467
rect 43562 3455 43568 3467
rect 44752 3455 44758 3467
rect 43562 3427 44758 3455
rect 43562 3415 43568 3427
rect 44752 3415 44758 3427
rect 44810 3415 44816 3467
rect 55216 3415 55222 3467
rect 55274 3455 55280 3467
rect 56002 3455 56030 3640
rect 56272 3563 56278 3615
rect 56330 3603 56336 3615
rect 57538 3603 57566 3640
rect 58192 3637 58198 3689
rect 58250 3677 58256 3689
rect 59728 3677 59734 3689
rect 58250 3649 59734 3677
rect 58250 3637 58256 3649
rect 59728 3637 59734 3649
rect 59786 3637 59792 3689
rect 56330 3575 57566 3603
rect 56330 3563 56336 3575
rect 55274 3427 56030 3455
rect 55274 3415 55280 3427
rect 56368 3415 56374 3467
rect 56426 3455 56432 3467
rect 59440 3455 59446 3467
rect 56426 3427 59446 3455
rect 56426 3415 56432 3427
rect 59440 3415 59446 3427
rect 59498 3415 59504 3467
rect 1152 3356 58848 3378
rect 1152 3304 19654 3356
rect 19706 3304 19718 3356
rect 19770 3304 19782 3356
rect 19834 3304 19846 3356
rect 19898 3304 50374 3356
rect 50426 3304 50438 3356
rect 50490 3304 50502 3356
rect 50554 3304 50566 3356
rect 50618 3304 58848 3356
rect 1152 3282 58848 3304
rect 3952 3193 3958 3245
rect 4010 3233 4016 3245
rect 5104 3233 5110 3245
rect 4010 3205 5110 3233
rect 4010 3193 4016 3205
rect 5104 3193 5110 3205
rect 5162 3193 5168 3245
rect 13264 3233 13270 3245
rect 13225 3205 13270 3233
rect 13264 3193 13270 3205
rect 13322 3193 13328 3245
rect 14032 3233 14038 3245
rect 13993 3205 14038 3233
rect 14032 3193 14038 3205
rect 14090 3193 14096 3245
rect 15088 3193 15094 3245
rect 15146 3233 15152 3245
rect 15379 3236 15437 3242
rect 15379 3233 15391 3236
rect 15146 3205 15391 3233
rect 15146 3193 15152 3205
rect 15379 3202 15391 3205
rect 15425 3202 15437 3236
rect 16816 3233 16822 3245
rect 16777 3205 16822 3233
rect 15379 3196 15437 3202
rect 16816 3193 16822 3205
rect 16874 3193 16880 3245
rect 18064 3233 18070 3245
rect 18025 3205 18070 3233
rect 18064 3193 18070 3205
rect 18122 3193 18128 3245
rect 18832 3233 18838 3245
rect 18793 3205 18838 3233
rect 18832 3193 18838 3205
rect 18890 3193 18896 3245
rect 19696 3193 19702 3245
rect 19754 3233 19760 3245
rect 20368 3233 20374 3245
rect 19754 3205 20374 3233
rect 19754 3193 19760 3205
rect 20368 3193 20374 3205
rect 20426 3193 20432 3245
rect 23344 3193 23350 3245
rect 23402 3233 23408 3245
rect 23920 3233 23926 3245
rect 23402 3205 23926 3233
rect 23402 3193 23408 3205
rect 23920 3193 23926 3205
rect 23978 3193 23984 3245
rect 24976 3193 24982 3245
rect 25034 3233 25040 3245
rect 26608 3233 26614 3245
rect 25034 3205 26614 3233
rect 25034 3193 25040 3205
rect 26608 3193 26614 3205
rect 26666 3193 26672 3245
rect 28816 3193 28822 3245
rect 28874 3233 28880 3245
rect 29776 3233 29782 3245
rect 28874 3205 29782 3233
rect 28874 3193 28880 3205
rect 29776 3193 29782 3205
rect 29834 3193 29840 3245
rect 30448 3193 30454 3245
rect 30506 3233 30512 3245
rect 31888 3233 31894 3245
rect 30506 3205 31894 3233
rect 30506 3193 30512 3205
rect 31888 3193 31894 3205
rect 31946 3193 31952 3245
rect 32656 3193 32662 3245
rect 32714 3233 32720 3245
rect 34096 3233 34102 3245
rect 32714 3205 34102 3233
rect 32714 3193 32720 3205
rect 34096 3193 34102 3205
rect 34154 3193 34160 3245
rect 44752 3193 44758 3245
rect 44810 3233 44816 3245
rect 46192 3233 46198 3245
rect 44810 3205 46198 3233
rect 44810 3193 44816 3205
rect 46192 3193 46198 3205
rect 46250 3193 46256 3245
rect 48496 3193 48502 3245
rect 48554 3233 48560 3245
rect 49648 3233 49654 3245
rect 48554 3205 49654 3233
rect 48554 3193 48560 3205
rect 49648 3193 49654 3205
rect 49706 3193 49712 3245
rect 56848 3193 56854 3245
rect 56906 3233 56912 3245
rect 58000 3233 58006 3245
rect 56906 3205 58006 3233
rect 56906 3193 56912 3205
rect 58000 3193 58006 3205
rect 58058 3193 58064 3245
rect 208 3119 214 3171
rect 266 3159 272 3171
rect 1744 3159 1750 3171
rect 266 3131 1750 3159
rect 266 3119 272 3131
rect 1744 3119 1750 3131
rect 1802 3119 1808 3171
rect 3088 3119 3094 3171
rect 3146 3159 3152 3171
rect 3568 3159 3574 3171
rect 3146 3131 3574 3159
rect 3146 3119 3152 3131
rect 3568 3119 3574 3131
rect 3626 3119 3632 3171
rect 12304 3119 12310 3171
rect 12362 3159 12368 3171
rect 12976 3159 12982 3171
rect 12362 3131 12982 3159
rect 12362 3119 12368 3131
rect 12976 3119 12982 3131
rect 13034 3119 13040 3171
rect 13840 3119 13846 3171
rect 13898 3159 13904 3171
rect 14512 3159 14518 3171
rect 13898 3131 14518 3159
rect 13898 3119 13904 3131
rect 14512 3119 14518 3131
rect 14570 3119 14576 3171
rect 17488 3119 17494 3171
rect 17546 3159 17552 3171
rect 18256 3159 18262 3171
rect 17546 3131 18262 3159
rect 17546 3119 17552 3131
rect 18256 3119 18262 3131
rect 18314 3119 18320 3171
rect 19888 3119 19894 3171
rect 19946 3159 19952 3171
rect 20464 3159 20470 3171
rect 19946 3131 20470 3159
rect 19946 3119 19952 3131
rect 20464 3119 20470 3131
rect 20522 3119 20528 3171
rect 21424 3119 21430 3171
rect 21482 3119 21488 3171
rect 23824 3119 23830 3171
rect 23882 3159 23888 3171
rect 25072 3159 25078 3171
rect 23882 3131 25078 3159
rect 23882 3119 23888 3131
rect 25072 3119 25078 3131
rect 25130 3119 25136 3171
rect 28240 3119 28246 3171
rect 28298 3159 28304 3171
rect 29296 3159 29302 3171
rect 28298 3131 29302 3159
rect 28298 3119 28304 3131
rect 29296 3119 29302 3131
rect 29354 3119 29360 3171
rect 29488 3119 29494 3171
rect 29546 3159 29552 3171
rect 29872 3159 29878 3171
rect 29546 3131 29878 3159
rect 29546 3119 29552 3131
rect 29872 3119 29878 3131
rect 29930 3119 29936 3171
rect 33808 3119 33814 3171
rect 33866 3159 33872 3171
rect 34672 3159 34678 3171
rect 33866 3131 34678 3159
rect 33866 3119 33872 3131
rect 34672 3119 34678 3131
rect 34730 3119 34736 3171
rect 35920 3119 35926 3171
rect 35978 3159 35984 3171
rect 36880 3159 36886 3171
rect 35978 3131 36886 3159
rect 35978 3119 35984 3131
rect 36880 3119 36886 3131
rect 36938 3119 36944 3171
rect 37072 3119 37078 3171
rect 37130 3159 37136 3171
rect 38608 3159 38614 3171
rect 37130 3131 38614 3159
rect 37130 3119 37136 3131
rect 38608 3119 38614 3131
rect 38666 3119 38672 3171
rect 44080 3119 44086 3171
rect 44138 3159 44144 3171
rect 45424 3159 45430 3171
rect 44138 3131 45430 3159
rect 44138 3119 44144 3131
rect 45424 3119 45430 3131
rect 45482 3119 45488 3171
rect 46288 3159 46294 3171
rect 45538 3131 46294 3159
rect 16720 3045 16726 3097
rect 16778 3085 16784 3097
rect 17584 3085 17590 3097
rect 16778 3057 17590 3085
rect 16778 3045 16784 3057
rect 17584 3045 17590 3057
rect 17642 3045 17648 3097
rect 18352 3045 18358 3097
rect 18410 3085 18416 3097
rect 19024 3085 19030 3097
rect 18410 3057 19030 3085
rect 18410 3045 18416 3057
rect 19024 3045 19030 3057
rect 19082 3045 19088 3097
rect 21139 3088 21197 3094
rect 19138 3057 20510 3085
rect 16 2971 22 3023
rect 74 3011 80 3023
rect 1555 3014 1613 3020
rect 1555 3011 1567 3014
rect 74 2983 1567 3011
rect 74 2971 80 2983
rect 1555 2980 1567 2983
rect 1601 2980 1613 3014
rect 2323 3014 2381 3020
rect 2323 3011 2335 3014
rect 1555 2974 1613 2980
rect 1666 2983 2335 3011
rect 688 2897 694 2949
rect 746 2937 752 2949
rect 1666 2937 1694 2983
rect 2323 2980 2335 2983
rect 2369 2980 2381 3014
rect 3091 3014 3149 3020
rect 3091 3011 3103 3014
rect 2323 2974 2381 2980
rect 2866 2983 3103 3011
rect 746 2909 1694 2937
rect 746 2897 752 2909
rect 2128 2897 2134 2949
rect 2186 2937 2192 2949
rect 2866 2937 2894 2983
rect 3091 2980 3103 2983
rect 3137 2980 3149 3014
rect 4912 3011 4918 3023
rect 4873 2983 4918 3011
rect 3091 2974 3149 2980
rect 4912 2971 4918 2983
rect 4970 2971 4976 3023
rect 5200 2971 5206 3023
rect 5258 3011 5264 3023
rect 5683 3014 5741 3020
rect 5683 3011 5695 3014
rect 5258 2983 5695 3011
rect 5258 2971 5264 2983
rect 5683 2980 5695 2983
rect 5729 2980 5741 3014
rect 5683 2974 5741 2980
rect 5968 2971 5974 3023
rect 6026 3011 6032 3023
rect 7027 3014 7085 3020
rect 7027 3011 7039 3014
rect 6026 2983 7039 3011
rect 6026 2971 6032 2983
rect 7027 2980 7039 2983
rect 7073 2980 7085 3014
rect 7027 2974 7085 2980
rect 7795 3014 7853 3020
rect 7795 2980 7807 3014
rect 7841 2980 7853 3014
rect 7795 2974 7853 2980
rect 5776 2937 5782 2949
rect 2186 2909 2894 2937
rect 5218 2909 5782 2937
rect 2186 2897 2192 2909
rect 5104 2749 5110 2801
rect 5162 2789 5168 2801
rect 5218 2789 5246 2909
rect 5776 2897 5782 2909
rect 5834 2897 5840 2949
rect 6736 2897 6742 2949
rect 6794 2937 6800 2949
rect 7810 2937 7838 2974
rect 8176 2971 8182 3023
rect 8234 3011 8240 3023
rect 9715 3014 9773 3020
rect 9715 3011 9727 3014
rect 8234 2983 9727 3011
rect 8234 2971 8240 2983
rect 9715 2980 9727 2983
rect 9761 2980 9773 3014
rect 9715 2974 9773 2980
rect 10483 3014 10541 3020
rect 10483 2980 10495 3014
rect 10529 2980 10541 3014
rect 12976 3011 12982 3023
rect 12937 2983 12982 3011
rect 10483 2974 10541 2980
rect 6794 2909 7838 2937
rect 8467 2940 8525 2946
rect 6794 2897 6800 2909
rect 8467 2906 8479 2940
rect 8513 2937 8525 2940
rect 8513 2909 8798 2937
rect 8513 2906 8525 2909
rect 8467 2900 8525 2906
rect 8770 2875 8798 2909
rect 8944 2897 8950 2949
rect 9002 2937 9008 2949
rect 10498 2937 10526 2974
rect 12976 2971 12982 2983
rect 13034 2971 13040 3023
rect 13360 2971 13366 3023
rect 13418 3011 13424 3023
rect 13747 3014 13805 3020
rect 13747 3011 13759 3014
rect 13418 2983 13759 3011
rect 13418 2971 13424 2983
rect 13747 2980 13759 2983
rect 13793 2980 13805 3014
rect 13747 2974 13805 2980
rect 14512 2971 14518 3023
rect 14570 3011 14576 3023
rect 15091 3014 15149 3020
rect 15091 3011 15103 3014
rect 14570 2983 15103 3011
rect 14570 2971 14576 2983
rect 15091 2980 15103 2983
rect 15137 2980 15149 3014
rect 16624 3011 16630 3023
rect 16585 2983 16630 3011
rect 15091 2974 15149 2980
rect 16624 2971 16630 2983
rect 16682 2971 16688 3023
rect 17008 2971 17014 3023
rect 17066 3011 17072 3023
rect 17779 3014 17837 3020
rect 17779 3011 17791 3014
rect 17066 2983 17791 3011
rect 17066 2971 17072 2983
rect 17779 2980 17791 2983
rect 17825 2980 17837 3014
rect 17779 2974 17837 2980
rect 18547 3014 18605 3020
rect 18547 2980 18559 3014
rect 18593 2980 18605 3014
rect 18547 2974 18605 2980
rect 9002 2909 10526 2937
rect 9002 2897 9008 2909
rect 15376 2897 15382 2949
rect 15434 2937 15440 2949
rect 16432 2937 16438 2949
rect 15434 2909 16438 2937
rect 15434 2897 15440 2909
rect 16432 2897 16438 2909
rect 16490 2897 16496 2949
rect 17680 2897 17686 2949
rect 17738 2937 17744 2949
rect 18562 2937 18590 2974
rect 18832 2971 18838 3023
rect 18890 3011 18896 3023
rect 19138 3011 19166 3057
rect 18890 2983 19166 3011
rect 18890 2971 18896 2983
rect 19312 2971 19318 3023
rect 19370 2971 19376 3023
rect 19600 2971 19606 3023
rect 19658 3011 19664 3023
rect 20482 3020 20510 3057
rect 21139 3054 21151 3088
rect 21185 3085 21197 3088
rect 21442 3085 21470 3119
rect 21185 3057 21470 3085
rect 21185 3054 21197 3057
rect 21139 3048 21197 3054
rect 22384 3045 22390 3097
rect 22442 3085 22448 3097
rect 23536 3085 23542 3097
rect 22442 3057 23542 3085
rect 22442 3045 22448 3057
rect 23536 3045 23542 3057
rect 23594 3045 23600 3097
rect 24595 3088 24653 3094
rect 24595 3054 24607 3088
rect 24641 3085 24653 3088
rect 24880 3085 24886 3097
rect 24641 3057 24886 3085
rect 24641 3054 24653 3057
rect 24595 3048 24653 3054
rect 24880 3045 24886 3057
rect 24938 3045 24944 3097
rect 25360 3045 25366 3097
rect 25418 3085 25424 3097
rect 26224 3085 26230 3097
rect 25418 3057 26230 3085
rect 25418 3045 25424 3057
rect 26224 3045 26230 3057
rect 26282 3045 26288 3097
rect 27472 3045 27478 3097
rect 27530 3085 27536 3097
rect 28912 3085 28918 3097
rect 27530 3057 28918 3085
rect 27530 3045 27536 3057
rect 28912 3045 28918 3057
rect 28970 3045 28976 3097
rect 29392 3045 29398 3097
rect 29450 3085 29456 3097
rect 31120 3085 31126 3097
rect 29450 3057 31126 3085
rect 29450 3045 29456 3057
rect 31120 3045 31126 3057
rect 31178 3045 31184 3097
rect 31888 3045 31894 3097
rect 31946 3085 31952 3097
rect 33328 3085 33334 3097
rect 31946 3057 33334 3085
rect 31946 3045 31952 3057
rect 33328 3045 33334 3057
rect 33386 3045 33392 3097
rect 35632 3045 35638 3097
rect 35690 3085 35696 3097
rect 36112 3085 36118 3097
rect 35690 3057 36118 3085
rect 35690 3045 35696 3057
rect 36112 3045 36118 3057
rect 36170 3045 36176 3097
rect 36688 3045 36694 3097
rect 36746 3085 36752 3097
rect 37552 3085 37558 3097
rect 36746 3057 37558 3085
rect 36746 3045 36752 3057
rect 37552 3045 37558 3057
rect 37610 3045 37616 3097
rect 38320 3045 38326 3097
rect 38378 3085 38384 3097
rect 38378 3057 39422 3085
rect 38378 3045 38384 3057
rect 20467 3014 20525 3020
rect 19658 2983 20318 3011
rect 19658 2971 19664 2983
rect 19330 2937 19358 2971
rect 17738 2909 18590 2937
rect 18658 2909 19358 2937
rect 17738 2897 17744 2909
rect 8752 2863 8758 2875
rect 8713 2835 8758 2863
rect 8752 2823 8758 2835
rect 8810 2823 8816 2875
rect 11443 2866 11501 2872
rect 11443 2832 11455 2866
rect 11489 2863 11501 2866
rect 11489 2835 17294 2863
rect 11489 2832 11501 2835
rect 11443 2826 11501 2832
rect 5162 2761 5246 2789
rect 17266 2789 17294 2835
rect 18256 2823 18262 2875
rect 18314 2863 18320 2875
rect 18658 2863 18686 2909
rect 19792 2897 19798 2949
rect 19850 2937 19856 2949
rect 20176 2937 20182 2949
rect 19850 2909 20182 2937
rect 19850 2897 19856 2909
rect 20176 2897 20182 2909
rect 20234 2897 20240 2949
rect 20290 2937 20318 2983
rect 20467 2980 20479 3014
rect 20513 2980 20525 3014
rect 21235 3014 21293 3020
rect 21235 3011 21247 3014
rect 20467 2974 20525 2980
rect 20578 2983 21247 3011
rect 20578 2937 20606 2983
rect 21235 2980 21247 2983
rect 21281 2980 21293 3014
rect 21235 2974 21293 2980
rect 21424 2971 21430 3023
rect 21482 3011 21488 3023
rect 23155 3014 23213 3020
rect 23155 3011 23167 3014
rect 21482 2983 23167 3011
rect 21482 2971 21488 2983
rect 23155 2980 23167 2983
rect 23201 2980 23213 3014
rect 23155 2974 23213 2980
rect 23923 3014 23981 3020
rect 23923 2980 23935 3014
rect 23969 2980 23981 3014
rect 23923 2974 23981 2980
rect 20848 2937 20854 2949
rect 20290 2909 20606 2937
rect 20674 2909 20854 2937
rect 18314 2835 18686 2863
rect 18314 2823 18320 2835
rect 20464 2823 20470 2875
rect 20522 2863 20528 2875
rect 20674 2863 20702 2909
rect 20848 2897 20854 2909
rect 20906 2897 20912 2949
rect 20944 2897 20950 2949
rect 21002 2937 21008 2949
rect 21712 2937 21718 2949
rect 21002 2909 21718 2937
rect 21002 2897 21008 2909
rect 21712 2897 21718 2909
rect 21770 2897 21776 2949
rect 22480 2897 22486 2949
rect 22538 2937 22544 2949
rect 23938 2937 23966 2974
rect 24016 2971 24022 3023
rect 24074 3011 24080 3023
rect 25843 3014 25901 3020
rect 25843 3011 25855 3014
rect 24074 2983 25855 3011
rect 24074 2971 24080 2983
rect 25843 2980 25855 2983
rect 25889 2980 25901 3014
rect 25843 2974 25901 2980
rect 26611 3014 26669 3020
rect 26611 2980 26623 3014
rect 26657 2980 26669 3014
rect 26611 2974 26669 2980
rect 22538 2909 23966 2937
rect 22538 2897 22544 2909
rect 25072 2897 25078 2949
rect 25130 2937 25136 2949
rect 26626 2937 26654 2974
rect 26896 2971 26902 3023
rect 26954 3011 26960 3023
rect 28531 3014 28589 3020
rect 28531 3011 28543 3014
rect 26954 2983 28543 3011
rect 26954 2971 26960 2983
rect 28531 2980 28543 2983
rect 28577 2980 28589 3014
rect 28531 2974 28589 2980
rect 29299 3014 29357 3020
rect 29299 2980 29311 3014
rect 29345 2980 29357 3014
rect 29299 2974 29357 2980
rect 25130 2909 26654 2937
rect 27283 2940 27341 2946
rect 25130 2897 25136 2909
rect 27283 2906 27295 2940
rect 27329 2937 27341 2940
rect 27329 2909 27614 2937
rect 27329 2906 27341 2909
rect 27283 2900 27341 2906
rect 27586 2872 27614 2909
rect 27664 2897 27670 2949
rect 27722 2937 27728 2949
rect 29314 2937 29342 2974
rect 29872 2971 29878 3023
rect 29930 3011 29936 3023
rect 31219 3014 31277 3020
rect 31219 3011 31231 3014
rect 29930 2983 31231 3011
rect 29930 2971 29936 2983
rect 31219 2980 31231 2983
rect 31265 2980 31277 3014
rect 31219 2974 31277 2980
rect 31987 3014 32045 3020
rect 31987 2980 31999 3014
rect 32033 2980 32045 3014
rect 31987 2974 32045 2980
rect 27722 2909 29342 2937
rect 27722 2897 27728 2909
rect 30544 2897 30550 2949
rect 30602 2937 30608 2949
rect 32002 2937 32030 2974
rect 32080 2971 32086 3023
rect 32138 3011 32144 3023
rect 33907 3014 33965 3020
rect 33907 3011 33919 3014
rect 32138 2983 33919 3011
rect 32138 2971 32144 2983
rect 33907 2980 33919 2983
rect 33953 2980 33965 3014
rect 33907 2974 33965 2980
rect 34675 3014 34733 3020
rect 34675 2980 34687 3014
rect 34721 2980 34733 3014
rect 34675 2974 34733 2980
rect 30602 2909 32030 2937
rect 30602 2897 30608 2909
rect 32272 2897 32278 2949
rect 32330 2937 32336 2949
rect 33136 2937 33142 2949
rect 32330 2909 33142 2937
rect 32330 2897 32336 2909
rect 33136 2897 33142 2909
rect 33194 2897 33200 2949
rect 33328 2897 33334 2949
rect 33386 2937 33392 2949
rect 34690 2937 34718 2974
rect 35440 2971 35446 3023
rect 35498 3011 35504 3023
rect 36595 3014 36653 3020
rect 36595 3011 36607 3014
rect 35498 2983 36607 3011
rect 35498 2971 35504 2983
rect 36595 2980 36607 2983
rect 36641 2980 36653 3014
rect 36595 2974 36653 2980
rect 37363 3014 37421 3020
rect 37363 2980 37375 3014
rect 37409 2980 37421 3014
rect 39283 3014 39341 3020
rect 39283 3011 39295 3014
rect 37363 2974 37421 2980
rect 37570 2983 39295 3011
rect 33386 2909 34718 2937
rect 33386 2897 33392 2909
rect 35344 2897 35350 2949
rect 35402 2937 35408 2949
rect 36016 2937 36022 2949
rect 35402 2909 36022 2937
rect 35402 2897 35408 2909
rect 36016 2897 36022 2909
rect 36074 2897 36080 2949
rect 36112 2897 36118 2949
rect 36170 2937 36176 2949
rect 37378 2937 37406 2974
rect 37570 2949 37598 2983
rect 39283 2980 39295 2983
rect 39329 2980 39341 3014
rect 39394 3011 39422 3057
rect 39664 3045 39670 3097
rect 39722 3085 39728 3097
rect 40912 3085 40918 3097
rect 39722 3057 40918 3085
rect 39722 3045 39728 3057
rect 40912 3045 40918 3057
rect 40970 3045 40976 3097
rect 41104 3045 41110 3097
rect 41162 3085 41168 3097
rect 42064 3085 42070 3097
rect 41162 3057 42070 3085
rect 41162 3045 41168 3057
rect 42064 3045 42070 3057
rect 42122 3045 42128 3097
rect 42544 3045 42550 3097
rect 42602 3085 42608 3097
rect 43312 3085 43318 3097
rect 42602 3057 43318 3085
rect 42602 3045 42608 3057
rect 43312 3045 43318 3057
rect 43370 3045 43376 3097
rect 44464 3045 44470 3097
rect 44522 3085 44528 3097
rect 45136 3085 45142 3097
rect 44522 3057 45142 3085
rect 44522 3045 44528 3057
rect 45136 3045 45142 3057
rect 45194 3045 45200 3097
rect 40051 3014 40109 3020
rect 40051 3011 40063 3014
rect 39394 2983 40063 3011
rect 39283 2974 39341 2980
rect 40051 2980 40063 2983
rect 40097 2980 40109 3014
rect 40051 2974 40109 2980
rect 40528 2971 40534 3023
rect 40586 3011 40592 3023
rect 41971 3014 42029 3020
rect 41971 3011 41983 3014
rect 40586 2983 41983 3011
rect 40586 2971 40592 2983
rect 41971 2980 41983 2983
rect 42017 2980 42029 3014
rect 41971 2974 42029 2980
rect 42739 3014 42797 3020
rect 42739 2980 42751 3014
rect 42785 2980 42797 3014
rect 44659 3014 44717 3020
rect 44659 3011 44671 3014
rect 42739 2974 42797 2980
rect 43042 2983 44671 3011
rect 36170 2909 37406 2937
rect 36170 2897 36176 2909
rect 37552 2897 37558 2949
rect 37610 2897 37616 2949
rect 38128 2897 38134 2949
rect 38186 2937 38192 2949
rect 39088 2937 39094 2949
rect 38186 2909 39094 2937
rect 38186 2897 38192 2909
rect 39088 2897 39094 2909
rect 39146 2897 39152 2949
rect 41200 2897 41206 2949
rect 41258 2937 41264 2949
rect 42754 2937 42782 2974
rect 41258 2909 42782 2937
rect 41258 2897 41264 2909
rect 20522 2835 20702 2863
rect 21139 2866 21197 2872
rect 20522 2823 20528 2835
rect 21139 2832 21151 2866
rect 21185 2832 21197 2866
rect 21139 2826 21197 2832
rect 27571 2866 27629 2872
rect 27571 2832 27583 2866
rect 27617 2863 27629 2866
rect 27952 2863 27958 2875
rect 27617 2835 27958 2863
rect 27617 2832 27629 2835
rect 27571 2826 27629 2832
rect 21154 2789 21182 2826
rect 27952 2823 27958 2835
rect 28010 2823 28016 2875
rect 30259 2866 30317 2872
rect 30259 2832 30271 2866
rect 30305 2863 30317 2866
rect 33040 2863 33046 2875
rect 30305 2835 33046 2863
rect 30305 2832 30317 2835
rect 30259 2826 30317 2832
rect 33040 2823 33046 2835
rect 33098 2823 33104 2875
rect 35248 2823 35254 2875
rect 35306 2863 35312 2875
rect 38323 2866 38381 2872
rect 38323 2863 38335 2866
rect 35306 2835 38335 2863
rect 35306 2823 35312 2835
rect 38323 2832 38335 2835
rect 38369 2832 38381 2866
rect 38323 2826 38381 2832
rect 43042 2801 43070 2983
rect 44659 2980 44671 2983
rect 44705 2980 44717 3014
rect 44659 2974 44717 2980
rect 45427 3014 45485 3020
rect 45427 2980 45439 3014
rect 45473 2980 45485 3014
rect 45427 2974 45485 2980
rect 43312 2897 43318 2949
rect 43370 2937 43376 2949
rect 43504 2937 43510 2949
rect 43370 2909 43510 2937
rect 43370 2897 43376 2909
rect 43504 2897 43510 2909
rect 43562 2897 43568 2949
rect 43984 2937 43990 2949
rect 43618 2909 43990 2937
rect 41008 2789 41014 2801
rect 17266 2761 21182 2789
rect 40969 2761 41014 2789
rect 5162 2749 5168 2761
rect 41008 2749 41014 2761
rect 41066 2749 41072 2801
rect 43024 2749 43030 2801
rect 43082 2749 43088 2801
rect 43216 2749 43222 2801
rect 43274 2789 43280 2801
rect 43618 2789 43646 2909
rect 43984 2897 43990 2909
rect 44042 2897 44048 2949
rect 44176 2897 44182 2949
rect 44234 2937 44240 2949
rect 45442 2937 45470 2974
rect 44234 2909 45470 2937
rect 44234 2897 44240 2909
rect 45136 2823 45142 2875
rect 45194 2863 45200 2875
rect 45538 2863 45566 3131
rect 46288 3119 46294 3131
rect 46346 3119 46352 3171
rect 48112 3119 48118 3171
rect 48170 3159 48176 3171
rect 48976 3159 48982 3171
rect 48170 3131 48982 3159
rect 48170 3119 48176 3131
rect 48976 3119 48982 3131
rect 49034 3119 49040 3171
rect 46192 3045 46198 3097
rect 46250 3085 46256 3097
rect 47632 3085 47638 3097
rect 46250 3057 47638 3085
rect 46250 3045 46256 3057
rect 47632 3045 47638 3057
rect 47690 3045 47696 3097
rect 51760 3045 51766 3097
rect 51818 3085 51824 3097
rect 52240 3085 52246 3097
rect 51818 3057 52246 3085
rect 51818 3045 51824 3057
rect 52240 3045 52246 3057
rect 52298 3045 52304 3097
rect 45616 2971 45622 3023
rect 45674 3011 45680 3023
rect 47347 3014 47405 3020
rect 47347 3011 47359 3014
rect 45674 2983 47359 3011
rect 45674 2971 45680 2983
rect 47347 2980 47359 2983
rect 47393 2980 47405 3014
rect 48115 3014 48173 3020
rect 48115 3011 48127 3014
rect 47347 2974 47405 2980
rect 47506 2983 48127 3011
rect 46288 2897 46294 2949
rect 46346 2937 46352 2949
rect 47506 2937 47534 2983
rect 48115 2980 48127 2983
rect 48161 2980 48173 3014
rect 48115 2974 48173 2980
rect 49648 2971 49654 3023
rect 49706 3011 49712 3023
rect 50035 3014 50093 3020
rect 50035 3011 50047 3014
rect 49706 2983 50047 3011
rect 49706 2971 49712 2983
rect 50035 2980 50047 2983
rect 50081 2980 50093 3014
rect 50035 2974 50093 2980
rect 50803 3014 50861 3020
rect 50803 2980 50815 3014
rect 50849 2980 50861 3014
rect 50803 2974 50861 2980
rect 46346 2909 47534 2937
rect 46346 2897 46352 2909
rect 47632 2897 47638 2949
rect 47690 2937 47696 2949
rect 48880 2937 48886 2949
rect 47690 2909 48886 2937
rect 47690 2897 47696 2909
rect 48880 2897 48886 2909
rect 48938 2897 48944 2949
rect 48976 2897 48982 2949
rect 49034 2937 49040 2949
rect 49840 2937 49846 2949
rect 49034 2909 49846 2937
rect 49034 2897 49040 2909
rect 49840 2897 49846 2909
rect 49898 2897 49904 2949
rect 50818 2937 50846 2974
rect 51472 2971 51478 3023
rect 51530 3011 51536 3023
rect 52723 3014 52781 3020
rect 52723 3011 52735 3014
rect 51530 2983 52735 3011
rect 51530 2971 51536 2983
rect 52723 2980 52735 2983
rect 52769 2980 52781 3014
rect 53491 3014 53549 3020
rect 53491 3011 53503 3014
rect 52723 2974 52781 2980
rect 52834 2983 53503 3011
rect 50050 2909 50846 2937
rect 50050 2875 50078 2909
rect 51376 2897 51382 2949
rect 51434 2937 51440 2949
rect 51856 2937 51862 2949
rect 51434 2909 51862 2937
rect 51434 2897 51440 2909
rect 51856 2897 51862 2909
rect 51914 2897 51920 2949
rect 52240 2897 52246 2949
rect 52298 2937 52304 2949
rect 52834 2937 52862 2983
rect 53491 2980 53503 2983
rect 53537 2980 53549 3014
rect 53491 2974 53549 2980
rect 53776 2971 53782 3023
rect 53834 3011 53840 3023
rect 55411 3014 55469 3020
rect 55411 3011 55423 3014
rect 53834 2983 55423 3011
rect 53834 2971 53840 2983
rect 55411 2980 55423 2983
rect 55457 2980 55469 3014
rect 55411 2974 55469 2980
rect 56179 3014 56237 3020
rect 56179 2980 56191 3014
rect 56225 2980 56237 3014
rect 56179 2974 56237 2980
rect 52298 2909 52862 2937
rect 52298 2897 52304 2909
rect 52912 2897 52918 2949
rect 52970 2937 52976 2949
rect 53680 2937 53686 2949
rect 52970 2909 53686 2937
rect 52970 2897 52976 2909
rect 53680 2897 53686 2909
rect 53738 2897 53744 2949
rect 54832 2897 54838 2949
rect 54890 2937 54896 2949
rect 56194 2937 56222 2974
rect 54890 2909 56222 2937
rect 54890 2897 54896 2909
rect 45194 2835 45566 2863
rect 45194 2823 45200 2835
rect 50032 2823 50038 2875
rect 50090 2823 50096 2875
rect 46384 2789 46390 2801
rect 43274 2761 43646 2789
rect 46345 2761 46390 2789
rect 43274 2749 43280 2761
rect 46384 2749 46390 2761
rect 46442 2749 46448 2801
rect 49075 2792 49133 2798
rect 49075 2758 49087 2792
rect 49121 2789 49133 2792
rect 52432 2789 52438 2801
rect 49121 2761 52438 2789
rect 49121 2758 49133 2761
rect 49075 2752 49133 2758
rect 52432 2749 52438 2761
rect 52490 2749 52496 2801
rect 1152 2690 58848 2712
rect 1152 2638 4294 2690
rect 4346 2638 4358 2690
rect 4410 2638 4422 2690
rect 4474 2638 4486 2690
rect 4538 2638 35014 2690
rect 35066 2638 35078 2690
rect 35130 2638 35142 2690
rect 35194 2638 35206 2690
rect 35258 2638 58848 2690
rect 1152 2616 58848 2638
rect 3952 2527 3958 2579
rect 4010 2567 4016 2579
rect 4240 2567 4246 2579
rect 4010 2539 4246 2567
rect 4010 2527 4016 2539
rect 4240 2527 4246 2539
rect 4298 2527 4304 2579
rect 4336 2527 4342 2579
rect 4394 2567 4400 2579
rect 4816 2567 4822 2579
rect 4394 2539 4822 2567
rect 4394 2527 4400 2539
rect 4816 2527 4822 2539
rect 4874 2527 4880 2579
rect 13744 2527 13750 2579
rect 13802 2567 13808 2579
rect 46384 2567 46390 2579
rect 13802 2539 46390 2567
rect 13802 2527 13808 2539
rect 46384 2527 46390 2539
rect 46442 2527 46448 2579
rect 19408 2453 19414 2505
rect 19466 2493 19472 2505
rect 19888 2493 19894 2505
rect 19466 2465 19894 2493
rect 19466 2453 19472 2465
rect 19888 2453 19894 2465
rect 19946 2453 19952 2505
rect 46096 2453 46102 2505
rect 46154 2493 46160 2505
rect 47056 2493 47062 2505
rect 46154 2465 47062 2493
rect 46154 2453 46160 2465
rect 47056 2453 47062 2465
rect 47114 2453 47120 2505
rect 41008 2379 41014 2431
rect 41066 2419 41072 2431
rect 49264 2419 49270 2431
rect 41066 2391 49270 2419
rect 41066 2379 41072 2391
rect 49264 2379 49270 2391
rect 49322 2379 49328 2431
rect 4720 2009 4726 2061
rect 4778 2049 4784 2061
rect 5296 2049 5302 2061
rect 4778 2021 5302 2049
rect 4778 2009 4784 2021
rect 5296 2009 5302 2021
rect 5354 2009 5360 2061
rect 4528 1861 4534 1913
rect 4586 1901 4592 1913
rect 4816 1901 4822 1913
rect 4586 1873 4822 1901
rect 4586 1861 4592 1873
rect 4816 1861 4822 1873
rect 4874 1861 4880 1913
rect 20176 1787 20182 1839
rect 20234 1827 20240 1839
rect 21232 1827 21238 1839
rect 20234 1799 21238 1827
rect 20234 1787 20240 1799
rect 21232 1787 21238 1799
rect 21290 1787 21296 1839
rect 30352 1713 30358 1765
rect 30410 1753 30416 1765
rect 30640 1753 30646 1765
rect 30410 1725 30646 1753
rect 30410 1713 30416 1725
rect 30640 1713 30646 1725
rect 30698 1713 30704 1765
rect 50512 1713 50518 1765
rect 50570 1753 50576 1765
rect 51088 1753 51094 1765
rect 50570 1725 51094 1753
rect 50570 1713 50576 1725
rect 51088 1713 51094 1725
rect 51146 1713 51152 1765
rect 36112 1639 36118 1691
rect 36170 1639 36176 1691
rect 35632 1565 35638 1617
rect 35690 1565 35696 1617
rect 35650 1531 35678 1565
rect 34882 1503 35678 1531
rect 34882 1321 34910 1503
rect 35152 1417 35158 1469
rect 35210 1457 35216 1469
rect 35536 1457 35542 1469
rect 35210 1429 35542 1457
rect 35210 1417 35216 1429
rect 35536 1417 35542 1429
rect 35594 1417 35600 1469
rect 35632 1417 35638 1469
rect 35690 1457 35696 1469
rect 35920 1457 35926 1469
rect 35690 1429 35926 1457
rect 35690 1417 35696 1429
rect 35920 1417 35926 1429
rect 35978 1417 35984 1469
rect 36130 1321 36158 1639
rect 50704 1565 50710 1617
rect 50762 1605 50768 1617
rect 50896 1605 50902 1617
rect 50762 1577 50902 1605
rect 50762 1565 50768 1577
rect 50896 1565 50902 1577
rect 50954 1565 50960 1617
rect 36304 1491 36310 1543
rect 36362 1491 36368 1543
rect 33232 1269 33238 1321
rect 33290 1309 33296 1321
rect 33712 1309 33718 1321
rect 33290 1281 33718 1309
rect 33290 1269 33296 1281
rect 33712 1269 33718 1281
rect 33770 1269 33776 1321
rect 34864 1269 34870 1321
rect 34922 1269 34928 1321
rect 36112 1269 36118 1321
rect 36170 1269 36176 1321
rect 36322 1173 36350 1491
rect 41008 1417 41014 1469
rect 41066 1457 41072 1469
rect 41296 1457 41302 1469
rect 41066 1429 41302 1457
rect 41066 1417 41072 1429
rect 41296 1417 41302 1429
rect 41354 1417 41360 1469
rect 50896 1417 50902 1469
rect 50954 1457 50960 1469
rect 51568 1457 51574 1469
rect 50954 1429 51574 1457
rect 50954 1417 50960 1429
rect 51568 1417 51574 1429
rect 51626 1417 51632 1469
rect 36304 1121 36310 1173
rect 36362 1121 36368 1173
rect 35440 1047 35446 1099
rect 35498 1087 35504 1099
rect 37264 1087 37270 1099
rect 35498 1059 37270 1087
rect 35498 1047 35504 1059
rect 37264 1047 37270 1059
rect 37322 1047 37328 1099
<< via1 >>
rect 4294 57250 4346 57302
rect 4358 57250 4410 57302
rect 4422 57250 4474 57302
rect 4486 57250 4538 57302
rect 35014 57250 35066 57302
rect 35078 57250 35130 57302
rect 35142 57250 35194 57302
rect 35206 57250 35258 57302
rect 1750 56991 1802 57043
rect 214 56917 266 56969
rect 3286 56991 3338 57043
rect 4918 56917 4970 56969
rect 9622 56991 9674 57043
rect 11254 56991 11306 57043
rect 6454 56917 6506 56969
rect 8086 56960 8138 56969
rect 8086 56926 8095 56960
rect 8095 56926 8129 56960
rect 8129 56926 8138 56960
rect 8086 56917 8138 56926
rect 16438 56991 16490 57043
rect 29110 56991 29162 57043
rect 12790 56917 12842 56969
rect 14422 56917 14474 56969
rect 15958 56917 16010 56969
rect 17494 56917 17546 56969
rect 19126 56917 19178 56969
rect 20662 56917 20714 56969
rect 22294 56917 22346 56969
rect 23830 56917 23882 56969
rect 25462 56917 25514 56969
rect 26998 56917 27050 56969
rect 28630 56960 28682 56969
rect 28630 56926 28639 56960
rect 28639 56926 28673 56960
rect 28673 56926 28682 56960
rect 28630 56917 28682 56926
rect 30262 56960 30314 56969
rect 30262 56926 30271 56960
rect 30271 56926 30305 56960
rect 30305 56926 30314 56960
rect 30262 56917 30314 56926
rect 31702 56960 31754 56969
rect 31702 56926 31711 56960
rect 31711 56926 31745 56960
rect 31745 56926 31754 56960
rect 31702 56917 31754 56926
rect 33334 56917 33386 56969
rect 34870 56960 34922 56969
rect 34870 56926 34879 56960
rect 34879 56926 34913 56960
rect 34913 56926 34922 56960
rect 34870 56917 34922 56926
rect 38038 56960 38090 56969
rect 38038 56926 38047 56960
rect 38047 56926 38081 56960
rect 38081 56926 38090 56960
rect 38038 56917 38090 56926
rect 41206 56917 41258 56969
rect 44374 56917 44426 56969
rect 47542 56960 47594 56969
rect 47542 56926 47551 56960
rect 47551 56926 47585 56960
rect 47585 56926 47594 56960
rect 47542 56917 47594 56926
rect 53878 56960 53930 56969
rect 53878 56926 53887 56960
rect 53887 56926 53921 56960
rect 53921 56926 53930 56960
rect 53878 56917 53930 56926
rect 3670 56843 3722 56895
rect 5110 56886 5162 56895
rect 5110 56852 5119 56886
rect 5119 56852 5153 56886
rect 5153 56852 5162 56886
rect 5110 56843 5162 56852
rect 8278 56843 8330 56895
rect 11254 56886 11306 56895
rect 11254 56852 11263 56886
rect 11263 56852 11297 56886
rect 11297 56852 11306 56886
rect 11254 56843 11306 56852
rect 12982 56886 13034 56895
rect 12982 56852 12991 56886
rect 12991 56852 13025 56886
rect 13025 56852 13034 56886
rect 12982 56843 13034 56852
rect 13654 56843 13706 56895
rect 16150 56886 16202 56895
rect 16150 56852 16159 56886
rect 16159 56852 16193 56886
rect 16193 56852 16202 56886
rect 16150 56843 16202 56852
rect 17974 56886 18026 56895
rect 17974 56852 17983 56886
rect 17983 56852 18017 56886
rect 18017 56852 18026 56886
rect 17974 56843 18026 56852
rect 19318 56886 19370 56895
rect 19318 56852 19327 56886
rect 19327 56852 19361 56886
rect 19361 56852 19370 56886
rect 19318 56843 19370 56852
rect 24022 56886 24074 56895
rect 3574 56769 3626 56821
rect 10774 56769 10826 56821
rect 24022 56852 24031 56886
rect 24031 56852 24065 56886
rect 24065 56852 24074 56886
rect 24022 56843 24074 56852
rect 27190 56886 27242 56895
rect 27190 56852 27199 56886
rect 27199 56852 27233 56886
rect 27233 56852 27242 56886
rect 27190 56843 27242 56852
rect 29974 56843 30026 56895
rect 34102 56886 34154 56895
rect 34102 56852 34111 56886
rect 34111 56852 34145 56886
rect 34145 56852 34154 56886
rect 34102 56843 34154 56852
rect 36502 56843 36554 56895
rect 39670 56843 39722 56895
rect 40630 56843 40682 56895
rect 42838 56843 42890 56895
rect 46102 56843 46154 56895
rect 49078 56843 49130 56895
rect 50710 56843 50762 56895
rect 52246 56843 52298 56895
rect 55414 56843 55466 56895
rect 57046 56886 57098 56895
rect 57046 56852 57055 56886
rect 57055 56852 57089 56886
rect 57089 56852 57098 56886
rect 57046 56843 57098 56852
rect 40342 56769 40394 56821
rect 9814 56738 9866 56747
rect 9814 56704 9823 56738
rect 9823 56704 9857 56738
rect 9857 56704 9866 56738
rect 9814 56695 9866 56704
rect 13654 56738 13706 56747
rect 13654 56704 13663 56738
rect 13663 56704 13697 56738
rect 13697 56704 13706 56738
rect 13654 56695 13706 56704
rect 36694 56738 36746 56747
rect 36694 56704 36703 56738
rect 36703 56704 36737 56738
rect 36737 56704 36746 56738
rect 36694 56695 36746 56704
rect 39766 56738 39818 56747
rect 39766 56704 39775 56738
rect 39775 56704 39809 56738
rect 39809 56704 39818 56738
rect 39766 56695 39818 56704
rect 40822 56738 40874 56747
rect 40822 56704 40831 56738
rect 40831 56704 40865 56738
rect 40865 56704 40874 56738
rect 40822 56695 40874 56704
rect 42934 56738 42986 56747
rect 42934 56704 42943 56738
rect 42943 56704 42977 56738
rect 42977 56704 42986 56738
rect 42934 56695 42986 56704
rect 46102 56695 46154 56747
rect 48694 56738 48746 56747
rect 48694 56704 48703 56738
rect 48703 56704 48737 56738
rect 48737 56704 48746 56738
rect 48694 56695 48746 56704
rect 50806 56738 50858 56747
rect 50806 56704 50815 56738
rect 50815 56704 50849 56738
rect 50849 56704 50858 56738
rect 50806 56695 50858 56704
rect 52822 56738 52874 56747
rect 52822 56704 52831 56738
rect 52831 56704 52865 56738
rect 52865 56704 52874 56738
rect 52822 56695 52874 56704
rect 55414 56695 55466 56747
rect 56758 56738 56810 56747
rect 56758 56704 56767 56738
rect 56767 56704 56801 56738
rect 56801 56704 56810 56738
rect 56758 56695 56810 56704
rect 19654 56584 19706 56636
rect 19718 56584 19770 56636
rect 19782 56584 19834 56636
rect 19846 56584 19898 56636
rect 50374 56584 50426 56636
rect 50438 56584 50490 56636
rect 50502 56584 50554 56636
rect 50566 56584 50618 56636
rect 694 56473 746 56525
rect 2230 56473 2282 56525
rect 2806 56473 2858 56525
rect 3862 56473 3914 56525
rect 5398 56473 5450 56525
rect 5974 56473 6026 56525
rect 7030 56473 7082 56525
rect 8566 56516 8618 56525
rect 8566 56482 8575 56516
rect 8575 56482 8609 56516
rect 8609 56482 8618 56516
rect 8566 56473 8618 56482
rect 10198 56473 10250 56525
rect 10678 56473 10730 56525
rect 11734 56473 11786 56525
rect 12310 56473 12362 56525
rect 13366 56473 13418 56525
rect 14902 56473 14954 56525
rect 17014 56473 17066 56525
rect 18070 56473 18122 56525
rect 18550 56473 18602 56525
rect 19990 56473 20042 56525
rect 21238 56473 21290 56525
rect 21718 56473 21770 56525
rect 22774 56473 22826 56525
rect 24406 56473 24458 56525
rect 25942 56473 25994 56525
rect 26518 56473 26570 56525
rect 27574 56473 27626 56525
rect 28054 56473 28106 56525
rect 29686 56516 29738 56525
rect 29686 56482 29695 56516
rect 29695 56482 29729 56516
rect 29729 56482 29738 56516
rect 29686 56473 29738 56482
rect 30646 56473 30698 56525
rect 31222 56473 31274 56525
rect 32278 56473 32330 56525
rect 33814 56473 33866 56525
rect 34582 56473 34634 56525
rect 36022 56473 36074 56525
rect 37558 56473 37610 56525
rect 38614 56473 38666 56525
rect 40150 56516 40202 56525
rect 40150 56482 40159 56516
rect 40159 56482 40193 56516
rect 40193 56482 40202 56516
rect 40150 56473 40202 56482
rect 41782 56473 41834 56525
rect 42262 56473 42314 56525
rect 43318 56473 43370 56525
rect 43894 56473 43946 56525
rect 44950 56473 45002 56525
rect 46486 56473 46538 56525
rect 48022 56473 48074 56525
rect 49654 56473 49706 56525
rect 50134 56473 50186 56525
rect 52918 56473 52970 56525
rect 53302 56473 53354 56525
rect 54358 56473 54410 56525
rect 54934 56473 54986 56525
rect 55990 56473 56042 56525
rect 26614 56399 26666 56451
rect 56758 56399 56810 56451
rect 11446 56325 11498 56377
rect 12214 56325 12266 56377
rect 28726 56325 28778 56377
rect 43894 56325 43946 56377
rect 2710 56251 2762 56303
rect 2806 56251 2858 56303
rect 42550 56251 42602 56303
rect 58582 56251 58634 56303
rect 2614 56177 2666 56229
rect 3286 56220 3338 56229
rect 3286 56186 3295 56220
rect 3295 56186 3329 56220
rect 3329 56186 3338 56220
rect 3286 56177 3338 56186
rect 5590 56220 5642 56229
rect 5590 56186 5599 56220
rect 5599 56186 5633 56220
rect 5633 56186 5642 56220
rect 5590 56177 5642 56186
rect 5974 56220 6026 56229
rect 5974 56186 5983 56220
rect 5983 56186 6017 56220
rect 6017 56186 6026 56220
rect 5974 56177 6026 56186
rect 7222 56220 7274 56229
rect 7222 56186 7231 56220
rect 7231 56186 7265 56220
rect 7265 56186 7274 56220
rect 8182 56220 8234 56229
rect 7222 56177 7274 56186
rect 8182 56186 8191 56220
rect 8191 56186 8225 56220
rect 8225 56186 8234 56220
rect 8182 56177 8234 56186
rect 10102 56220 10154 56229
rect 10102 56186 10111 56220
rect 10111 56186 10145 56220
rect 10145 56186 10154 56220
rect 10102 56177 10154 56186
rect 11158 56220 11210 56229
rect 11158 56186 11167 56220
rect 11167 56186 11201 56220
rect 11201 56186 11210 56220
rect 11158 56177 11210 56186
rect 11926 56220 11978 56229
rect 11926 56186 11935 56220
rect 11935 56186 11969 56220
rect 11969 56186 11978 56220
rect 11926 56177 11978 56186
rect 12694 56220 12746 56229
rect 12694 56186 12703 56220
rect 12703 56186 12737 56220
rect 12737 56186 12746 56220
rect 12694 56177 12746 56186
rect 13270 56220 13322 56229
rect 13270 56186 13279 56220
rect 13279 56186 13313 56220
rect 13313 56186 13322 56220
rect 13270 56177 13322 56186
rect 15094 56220 15146 56229
rect 15094 56186 15103 56220
rect 15103 56186 15137 56220
rect 15137 56186 15146 56220
rect 15094 56177 15146 56186
rect 17206 56220 17258 56229
rect 15382 56103 15434 56155
rect 17206 56186 17215 56220
rect 17215 56186 17249 56220
rect 17249 56186 17258 56220
rect 17206 56177 17258 56186
rect 18262 56220 18314 56229
rect 18262 56186 18271 56220
rect 18271 56186 18305 56220
rect 18305 56186 18314 56220
rect 18262 56177 18314 56186
rect 20374 56220 20426 56229
rect 20374 56186 20383 56220
rect 20383 56186 20417 56220
rect 20417 56186 20426 56220
rect 20374 56177 20426 56186
rect 21430 56220 21482 56229
rect 21430 56186 21439 56220
rect 21439 56186 21473 56220
rect 21473 56186 21482 56220
rect 21430 56177 21482 56186
rect 22198 56220 22250 56229
rect 22198 56186 22207 56220
rect 22207 56186 22241 56220
rect 22241 56186 22250 56220
rect 22198 56177 22250 56186
rect 22966 56220 23018 56229
rect 22966 56186 22975 56220
rect 22975 56186 23009 56220
rect 23009 56186 23018 56220
rect 26134 56220 26186 56229
rect 22966 56177 23018 56186
rect 26134 56186 26143 56220
rect 26143 56186 26177 56220
rect 26177 56186 26186 56220
rect 26134 56177 26186 56186
rect 26806 56220 26858 56229
rect 26806 56186 26815 56220
rect 26815 56186 26849 56220
rect 26849 56186 26858 56220
rect 26806 56177 26858 56186
rect 27478 56220 27530 56229
rect 27478 56186 27487 56220
rect 27487 56186 27521 56220
rect 27521 56186 27530 56220
rect 27478 56177 27530 56186
rect 28150 56220 28202 56229
rect 28150 56186 28159 56220
rect 28159 56186 28193 56220
rect 28193 56186 28202 56220
rect 28150 56177 28202 56186
rect 29302 56220 29354 56229
rect 29302 56186 29311 56220
rect 29311 56186 29345 56220
rect 29345 56186 29354 56220
rect 29302 56177 29354 56186
rect 30934 56220 30986 56229
rect 30934 56186 30943 56220
rect 30943 56186 30977 56220
rect 30977 56186 30986 56220
rect 30934 56177 30986 56186
rect 31702 56220 31754 56229
rect 31702 56186 31711 56220
rect 31711 56186 31745 56220
rect 31745 56186 31754 56220
rect 31702 56177 31754 56186
rect 32470 56220 32522 56229
rect 32470 56186 32479 56220
rect 32479 56186 32513 56220
rect 32513 56186 32522 56220
rect 32470 56177 32522 56186
rect 32854 56220 32906 56229
rect 32854 56186 32863 56220
rect 32863 56186 32897 56220
rect 32897 56186 32906 56220
rect 32854 56177 32906 56186
rect 34006 56220 34058 56229
rect 32758 56103 32810 56155
rect 34006 56186 34015 56220
rect 34015 56186 34049 56220
rect 34049 56186 34058 56220
rect 34006 56177 34058 56186
rect 34390 56220 34442 56229
rect 34390 56186 34399 56220
rect 34399 56186 34433 56220
rect 34433 56186 34442 56220
rect 34390 56177 34442 56186
rect 35830 56220 35882 56229
rect 35830 56186 35839 56220
rect 35839 56186 35873 56220
rect 35873 56186 35882 56220
rect 35830 56177 35882 56186
rect 35446 56103 35498 56155
rect 36790 56177 36842 56229
rect 37750 56220 37802 56229
rect 37750 56186 37759 56220
rect 37759 56186 37793 56220
rect 37793 56186 37802 56220
rect 37750 56177 37802 56186
rect 38710 56220 38762 56229
rect 38710 56186 38719 56220
rect 38719 56186 38753 56220
rect 38753 56186 38762 56220
rect 38710 56177 38762 56186
rect 39862 56220 39914 56229
rect 39862 56186 39871 56220
rect 39871 56186 39905 56220
rect 39905 56186 39914 56220
rect 39862 56177 39914 56186
rect 41974 56220 42026 56229
rect 41974 56186 41983 56220
rect 41983 56186 42017 56220
rect 42017 56186 42026 56220
rect 41974 56177 42026 56186
rect 42646 56220 42698 56229
rect 42646 56186 42655 56220
rect 42655 56186 42689 56220
rect 42689 56186 42698 56220
rect 42646 56177 42698 56186
rect 43606 56177 43658 56229
rect 44182 56220 44234 56229
rect 44182 56186 44191 56220
rect 44191 56186 44225 56220
rect 44225 56186 44234 56220
rect 44182 56177 44234 56186
rect 45046 56220 45098 56229
rect 45046 56186 45055 56220
rect 45055 56186 45089 56220
rect 45089 56186 45098 56220
rect 45046 56177 45098 56186
rect 46774 56220 46826 56229
rect 46774 56186 46783 56220
rect 46783 56186 46817 56220
rect 46817 56186 46826 56220
rect 46774 56177 46826 56186
rect 48214 56220 48266 56229
rect 48214 56186 48223 56220
rect 48223 56186 48257 56220
rect 48257 56186 48266 56220
rect 48214 56177 48266 56186
rect 48790 56177 48842 56229
rect 37078 56103 37130 56155
rect 40822 56103 40874 56155
rect 48598 56103 48650 56155
rect 38806 56029 38858 56081
rect 49942 56177 49994 56229
rect 51670 56220 51722 56229
rect 51670 56186 51679 56220
rect 51679 56186 51713 56220
rect 51713 56186 51722 56220
rect 51670 56177 51722 56186
rect 53686 56220 53738 56229
rect 51190 56103 51242 56155
rect 53686 56186 53695 56220
rect 53695 56186 53729 56220
rect 53729 56186 53738 56220
rect 53686 56177 53738 56186
rect 54550 56220 54602 56229
rect 54550 56186 54559 56220
rect 54559 56186 54593 56220
rect 54593 56186 54602 56220
rect 54550 56177 54602 56186
rect 55510 56220 55562 56229
rect 55510 56186 55519 56220
rect 55519 56186 55553 56220
rect 55553 56186 55562 56220
rect 55510 56177 55562 56186
rect 4294 55918 4346 55970
rect 4358 55918 4410 55970
rect 4422 55918 4474 55970
rect 4486 55918 4538 55970
rect 35014 55918 35066 55970
rect 35078 55918 35130 55970
rect 35142 55918 35194 55970
rect 35206 55918 35258 55970
rect 3766 55733 3818 55785
rect 11926 55733 11978 55785
rect 1174 55659 1226 55711
rect 4630 55659 4682 55711
rect 7510 55659 7562 55711
rect 9142 55659 9194 55711
rect 13846 55659 13898 55711
rect 5014 55585 5066 55637
rect 20182 55659 20234 55711
rect 23350 55659 23402 55711
rect 24886 55659 24938 55711
rect 39094 55659 39146 55711
rect 40726 55659 40778 55711
rect 45430 55659 45482 55711
rect 46966 55659 47018 55711
rect 51766 55659 51818 55711
rect 56470 55659 56522 55711
rect 57526 55659 57578 55711
rect 1750 55554 1802 55563
rect 1750 55520 1759 55554
rect 1759 55520 1793 55554
rect 1793 55520 1802 55554
rect 1750 55511 1802 55520
rect 4630 55511 4682 55563
rect 7702 55554 7754 55563
rect 7702 55520 7711 55554
rect 7711 55520 7745 55554
rect 7745 55520 7754 55554
rect 7702 55511 7754 55520
rect 12790 55554 12842 55563
rect 12790 55520 12799 55554
rect 12799 55520 12833 55554
rect 12833 55520 12842 55554
rect 12790 55511 12842 55520
rect 16534 55511 16586 55563
rect 20278 55511 20330 55563
rect 23158 55511 23210 55563
rect 24886 55511 24938 55563
rect 25654 55554 25706 55563
rect 25654 55520 25663 55554
rect 25663 55520 25697 55554
rect 25697 55520 25706 55554
rect 25654 55511 25706 55520
rect 52630 55585 52682 55637
rect 38806 55437 38858 55489
rect 8950 55406 9002 55415
rect 8950 55372 8959 55406
rect 8959 55372 8993 55406
rect 8993 55372 9002 55406
rect 8950 55363 9002 55372
rect 23158 55406 23210 55415
rect 23158 55372 23167 55406
rect 23167 55372 23201 55406
rect 23201 55372 23210 55406
rect 23158 55363 23210 55372
rect 24886 55363 24938 55415
rect 25654 55363 25706 55415
rect 38902 55406 38954 55415
rect 38902 55372 38911 55406
rect 38911 55372 38945 55406
rect 38945 55372 38954 55406
rect 38902 55363 38954 55372
rect 40438 55363 40490 55415
rect 42166 55406 42218 55415
rect 42166 55372 42175 55406
rect 42175 55372 42209 55406
rect 42209 55372 42218 55406
rect 45238 55406 45290 55415
rect 42166 55363 42218 55372
rect 45238 55372 45247 55406
rect 45247 55372 45281 55406
rect 45281 55372 45290 55406
rect 45238 55363 45290 55372
rect 46582 55363 46634 55415
rect 51574 55406 51626 55415
rect 51574 55372 51583 55406
rect 51583 55372 51617 55406
rect 51617 55372 51626 55406
rect 51574 55363 51626 55372
rect 55606 55406 55658 55415
rect 55606 55372 55615 55406
rect 55615 55372 55649 55406
rect 55649 55372 55658 55406
rect 55606 55363 55658 55372
rect 56278 55406 56330 55415
rect 56278 55372 56287 55406
rect 56287 55372 56321 55406
rect 56321 55372 56330 55406
rect 57334 55406 57386 55415
rect 56278 55363 56330 55372
rect 57334 55372 57343 55406
rect 57343 55372 57377 55406
rect 57377 55372 57386 55406
rect 57334 55363 57386 55372
rect 19654 55252 19706 55304
rect 19718 55252 19770 55304
rect 19782 55252 19834 55304
rect 19846 55252 19898 55304
rect 50374 55252 50426 55304
rect 50438 55252 50490 55304
rect 50502 55252 50554 55304
rect 50566 55252 50618 55304
rect 19990 55141 20042 55193
rect 55606 55141 55658 55193
rect 59158 55141 59210 55193
rect 11446 54993 11498 55045
rect 58006 54845 58058 54897
rect 30070 54697 30122 54749
rect 44662 54740 44714 54749
rect 44662 54706 44671 54740
rect 44671 54706 44705 54740
rect 44705 54706 44714 54740
rect 44662 54697 44714 54706
rect 55798 54740 55850 54749
rect 55798 54706 55807 54740
rect 55807 54706 55841 54740
rect 55841 54706 55850 54740
rect 55798 54697 55850 54706
rect 4294 54586 4346 54638
rect 4358 54586 4410 54638
rect 4422 54586 4474 54638
rect 4486 54586 4538 54638
rect 35014 54586 35066 54638
rect 35078 54586 35130 54638
rect 35142 54586 35194 54638
rect 35206 54586 35258 54638
rect 58102 54327 58154 54379
rect 53014 54179 53066 54231
rect 57622 54222 57674 54231
rect 57622 54188 57631 54222
rect 57631 54188 57665 54222
rect 57665 54188 57674 54222
rect 57622 54179 57674 54188
rect 36502 54105 36554 54157
rect 36886 54105 36938 54157
rect 55798 54105 55850 54157
rect 19654 53920 19706 53972
rect 19718 53920 19770 53972
rect 19782 53920 19834 53972
rect 19846 53920 19898 53972
rect 50374 53920 50426 53972
rect 50438 53920 50490 53972
rect 50502 53920 50554 53972
rect 50566 53920 50618 53972
rect 10870 53809 10922 53861
rect 57622 53809 57674 53861
rect 59638 53809 59690 53861
rect 6454 53365 6506 53417
rect 57622 53408 57674 53417
rect 57622 53374 57631 53408
rect 57631 53374 57665 53408
rect 57665 53374 57674 53408
rect 57622 53365 57674 53374
rect 4294 53254 4346 53306
rect 4358 53254 4410 53306
rect 4422 53254 4474 53306
rect 4486 53254 4538 53306
rect 35014 53254 35066 53306
rect 35078 53254 35130 53306
rect 35142 53254 35194 53306
rect 35206 53254 35258 53306
rect 48886 52847 48938 52899
rect 30934 52773 30986 52825
rect 22678 52699 22730 52751
rect 19654 52588 19706 52640
rect 19718 52588 19770 52640
rect 19782 52588 19834 52640
rect 19846 52588 19898 52640
rect 50374 52588 50426 52640
rect 50438 52588 50490 52640
rect 50502 52588 50554 52640
rect 50566 52588 50618 52640
rect 46774 52181 46826 52233
rect 42838 52076 42890 52085
rect 42838 52042 42847 52076
rect 42847 52042 42881 52076
rect 42881 52042 42890 52076
rect 42838 52033 42890 52042
rect 4294 51922 4346 51974
rect 4358 51922 4410 51974
rect 4422 51922 4474 51974
rect 4486 51922 4538 51974
rect 35014 51922 35066 51974
rect 35078 51922 35130 51974
rect 35142 51922 35194 51974
rect 35206 51922 35258 51974
rect 1942 51558 1994 51567
rect 1942 51524 1951 51558
rect 1951 51524 1985 51558
rect 1985 51524 1994 51558
rect 1942 51515 1994 51524
rect 52918 51515 52970 51567
rect 48598 51441 48650 51493
rect 19654 51256 19706 51308
rect 19718 51256 19770 51308
rect 19782 51256 19834 51308
rect 19846 51256 19898 51308
rect 50374 51256 50426 51308
rect 50438 51256 50490 51308
rect 50502 51256 50554 51308
rect 50566 51256 50618 51308
rect 1942 51145 1994 51197
rect 32374 51145 32426 51197
rect 31318 50701 31370 50753
rect 31510 50744 31562 50753
rect 31510 50710 31519 50744
rect 31519 50710 31553 50744
rect 31553 50710 31562 50744
rect 31510 50701 31562 50710
rect 4294 50590 4346 50642
rect 4358 50590 4410 50642
rect 4422 50590 4474 50642
rect 4486 50590 4538 50642
rect 35014 50590 35066 50642
rect 35078 50590 35130 50642
rect 35142 50590 35194 50642
rect 35206 50590 35258 50642
rect 23830 50479 23882 50531
rect 31510 50479 31562 50531
rect 31318 50405 31370 50457
rect 42262 50405 42314 50457
rect 56854 50257 56906 50309
rect 49174 50226 49226 50235
rect 49174 50192 49183 50226
rect 49183 50192 49217 50226
rect 49217 50192 49226 50226
rect 49174 50183 49226 50192
rect 31798 50109 31850 50161
rect 49174 50035 49226 50087
rect 19654 49924 19706 49976
rect 19718 49924 19770 49976
rect 19782 49924 19834 49976
rect 19846 49924 19898 49976
rect 50374 49924 50426 49976
rect 50438 49924 50490 49976
rect 50502 49924 50554 49976
rect 50566 49924 50618 49976
rect 38422 49412 38474 49421
rect 38422 49378 38431 49412
rect 38431 49378 38465 49412
rect 38465 49378 38474 49412
rect 38422 49369 38474 49378
rect 51286 49369 51338 49421
rect 52054 49412 52106 49421
rect 52054 49378 52063 49412
rect 52063 49378 52097 49412
rect 52097 49378 52106 49412
rect 52054 49369 52106 49378
rect 4294 49258 4346 49310
rect 4358 49258 4410 49310
rect 4422 49258 4474 49310
rect 4486 49258 4538 49310
rect 35014 49258 35066 49310
rect 35078 49258 35130 49310
rect 35142 49258 35194 49310
rect 35206 49258 35258 49310
rect 40342 49147 40394 49199
rect 30934 49073 30986 49125
rect 52054 49073 52106 49125
rect 38422 48999 38474 49051
rect 48982 48999 49034 49051
rect 55606 48925 55658 48977
rect 47830 48703 47882 48755
rect 19654 48592 19706 48644
rect 19718 48592 19770 48644
rect 19782 48592 19834 48644
rect 19846 48592 19898 48644
rect 50374 48592 50426 48644
rect 50438 48592 50490 48644
rect 50502 48592 50554 48644
rect 50566 48592 50618 48644
rect 10966 48037 11018 48089
rect 4294 47926 4346 47978
rect 4358 47926 4410 47978
rect 4422 47926 4474 47978
rect 4486 47926 4538 47978
rect 35014 47926 35066 47978
rect 35078 47926 35130 47978
rect 35142 47926 35194 47978
rect 35206 47926 35258 47978
rect 28726 47815 28778 47867
rect 34198 47593 34250 47645
rect 54262 47519 54314 47571
rect 19654 47260 19706 47312
rect 19718 47260 19770 47312
rect 19782 47260 19834 47312
rect 19846 47260 19898 47312
rect 50374 47260 50426 47312
rect 50438 47260 50490 47312
rect 50502 47260 50554 47312
rect 50566 47260 50618 47312
rect 2614 47149 2666 47201
rect 19126 46779 19178 46831
rect 10678 46705 10730 46757
rect 4294 46594 4346 46646
rect 4358 46594 4410 46646
rect 4422 46594 4474 46646
rect 4486 46594 4538 46646
rect 35014 46594 35066 46646
rect 35078 46594 35130 46646
rect 35142 46594 35194 46646
rect 35206 46594 35258 46646
rect 6070 46483 6122 46535
rect 10678 46483 10730 46535
rect 10870 46526 10922 46535
rect 10870 46492 10879 46526
rect 10879 46492 10913 46526
rect 10913 46492 10922 46526
rect 10870 46483 10922 46492
rect 33814 46261 33866 46313
rect 41974 46187 42026 46239
rect 7222 46039 7274 46091
rect 41110 46113 41162 46165
rect 19654 45928 19706 45980
rect 19718 45928 19770 45980
rect 19782 45928 19834 45980
rect 19846 45928 19898 45980
rect 50374 45928 50426 45980
rect 50438 45928 50490 45980
rect 50502 45928 50554 45980
rect 50566 45928 50618 45980
rect 6550 45416 6602 45425
rect 6550 45382 6559 45416
rect 6559 45382 6593 45416
rect 6593 45382 6602 45416
rect 6550 45373 6602 45382
rect 41014 45373 41066 45425
rect 4294 45262 4346 45314
rect 4358 45262 4410 45314
rect 4422 45262 4474 45314
rect 4486 45262 4538 45314
rect 35014 45262 35066 45314
rect 35078 45262 35130 45314
rect 35142 45262 35194 45314
rect 35206 45262 35258 45314
rect 6550 45151 6602 45203
rect 53206 45151 53258 45203
rect 37462 44707 37514 44759
rect 44854 44707 44906 44759
rect 19654 44596 19706 44648
rect 19718 44596 19770 44648
rect 19782 44596 19834 44648
rect 19846 44596 19898 44648
rect 50374 44596 50426 44648
rect 50438 44596 50490 44648
rect 50502 44596 50554 44648
rect 50566 44596 50618 44648
rect 26134 44115 26186 44167
rect 17110 44084 17162 44093
rect 17110 44050 17119 44084
rect 17119 44050 17153 44084
rect 17153 44050 17162 44084
rect 17110 44041 17162 44050
rect 4294 43930 4346 43982
rect 4358 43930 4410 43982
rect 4422 43930 4474 43982
rect 4486 43930 4538 43982
rect 35014 43930 35066 43982
rect 35078 43930 35130 43982
rect 35142 43930 35194 43982
rect 35206 43930 35258 43982
rect 12310 43375 12362 43427
rect 19654 43264 19706 43316
rect 19718 43264 19770 43316
rect 19782 43264 19834 43316
rect 19846 43264 19898 43316
rect 50374 43264 50426 43316
rect 50438 43264 50490 43316
rect 50502 43264 50554 43316
rect 50566 43264 50618 43316
rect 1846 42709 1898 42761
rect 4294 42598 4346 42650
rect 4358 42598 4410 42650
rect 4422 42598 4474 42650
rect 4486 42598 4538 42650
rect 35014 42598 35066 42650
rect 35078 42598 35130 42650
rect 35142 42598 35194 42650
rect 35206 42598 35258 42650
rect 39670 42191 39722 42243
rect 18262 42117 18314 42169
rect 5590 42043 5642 42095
rect 46294 42086 46346 42095
rect 46294 42052 46303 42086
rect 46303 42052 46337 42086
rect 46337 42052 46346 42086
rect 46294 42043 46346 42052
rect 19654 41932 19706 41984
rect 19718 41932 19770 41984
rect 19782 41932 19834 41984
rect 19846 41932 19898 41984
rect 50374 41932 50426 41984
rect 50438 41932 50490 41984
rect 50502 41932 50554 41984
rect 50566 41932 50618 41984
rect 17206 41377 17258 41429
rect 25750 41377 25802 41429
rect 4294 41266 4346 41318
rect 4358 41266 4410 41318
rect 4422 41266 4474 41318
rect 4486 41266 4538 41318
rect 35014 41266 35066 41318
rect 35078 41266 35130 41318
rect 35142 41266 35194 41318
rect 35206 41266 35258 41318
rect 25750 41155 25802 41207
rect 46198 41155 46250 41207
rect 42742 40859 42794 40911
rect 29110 40785 29162 40837
rect 45142 40711 45194 40763
rect 19654 40600 19706 40652
rect 19718 40600 19770 40652
rect 19782 40600 19834 40652
rect 19846 40600 19898 40652
rect 50374 40600 50426 40652
rect 50438 40600 50490 40652
rect 50502 40600 50554 40652
rect 50566 40600 50618 40652
rect 57334 40341 57386 40393
rect 32950 40088 33002 40097
rect 32950 40054 32959 40088
rect 32959 40054 32993 40088
rect 32993 40054 33002 40088
rect 32950 40045 33002 40054
rect 4294 39934 4346 39986
rect 4358 39934 4410 39986
rect 4422 39934 4474 39986
rect 4486 39934 4538 39986
rect 35014 39934 35066 39986
rect 35078 39934 35130 39986
rect 35142 39934 35194 39986
rect 35206 39934 35258 39986
rect 23926 39379 23978 39431
rect 19654 39268 19706 39320
rect 19718 39268 19770 39320
rect 19782 39268 19834 39320
rect 19846 39268 19898 39320
rect 50374 39268 50426 39320
rect 50438 39268 50490 39320
rect 50502 39268 50554 39320
rect 50566 39268 50618 39320
rect 11158 38787 11210 38839
rect 12598 38756 12650 38765
rect 12598 38722 12607 38756
rect 12607 38722 12641 38756
rect 12641 38722 12650 38756
rect 12598 38713 12650 38722
rect 24118 38756 24170 38765
rect 24118 38722 24127 38756
rect 24127 38722 24161 38756
rect 24161 38722 24170 38756
rect 24118 38713 24170 38722
rect 52342 38756 52394 38765
rect 52342 38722 52351 38756
rect 52351 38722 52385 38756
rect 52385 38722 52394 38756
rect 52342 38713 52394 38722
rect 4294 38602 4346 38654
rect 4358 38602 4410 38654
rect 4422 38602 4474 38654
rect 4486 38602 4538 38654
rect 35014 38602 35066 38654
rect 35078 38602 35130 38654
rect 35142 38602 35194 38654
rect 35206 38602 35258 38654
rect 12598 38491 12650 38543
rect 55990 38491 56042 38543
rect 11350 38417 11402 38469
rect 52342 38417 52394 38469
rect 4054 38047 4106 38099
rect 50230 38195 50282 38247
rect 19654 37936 19706 37988
rect 19718 37936 19770 37988
rect 19782 37936 19834 37988
rect 19846 37936 19898 37988
rect 50374 37936 50426 37988
rect 50438 37936 50490 37988
rect 50502 37936 50554 37988
rect 50566 37936 50618 37988
rect 11158 37381 11210 37433
rect 20278 37381 20330 37433
rect 29590 37424 29642 37433
rect 29590 37390 29599 37424
rect 29599 37390 29633 37424
rect 29633 37390 29642 37424
rect 29590 37381 29642 37390
rect 4294 37270 4346 37322
rect 4358 37270 4410 37322
rect 4422 37270 4474 37322
rect 4486 37270 4538 37322
rect 35014 37270 35066 37322
rect 35078 37270 35130 37322
rect 35142 37270 35194 37322
rect 35206 37270 35258 37322
rect 5014 37202 5066 37211
rect 5014 37168 5023 37202
rect 5023 37168 5057 37202
rect 5057 37168 5066 37202
rect 5014 37159 5066 37168
rect 11158 37159 11210 37211
rect 30262 37159 30314 37211
rect 51766 36863 51818 36915
rect 19654 36604 19706 36656
rect 19718 36604 19770 36656
rect 19782 36604 19834 36656
rect 19846 36604 19898 36656
rect 50374 36604 50426 36656
rect 50438 36604 50490 36656
rect 50502 36604 50554 36656
rect 50566 36604 50618 36656
rect 2806 36493 2858 36545
rect 16438 36092 16490 36101
rect 16438 36058 16447 36092
rect 16447 36058 16481 36092
rect 16481 36058 16490 36092
rect 16438 36049 16490 36058
rect 56278 36049 56330 36101
rect 4294 35938 4346 35990
rect 4358 35938 4410 35990
rect 4422 35938 4474 35990
rect 4486 35938 4538 35990
rect 35014 35938 35066 35990
rect 35078 35938 35130 35990
rect 35142 35938 35194 35990
rect 35206 35938 35258 35990
rect 13078 35531 13130 35583
rect 22966 35531 23018 35583
rect 5302 35383 5354 35435
rect 13078 35426 13130 35435
rect 13078 35392 13087 35426
rect 13087 35392 13121 35426
rect 13121 35392 13130 35426
rect 13078 35383 13130 35392
rect 19654 35272 19706 35324
rect 19718 35272 19770 35324
rect 19782 35272 19834 35324
rect 19846 35272 19898 35324
rect 50374 35272 50426 35324
rect 50438 35272 50490 35324
rect 50502 35272 50554 35324
rect 50566 35272 50618 35324
rect 32470 35013 32522 35065
rect 22294 34865 22346 34917
rect 12694 34791 12746 34843
rect 12598 34717 12650 34769
rect 36598 34791 36650 34843
rect 43414 34791 43466 34843
rect 28534 34760 28586 34769
rect 28534 34726 28543 34760
rect 28543 34726 28577 34760
rect 28577 34726 28586 34760
rect 28534 34717 28586 34726
rect 4294 34606 4346 34658
rect 4358 34606 4410 34658
rect 4422 34606 4474 34658
rect 4486 34606 4538 34658
rect 35014 34606 35066 34658
rect 35078 34606 35130 34658
rect 35142 34606 35194 34658
rect 35206 34606 35258 34658
rect 22966 34242 23018 34251
rect 22966 34208 22975 34242
rect 22975 34208 23009 34242
rect 23009 34208 23018 34242
rect 22966 34199 23018 34208
rect 56950 34199 57002 34251
rect 19654 33940 19706 33992
rect 19718 33940 19770 33992
rect 19782 33940 19834 33992
rect 19846 33940 19898 33992
rect 50374 33940 50426 33992
rect 50438 33940 50490 33992
rect 50502 33940 50554 33992
rect 50566 33940 50618 33992
rect 34582 33607 34634 33659
rect 12502 33533 12554 33585
rect 15958 33385 16010 33437
rect 48214 33533 48266 33585
rect 43126 33428 43178 33437
rect 43126 33394 43135 33428
rect 43135 33394 43169 33428
rect 43169 33394 43178 33428
rect 43126 33385 43178 33394
rect 4294 33274 4346 33326
rect 4358 33274 4410 33326
rect 4422 33274 4474 33326
rect 4486 33274 4538 33326
rect 35014 33274 35066 33326
rect 35078 33274 35130 33326
rect 35142 33274 35194 33326
rect 35206 33274 35258 33326
rect 13750 33163 13802 33215
rect 43126 33163 43178 33215
rect 49654 33163 49706 33215
rect 2710 33015 2762 33067
rect 29494 32941 29546 32993
rect 33238 32719 33290 32771
rect 19654 32608 19706 32660
rect 19718 32608 19770 32660
rect 19782 32608 19834 32660
rect 19846 32608 19898 32660
rect 50374 32608 50426 32660
rect 50438 32608 50490 32660
rect 50502 32608 50554 32660
rect 50566 32608 50618 32660
rect 53686 32127 53738 32179
rect 32182 32096 32234 32105
rect 32182 32062 32191 32096
rect 32191 32062 32225 32096
rect 32225 32062 32234 32096
rect 32182 32053 32234 32062
rect 39286 32053 39338 32105
rect 4294 31942 4346 31994
rect 4358 31942 4410 31994
rect 4422 31942 4474 31994
rect 4486 31942 4538 31994
rect 35014 31942 35066 31994
rect 35078 31942 35130 31994
rect 35142 31942 35194 31994
rect 35206 31942 35258 31994
rect 32182 31831 32234 31883
rect 52054 31831 52106 31883
rect 21238 31683 21290 31735
rect 36118 31683 36170 31735
rect 20374 31609 20426 31661
rect 19654 31276 19706 31328
rect 19718 31276 19770 31328
rect 19782 31276 19834 31328
rect 19846 31276 19898 31328
rect 50374 31276 50426 31328
rect 50438 31276 50490 31328
rect 50502 31276 50554 31328
rect 50566 31276 50618 31328
rect 54550 31017 54602 31069
rect 35446 30721 35498 30773
rect 4294 30610 4346 30662
rect 4358 30610 4410 30662
rect 4422 30610 4474 30662
rect 4486 30610 4538 30662
rect 35014 30610 35066 30662
rect 35078 30610 35130 30662
rect 35142 30610 35194 30662
rect 35206 30610 35258 30662
rect 16246 30277 16298 30329
rect 19654 29944 19706 29996
rect 19718 29944 19770 29996
rect 19782 29944 19834 29996
rect 19846 29944 19898 29996
rect 50374 29944 50426 29996
rect 50438 29944 50490 29996
rect 50502 29944 50554 29996
rect 50566 29944 50618 29996
rect 13270 29611 13322 29663
rect 8662 29537 8714 29589
rect 18838 29537 18890 29589
rect 8278 29463 8330 29515
rect 17878 29463 17930 29515
rect 18358 29432 18410 29441
rect 18358 29398 18367 29432
rect 18367 29398 18401 29432
rect 18401 29398 18410 29432
rect 18358 29389 18410 29398
rect 4294 29278 4346 29330
rect 4358 29278 4410 29330
rect 4422 29278 4474 29330
rect 4486 29278 4538 29330
rect 35014 29278 35066 29330
rect 35078 29278 35130 29330
rect 35142 29278 35194 29330
rect 35206 29278 35258 29330
rect 8230 28871 8282 28923
rect 8662 28871 8714 28923
rect 10102 28797 10154 28849
rect 8615 28723 8667 28775
rect 19654 28612 19706 28664
rect 19718 28612 19770 28664
rect 19782 28612 19834 28664
rect 19846 28612 19898 28664
rect 50374 28612 50426 28664
rect 50438 28612 50490 28664
rect 50502 28612 50554 28664
rect 50566 28612 50618 28664
rect 8615 28501 8667 28553
rect 18934 28501 18986 28553
rect 5974 28279 6026 28331
rect 14422 28279 14474 28331
rect 3286 28205 3338 28257
rect 8182 28131 8234 28183
rect 18070 28131 18122 28183
rect 6550 28057 6602 28109
rect 21334 28100 21386 28109
rect 21334 28066 21343 28100
rect 21343 28066 21377 28100
rect 21377 28066 21386 28100
rect 21334 28057 21386 28066
rect 29014 28057 29066 28109
rect 4294 27946 4346 27998
rect 4358 27946 4410 27998
rect 4422 27946 4474 27998
rect 4486 27946 4538 27998
rect 35014 27946 35066 27998
rect 35078 27946 35130 27998
rect 35142 27946 35194 27998
rect 35206 27946 35258 27998
rect 9334 27835 9386 27887
rect 12694 27835 12746 27887
rect 14422 27878 14474 27887
rect 14422 27844 14431 27878
rect 14431 27844 14465 27878
rect 14465 27844 14474 27878
rect 14422 27835 14474 27844
rect 21334 27835 21386 27887
rect 48118 27835 48170 27887
rect 5398 27539 5450 27591
rect 26230 27539 26282 27591
rect 8182 27465 8234 27517
rect 9334 27465 9386 27517
rect 9046 27391 9098 27443
rect 9622 27391 9674 27443
rect 16822 27391 16874 27443
rect 19654 27280 19706 27332
rect 19718 27280 19770 27332
rect 19782 27280 19834 27332
rect 19846 27280 19898 27332
rect 50374 27280 50426 27332
rect 50438 27280 50490 27332
rect 50502 27280 50554 27332
rect 50566 27280 50618 27332
rect 31702 27169 31754 27221
rect 1942 26873 1994 26925
rect 34870 26873 34922 26925
rect 18166 26799 18218 26851
rect 26422 26725 26474 26777
rect 36214 26768 36266 26777
rect 36214 26734 36223 26768
rect 36223 26734 36257 26768
rect 36257 26734 36266 26768
rect 36214 26725 36266 26734
rect 4294 26614 4346 26666
rect 4358 26614 4410 26666
rect 4422 26614 4474 26666
rect 4486 26614 4538 26666
rect 35014 26614 35066 26666
rect 35078 26614 35130 26666
rect 35142 26614 35194 26666
rect 35206 26614 35258 26666
rect 1942 26546 1994 26555
rect 1942 26512 1951 26546
rect 1951 26512 1985 26546
rect 1985 26512 1994 26546
rect 1942 26503 1994 26512
rect 10870 26503 10922 26555
rect 12118 26429 12170 26481
rect 37750 26207 37802 26259
rect 17014 26059 17066 26111
rect 19654 25948 19706 26000
rect 19718 25948 19770 26000
rect 19782 25948 19834 26000
rect 19846 25948 19898 26000
rect 50374 25948 50426 26000
rect 50438 25948 50490 26000
rect 50502 25948 50554 26000
rect 50566 25948 50618 26000
rect 40726 25541 40778 25593
rect 12022 25467 12074 25519
rect 4294 25282 4346 25334
rect 4358 25282 4410 25334
rect 4422 25282 4474 25334
rect 4486 25282 4538 25334
rect 35014 25282 35066 25334
rect 35078 25282 35130 25334
rect 35142 25282 35194 25334
rect 35206 25282 35258 25334
rect 11062 25171 11114 25223
rect 8086 24949 8138 25001
rect 26902 24875 26954 24927
rect 31702 24875 31754 24927
rect 51190 24875 51242 24927
rect 8758 24727 8810 24779
rect 19654 24616 19706 24668
rect 19718 24616 19770 24668
rect 19782 24616 19834 24668
rect 19846 24616 19898 24668
rect 50374 24616 50426 24668
rect 50438 24616 50490 24668
rect 50502 24616 50554 24668
rect 50566 24616 50618 24668
rect 8086 24505 8138 24557
rect 14134 24505 14186 24557
rect 35350 24135 35402 24187
rect 31990 24061 32042 24113
rect 44758 24061 44810 24113
rect 4294 23950 4346 24002
rect 4358 23950 4410 24002
rect 4422 23950 4474 24002
rect 4486 23950 4538 24002
rect 35014 23950 35066 24002
rect 35078 23950 35130 24002
rect 35142 23950 35194 24002
rect 35206 23950 35258 24002
rect 25462 23839 25514 23891
rect 31990 23839 32042 23891
rect 15478 23765 15530 23817
rect 34390 23617 34442 23669
rect 41878 23543 41930 23595
rect 46966 23586 47018 23595
rect 8086 23469 8138 23521
rect 13270 23469 13322 23521
rect 29398 23469 29450 23521
rect 46966 23552 46975 23586
rect 46975 23552 47009 23586
rect 47009 23552 47018 23586
rect 46966 23543 47018 23552
rect 8470 23395 8522 23447
rect 49750 23395 49802 23447
rect 19654 23284 19706 23336
rect 19718 23284 19770 23336
rect 19782 23284 19834 23336
rect 19846 23284 19898 23336
rect 50374 23284 50426 23336
rect 50438 23284 50490 23336
rect 50502 23284 50554 23336
rect 50566 23284 50618 23336
rect 8086 23173 8138 23225
rect 13174 23173 13226 23225
rect 8470 23099 8522 23151
rect 14038 23099 14090 23151
rect 10582 22877 10634 22929
rect 55414 22877 55466 22929
rect 8086 22803 8138 22855
rect 26614 22803 26666 22855
rect 46678 22803 46730 22855
rect 37558 22772 37610 22781
rect 37558 22738 37567 22772
rect 37567 22738 37601 22772
rect 37601 22738 37610 22772
rect 37558 22729 37610 22738
rect 4294 22618 4346 22670
rect 4358 22618 4410 22670
rect 4422 22618 4474 22670
rect 4486 22618 4538 22670
rect 35014 22618 35066 22670
rect 35078 22618 35130 22670
rect 35142 22618 35194 22670
rect 35206 22618 35258 22670
rect 25750 22507 25802 22559
rect 37558 22507 37610 22559
rect 57622 22433 57674 22485
rect 8086 22285 8138 22337
rect 10582 22137 10634 22189
rect 19654 21952 19706 22004
rect 19718 21952 19770 22004
rect 19782 21952 19834 22004
rect 19846 21952 19898 22004
rect 50374 21952 50426 22004
rect 50438 21952 50490 22004
rect 50502 21952 50554 22004
rect 50566 21952 50618 22004
rect 43894 21619 43946 21671
rect 8086 21545 8138 21597
rect 48694 21545 48746 21597
rect 8566 21397 8618 21449
rect 52822 21471 52874 21523
rect 33046 21397 33098 21449
rect 4294 21286 4346 21338
rect 4358 21286 4410 21338
rect 4422 21286 4474 21338
rect 4486 21286 4538 21338
rect 35014 21286 35066 21338
rect 35078 21286 35130 21338
rect 35142 21286 35194 21338
rect 35206 21286 35258 21338
rect 8086 20899 8138 20951
rect 50806 20879 50858 20931
rect 7606 20774 7658 20783
rect 7606 20740 7615 20774
rect 7615 20740 7649 20774
rect 7649 20740 7658 20774
rect 7606 20731 7658 20740
rect 8566 20731 8618 20783
rect 8758 20731 8810 20783
rect 9334 20731 9386 20783
rect 55510 20731 55562 20783
rect 19654 20620 19706 20672
rect 19718 20620 19770 20672
rect 19782 20620 19834 20672
rect 19846 20620 19898 20672
rect 50374 20620 50426 20672
rect 50438 20620 50490 20672
rect 50502 20620 50554 20672
rect 50566 20620 50618 20672
rect 7606 20509 7658 20561
rect 8758 20509 8810 20561
rect 9334 20509 9386 20561
rect 44182 20139 44234 20191
rect 7606 20065 7658 20117
rect 8758 20065 8810 20117
rect 16726 20065 16778 20117
rect 32566 20065 32618 20117
rect 4294 19954 4346 20006
rect 4358 19954 4410 20006
rect 4422 19954 4474 20006
rect 4486 19954 4538 20006
rect 35014 19954 35066 20006
rect 35078 19954 35130 20006
rect 35142 19954 35194 20006
rect 35206 19954 35258 20006
rect 7606 19886 7658 19895
rect 7606 19852 7615 19886
rect 7615 19852 7649 19886
rect 7649 19852 7658 19886
rect 7606 19843 7658 19852
rect 8758 19843 8810 19895
rect 48790 19843 48842 19895
rect 16726 19769 16778 19821
rect 40342 19769 40394 19821
rect 7126 19590 7178 19599
rect 7126 19556 7135 19590
rect 7135 19556 7169 19590
rect 7169 19556 7178 19590
rect 7126 19547 7178 19556
rect 34774 19590 34826 19599
rect 34774 19556 34783 19590
rect 34783 19556 34817 19590
rect 34817 19556 34826 19590
rect 34774 19547 34826 19556
rect 8278 19473 8330 19525
rect 9046 19473 9098 19525
rect 46102 19473 46154 19525
rect 19654 19288 19706 19340
rect 19718 19288 19770 19340
rect 19782 19288 19834 19340
rect 19846 19288 19898 19340
rect 50374 19288 50426 19340
rect 50438 19288 50490 19340
rect 50502 19288 50554 19340
rect 50566 19288 50618 19340
rect 7126 19177 7178 19229
rect 49846 19177 49898 19229
rect 2518 19103 2570 19155
rect 34774 19103 34826 19155
rect 39862 18881 39914 18933
rect 21238 18776 21290 18785
rect 21238 18742 21247 18776
rect 21247 18742 21281 18776
rect 21281 18742 21290 18776
rect 21238 18733 21290 18742
rect 47638 18733 47690 18785
rect 4294 18622 4346 18674
rect 4358 18622 4410 18674
rect 4422 18622 4474 18674
rect 4486 18622 4538 18674
rect 35014 18622 35066 18674
rect 35078 18622 35130 18674
rect 35142 18622 35194 18674
rect 35206 18622 35258 18674
rect 45238 18437 45290 18489
rect 7414 18215 7466 18267
rect 8086 18215 8138 18267
rect 47158 18289 47210 18341
rect 40726 18258 40778 18267
rect 40726 18224 40735 18258
rect 40735 18224 40769 18258
rect 40769 18224 40778 18258
rect 40726 18215 40778 18224
rect 51670 18289 51722 18341
rect 50998 18110 51050 18119
rect 50998 18076 51007 18110
rect 51007 18076 51041 18110
rect 51041 18076 51050 18110
rect 50998 18067 51050 18076
rect 19654 17956 19706 18008
rect 19718 17956 19770 18008
rect 19782 17956 19834 18008
rect 19846 17956 19898 18008
rect 50374 17956 50426 18008
rect 50438 17956 50490 18008
rect 50502 17956 50554 18008
rect 50566 17956 50618 18008
rect 7798 17845 7850 17897
rect 50998 17771 51050 17823
rect 8086 17697 8138 17749
rect 42934 17697 42986 17749
rect 35830 17623 35882 17675
rect 7414 17475 7466 17527
rect 8566 17475 8618 17527
rect 23734 17401 23786 17453
rect 4294 17290 4346 17342
rect 4358 17290 4410 17342
rect 4422 17290 4474 17342
rect 4486 17290 4538 17342
rect 35014 17290 35066 17342
rect 35078 17290 35130 17342
rect 35142 17290 35194 17342
rect 35206 17290 35258 17342
rect 15094 16957 15146 17009
rect 5974 16926 6026 16935
rect 5974 16892 5983 16926
rect 5983 16892 6017 16926
rect 6017 16892 6026 16926
rect 5974 16883 6026 16892
rect 7126 16926 7178 16935
rect 7126 16892 7135 16926
rect 7135 16892 7169 16926
rect 7169 16892 7178 16926
rect 7126 16883 7178 16892
rect 46870 16926 46922 16935
rect 46870 16892 46879 16926
rect 46879 16892 46913 16926
rect 46913 16892 46922 16926
rect 46870 16883 46922 16892
rect 55990 16926 56042 16935
rect 55990 16892 55999 16926
rect 55999 16892 56033 16926
rect 56033 16892 56042 16926
rect 55990 16883 56042 16892
rect 39766 16809 39818 16861
rect 42646 16735 42698 16787
rect 19654 16624 19706 16676
rect 19718 16624 19770 16676
rect 19782 16624 19834 16676
rect 19846 16624 19898 16676
rect 50374 16624 50426 16676
rect 50438 16624 50490 16676
rect 50502 16624 50554 16676
rect 50566 16624 50618 16676
rect 5974 16513 6026 16565
rect 13558 16513 13610 16565
rect 30166 16513 30218 16565
rect 46870 16513 46922 16565
rect 7126 16439 7178 16491
rect 54070 16439 54122 16491
rect 52438 16069 52490 16121
rect 4294 15958 4346 16010
rect 4358 15958 4410 16010
rect 4422 15958 4474 16010
rect 4486 15958 4538 16010
rect 35014 15958 35066 16010
rect 35078 15958 35130 16010
rect 35142 15958 35194 16010
rect 35206 15958 35258 16010
rect 21430 15551 21482 15603
rect 36694 15477 36746 15529
rect 38902 15403 38954 15455
rect 19654 15292 19706 15344
rect 19718 15292 19770 15344
rect 19782 15292 19834 15344
rect 19846 15292 19898 15344
rect 50374 15292 50426 15344
rect 50438 15292 50490 15344
rect 50502 15292 50554 15344
rect 50566 15292 50618 15344
rect 13654 15181 13706 15233
rect 22198 15181 22250 15233
rect 58006 15076 58058 15085
rect 58006 15042 58015 15076
rect 58015 15042 58049 15076
rect 58049 15042 58058 15076
rect 58006 15033 58058 15042
rect 17782 14885 17834 14937
rect 46582 14885 46634 14937
rect 7702 14811 7754 14863
rect 4294 14626 4346 14678
rect 4358 14626 4410 14678
rect 4422 14626 4474 14678
rect 4486 14626 4538 14678
rect 35014 14626 35066 14678
rect 35078 14626 35130 14678
rect 35142 14626 35194 14678
rect 35206 14626 35258 14678
rect 45046 14515 45098 14567
rect 45238 14441 45290 14493
rect 17782 14410 17834 14419
rect 17782 14376 17791 14410
rect 17791 14376 17825 14410
rect 17825 14376 17834 14410
rect 17782 14367 17834 14376
rect 34102 14145 34154 14197
rect 4726 14114 4778 14123
rect 4726 14080 4735 14114
rect 4735 14080 4769 14114
rect 4769 14080 4778 14114
rect 4726 14071 4778 14080
rect 36790 14071 36842 14123
rect 19654 13960 19706 14012
rect 19718 13960 19770 14012
rect 19782 13960 19834 14012
rect 19846 13960 19898 14012
rect 50374 13960 50426 14012
rect 50438 13960 50490 14012
rect 50502 13960 50554 14012
rect 50566 13960 50618 14012
rect 4726 13849 4778 13901
rect 27478 13849 27530 13901
rect 9238 13701 9290 13753
rect 25654 13701 25706 13753
rect 7606 13627 7658 13679
rect 9910 13627 9962 13679
rect 32854 13627 32906 13679
rect 8374 13479 8426 13531
rect 29974 13479 30026 13531
rect 8566 13405 8618 13457
rect 9814 13405 9866 13457
rect 15094 13448 15146 13457
rect 15094 13414 15103 13448
rect 15103 13414 15137 13448
rect 15137 13414 15146 13448
rect 15094 13405 15146 13414
rect 51574 13701 51626 13753
rect 4294 13294 4346 13346
rect 4358 13294 4410 13346
rect 4422 13294 4474 13346
rect 4486 13294 4538 13346
rect 35014 13294 35066 13346
rect 35078 13294 35130 13346
rect 35142 13294 35194 13346
rect 35206 13294 35258 13346
rect 7606 13226 7658 13235
rect 7606 13192 7615 13226
rect 7615 13192 7649 13226
rect 7649 13192 7658 13226
rect 7606 13183 7658 13192
rect 15094 13183 15146 13235
rect 48310 13183 48362 13235
rect 8374 13109 8426 13161
rect 36214 13109 36266 13161
rect 34006 13035 34058 13087
rect 28150 12961 28202 13013
rect 9910 12739 9962 12791
rect 19654 12628 19706 12680
rect 19718 12628 19770 12680
rect 19782 12628 19834 12680
rect 19846 12628 19898 12680
rect 50374 12628 50426 12680
rect 50438 12628 50490 12680
rect 50502 12628 50554 12680
rect 50566 12628 50618 12680
rect 8566 12517 8618 12569
rect 29302 12517 29354 12569
rect 6838 12369 6890 12421
rect 13078 12369 13130 12421
rect 56950 12369 57002 12421
rect 8086 12295 8138 12347
rect 27190 12295 27242 12347
rect 5206 12147 5258 12199
rect 12502 12221 12554 12273
rect 12790 12221 12842 12273
rect 15862 12147 15914 12199
rect 47542 12221 47594 12273
rect 57526 12221 57578 12273
rect 42454 12147 42506 12199
rect 15190 12116 15242 12125
rect 15190 12082 15199 12116
rect 15199 12082 15233 12116
rect 15233 12082 15242 12116
rect 15190 12073 15242 12082
rect 18742 12116 18794 12125
rect 18742 12082 18751 12116
rect 18751 12082 18785 12116
rect 18785 12082 18794 12116
rect 18742 12073 18794 12082
rect 33526 12073 33578 12125
rect 4294 11962 4346 12014
rect 4358 11962 4410 12014
rect 4422 11962 4474 12014
rect 4486 11962 4538 12014
rect 35014 11962 35066 12014
rect 35078 11962 35130 12014
rect 35142 11962 35194 12014
rect 35206 11962 35258 12014
rect 1750 11894 1802 11903
rect 1750 11860 1759 11894
rect 1759 11860 1793 11894
rect 1793 11860 1802 11894
rect 1750 11851 1802 11860
rect 5206 11894 5258 11903
rect 5206 11860 5215 11894
rect 5215 11860 5249 11894
rect 5249 11860 5258 11894
rect 5206 11851 5258 11860
rect 8374 11851 8426 11903
rect 15190 11851 15242 11903
rect 42934 11851 42986 11903
rect 8566 11777 8618 11829
rect 8086 11703 8138 11755
rect 24310 11703 24362 11755
rect 40438 11629 40490 11681
rect 38518 11555 38570 11607
rect 52534 11555 52586 11607
rect 54646 11598 54698 11607
rect 54646 11564 54655 11598
rect 54655 11564 54689 11598
rect 54689 11564 54698 11598
rect 54646 11555 54698 11564
rect 58198 11555 58250 11607
rect 57142 11407 57194 11459
rect 19654 11296 19706 11348
rect 19718 11296 19770 11348
rect 19782 11296 19834 11348
rect 19846 11296 19898 11348
rect 50374 11296 50426 11348
rect 50438 11296 50490 11348
rect 50502 11296 50554 11348
rect 50566 11296 50618 11348
rect 8662 11185 8714 11237
rect 16054 11185 16106 11237
rect 21334 11037 21386 11089
rect 8086 10963 8138 11015
rect 24214 10963 24266 11015
rect 24502 10963 24554 11015
rect 33814 10963 33866 11015
rect 56086 11037 56138 11089
rect 10582 10815 10634 10867
rect 26806 10815 26858 10867
rect 28438 10815 28490 10867
rect 29590 10815 29642 10867
rect 56758 10889 56810 10941
rect 58294 10815 58346 10867
rect 10870 10741 10922 10793
rect 11158 10741 11210 10793
rect 36022 10741 36074 10793
rect 40726 10741 40778 10793
rect 50902 10741 50954 10793
rect 4294 10630 4346 10682
rect 4358 10630 4410 10682
rect 4422 10630 4474 10682
rect 4486 10630 4538 10682
rect 35014 10630 35066 10682
rect 35078 10630 35130 10682
rect 35142 10630 35194 10682
rect 35206 10630 35258 10682
rect 56854 10562 56906 10571
rect 56854 10528 56863 10562
rect 56863 10528 56897 10562
rect 56897 10528 56906 10562
rect 56854 10519 56906 10528
rect 10582 10445 10634 10497
rect 12886 10371 12938 10423
rect 25174 10297 25226 10349
rect 55990 10371 56042 10423
rect 56086 10371 56138 10423
rect 26614 10223 26666 10275
rect 51574 10223 51626 10275
rect 8086 10149 8138 10201
rect 16246 10149 16298 10201
rect 56854 10223 56906 10275
rect 9430 10075 9482 10127
rect 17110 10075 17162 10127
rect 55702 10075 55754 10127
rect 56470 10075 56522 10127
rect 58582 10075 58634 10127
rect 19654 9964 19706 10016
rect 19718 9964 19770 10016
rect 19782 9964 19834 10016
rect 19846 9964 19898 10016
rect 50374 9964 50426 10016
rect 50438 9964 50490 10016
rect 50502 9964 50554 10016
rect 50566 9964 50618 10016
rect 8086 9853 8138 9905
rect 17974 9853 18026 9905
rect 18358 9853 18410 9905
rect 21526 9853 21578 9905
rect 7990 9779 8042 9831
rect 10966 9779 11018 9831
rect 20374 9779 20426 9831
rect 42838 9853 42890 9905
rect 55126 9853 55178 9905
rect 21718 9779 21770 9831
rect 49174 9779 49226 9831
rect 51670 9779 51722 9831
rect 20854 9705 20906 9757
rect 54646 9705 54698 9757
rect 8278 9631 8330 9683
rect 16150 9631 16202 9683
rect 17302 9631 17354 9683
rect 44662 9631 44714 9683
rect 46966 9631 47018 9683
rect 57622 9674 57674 9683
rect 57622 9640 57631 9674
rect 57631 9640 57665 9674
rect 57665 9640 57674 9674
rect 57622 9631 57674 9640
rect 18262 9557 18314 9609
rect 28246 9557 28298 9609
rect 28342 9557 28394 9609
rect 29494 9557 29546 9609
rect 54262 9557 54314 9609
rect 15094 9483 15146 9535
rect 43606 9483 43658 9535
rect 7798 9409 7850 9461
rect 12214 9409 12266 9461
rect 16534 9409 16586 9461
rect 20662 9409 20714 9461
rect 25846 9452 25898 9461
rect 25846 9418 25855 9452
rect 25855 9418 25889 9452
rect 25889 9418 25898 9452
rect 25846 9409 25898 9418
rect 34486 9409 34538 9461
rect 35446 9409 35498 9461
rect 41782 9409 41834 9461
rect 47734 9409 47786 9461
rect 54934 9557 54986 9609
rect 4294 9298 4346 9350
rect 4358 9298 4410 9350
rect 4422 9298 4474 9350
rect 4486 9298 4538 9350
rect 35014 9298 35066 9350
rect 35078 9298 35130 9350
rect 35142 9298 35194 9350
rect 35206 9298 35258 9350
rect 7894 9187 7946 9239
rect 13942 9187 13994 9239
rect 32950 9187 33002 9239
rect 33046 9187 33098 9239
rect 51670 9187 51722 9239
rect 53014 9230 53066 9239
rect 53014 9196 53023 9230
rect 53023 9196 53057 9230
rect 53057 9196 53066 9230
rect 53014 9187 53066 9196
rect 55606 9230 55658 9239
rect 16438 9113 16490 9165
rect 26806 9113 26858 9165
rect 28726 9113 28778 9165
rect 36310 9113 36362 9165
rect 8518 9039 8570 9091
rect 10774 9039 10826 9091
rect 17686 9039 17738 9091
rect 21718 9039 21770 9091
rect 8086 8965 8138 9017
rect 8230 8965 8282 9017
rect 8950 8965 9002 9017
rect 19318 8965 19370 9017
rect 54550 9039 54602 9091
rect 55222 8965 55274 9017
rect 55606 9196 55615 9230
rect 55615 9196 55649 9230
rect 55649 9196 55658 9230
rect 55606 9187 55658 9196
rect 57238 9008 57290 9017
rect 12694 8891 12746 8943
rect 18454 8891 18506 8943
rect 44086 8891 44138 8943
rect 57238 8974 57247 9008
rect 57247 8974 57281 9008
rect 57281 8974 57290 9008
rect 57238 8965 57290 8974
rect 16246 8817 16298 8869
rect 18166 8817 18218 8869
rect 7606 8786 7658 8795
rect 7606 8752 7615 8786
rect 7615 8752 7649 8786
rect 7649 8752 7658 8786
rect 7606 8743 7658 8752
rect 8854 8743 8906 8795
rect 9046 8743 9098 8795
rect 23158 8817 23210 8869
rect 26902 8817 26954 8869
rect 20950 8743 21002 8795
rect 22294 8743 22346 8795
rect 26998 8743 27050 8795
rect 30166 8743 30218 8795
rect 57334 8891 57386 8943
rect 53878 8743 53930 8795
rect 19654 8632 19706 8684
rect 19718 8632 19770 8684
rect 19782 8632 19834 8684
rect 19846 8632 19898 8684
rect 50374 8632 50426 8684
rect 50438 8632 50490 8684
rect 50502 8632 50554 8684
rect 50566 8632 50618 8684
rect 1846 8521 1898 8573
rect 5398 8521 5450 8573
rect 7606 8521 7658 8573
rect 8854 8521 8906 8573
rect 9910 8521 9962 8573
rect 12598 8521 12650 8573
rect 12790 8521 12842 8573
rect 48598 8564 48650 8573
rect 48598 8530 48607 8564
rect 48607 8530 48641 8564
rect 48641 8530 48650 8564
rect 48598 8521 48650 8530
rect 4918 8447 4970 8499
rect 2518 8416 2570 8425
rect 2518 8382 2527 8416
rect 2527 8382 2561 8416
rect 2561 8382 2570 8416
rect 2518 8373 2570 8382
rect 5110 8373 5162 8425
rect 7222 8373 7274 8425
rect 7990 8373 8042 8425
rect 8086 8373 8138 8425
rect 9718 8373 9770 8425
rect 9910 8373 9962 8425
rect 11350 8416 11402 8425
rect 11350 8382 11359 8416
rect 11359 8382 11393 8416
rect 11393 8382 11402 8416
rect 11350 8373 11402 8382
rect 13558 8373 13610 8425
rect 16246 8416 16298 8425
rect 16246 8382 16255 8416
rect 16255 8382 16289 8416
rect 16289 8382 16298 8416
rect 16246 8373 16298 8382
rect 17014 8416 17066 8425
rect 17014 8382 17023 8416
rect 17023 8382 17057 8416
rect 17057 8382 17066 8416
rect 17014 8373 17066 8382
rect 1654 8268 1706 8277
rect 1654 8234 1663 8268
rect 1663 8234 1697 8268
rect 1697 8234 1706 8268
rect 1654 8225 1706 8234
rect 2134 8225 2186 8277
rect 3190 8268 3242 8277
rect 3190 8234 3199 8268
rect 3199 8234 3233 8268
rect 3233 8234 3242 8268
rect 3190 8225 3242 8234
rect 4822 8151 4874 8203
rect 6838 8225 6890 8277
rect 13750 8299 13802 8351
rect 48118 8416 48170 8425
rect 48118 8382 48127 8416
rect 48127 8382 48161 8416
rect 48161 8382 48170 8416
rect 48118 8373 48170 8382
rect 58966 8521 59018 8573
rect 49750 8416 49802 8425
rect 49750 8382 49759 8416
rect 49759 8382 49793 8416
rect 49793 8382 49802 8416
rect 49750 8373 49802 8382
rect 51574 8373 51626 8425
rect 53206 8416 53258 8425
rect 53206 8382 53215 8416
rect 53215 8382 53249 8416
rect 53249 8382 53258 8416
rect 53206 8373 53258 8382
rect 54070 8416 54122 8425
rect 54070 8382 54079 8416
rect 54079 8382 54113 8416
rect 54113 8382 54122 8416
rect 54070 8373 54122 8382
rect 7702 8225 7754 8277
rect 9526 8225 9578 8277
rect 10294 8225 10346 8277
rect 5494 8120 5546 8129
rect 5494 8086 5503 8120
rect 5503 8086 5537 8120
rect 5537 8086 5546 8120
rect 5494 8077 5546 8086
rect 10678 8225 10730 8277
rect 11446 8225 11498 8277
rect 12214 8225 12266 8277
rect 51190 8299 51242 8351
rect 16054 8225 16106 8277
rect 16342 8225 16394 8277
rect 48022 8151 48074 8203
rect 48694 8225 48746 8277
rect 49462 8225 49514 8277
rect 53110 8151 53162 8203
rect 53494 8225 53546 8277
rect 56950 8299 57002 8351
rect 58390 8225 58442 8277
rect 59830 8151 59882 8203
rect 16246 8077 16298 8129
rect 31222 8077 31274 8129
rect 44950 8077 45002 8129
rect 4294 7966 4346 8018
rect 4358 7966 4410 8018
rect 4422 7966 4474 8018
rect 4486 7966 4538 8018
rect 35014 7966 35066 8018
rect 35078 7966 35130 8018
rect 35142 7966 35194 8018
rect 35206 7966 35258 8018
rect 8518 7855 8570 7907
rect 11254 7855 11306 7907
rect 36502 7898 36554 7907
rect 36502 7864 36511 7898
rect 36511 7864 36545 7898
rect 36545 7864 36554 7898
rect 36502 7855 36554 7864
rect 41014 7855 41066 7907
rect 42262 7898 42314 7907
rect 42262 7864 42271 7898
rect 42271 7864 42305 7898
rect 42305 7864 42314 7898
rect 42262 7855 42314 7864
rect 45238 7898 45290 7907
rect 45238 7864 45247 7898
rect 45247 7864 45281 7898
rect 45281 7864 45290 7898
rect 45238 7855 45290 7864
rect 46198 7855 46250 7907
rect 47542 7898 47594 7907
rect 47542 7864 47551 7898
rect 47551 7864 47585 7898
rect 47585 7864 47594 7898
rect 48982 7898 49034 7907
rect 47542 7855 47594 7864
rect 48982 7864 48991 7898
rect 48991 7864 49025 7898
rect 49025 7864 49034 7898
rect 48982 7855 49034 7864
rect 52918 7855 52970 7907
rect 3766 7781 3818 7833
rect 7798 7781 7850 7833
rect 5494 7707 5546 7759
rect 7942 7707 7994 7759
rect 9142 7707 9194 7759
rect 11734 7707 11786 7759
rect 1462 7633 1514 7685
rect 4054 7676 4106 7685
rect 4054 7642 4063 7676
rect 4063 7642 4097 7676
rect 4097 7642 4106 7676
rect 4054 7633 4106 7642
rect 4918 7633 4970 7685
rect 8518 7633 8570 7685
rect 9430 7676 9482 7685
rect 9430 7642 9439 7676
rect 9439 7642 9473 7676
rect 9473 7642 9482 7676
rect 9430 7633 9482 7642
rect 12022 7633 12074 7685
rect 12502 7633 12554 7685
rect 15094 7676 15146 7685
rect 15094 7642 15103 7676
rect 15103 7642 15137 7676
rect 15137 7642 15146 7676
rect 15094 7633 15146 7642
rect 15862 7676 15914 7685
rect 15862 7642 15871 7676
rect 15871 7642 15905 7676
rect 15905 7642 15914 7676
rect 15862 7633 15914 7642
rect 20950 7750 21002 7759
rect 20950 7716 20959 7750
rect 20959 7716 20993 7750
rect 20993 7716 21002 7750
rect 20950 7707 21002 7716
rect 24022 7707 24074 7759
rect 25462 7750 25514 7759
rect 25462 7716 25471 7750
rect 25471 7716 25505 7750
rect 25505 7716 25514 7750
rect 25462 7707 25514 7716
rect 26230 7750 26282 7759
rect 26230 7716 26239 7750
rect 26239 7716 26273 7750
rect 26273 7716 26282 7750
rect 26230 7707 26282 7716
rect 26998 7750 27050 7759
rect 26998 7716 27007 7750
rect 27007 7716 27041 7750
rect 27041 7716 27050 7750
rect 26998 7707 27050 7716
rect 54166 7781 54218 7833
rect 28438 7707 28490 7759
rect 29398 7750 29450 7759
rect 29398 7716 29407 7750
rect 29407 7716 29441 7750
rect 29441 7716 29450 7750
rect 29398 7707 29450 7716
rect 29590 7707 29642 7759
rect 31222 7750 31274 7759
rect 31222 7716 31231 7750
rect 31231 7716 31265 7750
rect 31265 7716 31274 7750
rect 31222 7707 31274 7716
rect 34582 7750 34634 7759
rect 34582 7716 34591 7750
rect 34591 7716 34625 7750
rect 34625 7716 34634 7750
rect 34582 7707 34634 7716
rect 35350 7750 35402 7759
rect 35350 7716 35359 7750
rect 35359 7716 35393 7750
rect 35393 7716 35402 7750
rect 35350 7707 35402 7716
rect 36118 7750 36170 7759
rect 36118 7716 36127 7750
rect 36127 7716 36161 7750
rect 36161 7716 36170 7750
rect 36118 7707 36170 7716
rect 36502 7707 36554 7759
rect 40342 7750 40394 7759
rect 40342 7716 40351 7750
rect 40351 7716 40385 7750
rect 40385 7716 40394 7750
rect 40342 7707 40394 7716
rect 41878 7750 41930 7759
rect 30070 7676 30122 7685
rect 30070 7642 30079 7676
rect 30079 7642 30113 7676
rect 30113 7642 30122 7676
rect 30070 7633 30122 7642
rect 40246 7633 40298 7685
rect 41878 7716 41887 7750
rect 41887 7716 41921 7750
rect 41921 7716 41930 7750
rect 41878 7707 41930 7716
rect 42262 7707 42314 7759
rect 44086 7750 44138 7759
rect 44086 7716 44095 7750
rect 44095 7716 44129 7750
rect 44129 7716 44138 7750
rect 44086 7707 44138 7716
rect 44854 7750 44906 7759
rect 44854 7716 44863 7750
rect 44863 7716 44897 7750
rect 44897 7716 44906 7750
rect 44854 7707 44906 7716
rect 45046 7707 45098 7759
rect 45814 7707 45866 7759
rect 47158 7750 47210 7759
rect 47158 7716 47167 7750
rect 47167 7716 47201 7750
rect 47201 7716 47210 7750
rect 47158 7707 47210 7716
rect 47542 7707 47594 7759
rect 48406 7707 48458 7759
rect 51766 7750 51818 7759
rect 51766 7716 51775 7750
rect 51775 7716 51809 7750
rect 51809 7716 51818 7750
rect 51766 7707 51818 7716
rect 52630 7750 52682 7759
rect 52630 7716 52639 7750
rect 52639 7716 52673 7750
rect 52673 7716 52682 7750
rect 52630 7707 52682 7716
rect 52726 7707 52778 7759
rect 42166 7633 42218 7685
rect 5590 7602 5642 7611
rect 5590 7568 5599 7602
rect 5599 7568 5633 7602
rect 5633 7568 5642 7602
rect 5590 7559 5642 7568
rect 8086 7559 8138 7611
rect 12310 7559 12362 7611
rect 9910 7485 9962 7537
rect 21238 7559 21290 7611
rect 33910 7559 33962 7611
rect 34486 7559 34538 7611
rect 2422 7454 2474 7463
rect 2422 7420 2431 7454
rect 2431 7420 2465 7454
rect 2465 7420 2474 7454
rect 2422 7411 2474 7420
rect 2998 7411 3050 7463
rect 3958 7454 4010 7463
rect 3958 7420 3967 7454
rect 3967 7420 4001 7454
rect 4001 7420 4010 7454
rect 3958 7411 4010 7420
rect 4054 7411 4106 7463
rect 5302 7411 5354 7463
rect 9334 7454 9386 7463
rect 9334 7420 9343 7454
rect 9343 7420 9377 7454
rect 9377 7420 9386 7454
rect 9334 7411 9386 7420
rect 22966 7485 23018 7537
rect 36214 7485 36266 7537
rect 41014 7559 41066 7611
rect 45238 7559 45290 7611
rect 46198 7633 46250 7685
rect 48982 7633 49034 7685
rect 49654 7633 49706 7685
rect 52918 7633 52970 7685
rect 58774 7707 58826 7759
rect 55798 7676 55850 7685
rect 55798 7642 55807 7676
rect 55807 7642 55841 7676
rect 55841 7642 55850 7676
rect 55798 7633 55850 7642
rect 56182 7633 56234 7685
rect 56662 7633 56714 7685
rect 10966 7411 11018 7463
rect 12502 7411 12554 7463
rect 15670 7411 15722 7463
rect 15862 7411 15914 7463
rect 16150 7411 16202 7463
rect 20758 7411 20810 7463
rect 23830 7454 23882 7463
rect 23830 7420 23839 7454
rect 23839 7420 23873 7454
rect 23873 7420 23882 7454
rect 23830 7411 23882 7420
rect 24118 7411 24170 7463
rect 24790 7411 24842 7463
rect 25558 7411 25610 7463
rect 26710 7411 26762 7463
rect 28150 7411 28202 7463
rect 29206 7411 29258 7463
rect 31030 7411 31082 7463
rect 33622 7411 33674 7463
rect 34390 7411 34442 7463
rect 34774 7411 34826 7463
rect 35830 7411 35882 7463
rect 36694 7411 36746 7463
rect 38038 7411 38090 7463
rect 38806 7411 38858 7463
rect 39574 7411 39626 7463
rect 41398 7411 41450 7463
rect 42454 7411 42506 7463
rect 43894 7411 43946 7463
rect 44662 7411 44714 7463
rect 46486 7411 46538 7463
rect 47254 7411 47306 7463
rect 49078 7485 49130 7537
rect 51670 7411 51722 7463
rect 52342 7411 52394 7463
rect 59350 7411 59402 7463
rect 19654 7300 19706 7352
rect 19718 7300 19770 7352
rect 19782 7300 19834 7352
rect 19846 7300 19898 7352
rect 50374 7300 50426 7352
rect 50438 7300 50490 7352
rect 50502 7300 50554 7352
rect 50566 7300 50618 7352
rect 5590 7189 5642 7241
rect 25846 7189 25898 7241
rect 6550 7115 6602 7167
rect 10582 7115 10634 7167
rect 12406 7115 12458 7167
rect 20662 7115 20714 7167
rect 23926 7158 23978 7167
rect 6070 7084 6122 7093
rect 6070 7050 6079 7084
rect 6079 7050 6113 7084
rect 6113 7050 6122 7084
rect 6070 7041 6122 7050
rect 7126 7041 7178 7093
rect 15862 7084 15914 7093
rect 1654 7010 1706 7019
rect 1654 6976 1663 7010
rect 1663 6976 1697 7010
rect 1697 6976 1706 7010
rect 1654 6967 1706 6976
rect 2518 7010 2570 7019
rect 2518 6976 2527 7010
rect 2527 6976 2561 7010
rect 2561 6976 2570 7010
rect 2518 6967 2570 6976
rect 3670 6967 3722 7019
rect 6358 6967 6410 7019
rect 7030 6967 7082 7019
rect 7606 7010 7658 7019
rect 7606 6976 7615 7010
rect 7615 6976 7649 7010
rect 7649 6976 7658 7010
rect 7606 6967 7658 6976
rect 5878 6893 5930 6945
rect 6550 6893 6602 6945
rect 6934 6893 6986 6945
rect 8854 6967 8906 7019
rect 10582 7010 10634 7019
rect 7318 6819 7370 6871
rect 9238 6893 9290 6945
rect 5206 6745 5258 6797
rect 8086 6745 8138 6797
rect 9814 6936 9866 6945
rect 9814 6902 9823 6936
rect 9823 6902 9857 6936
rect 9857 6902 9866 6936
rect 10582 6976 10591 7010
rect 10591 6976 10625 7010
rect 10625 6976 10634 7010
rect 10582 6967 10634 6976
rect 9814 6893 9866 6902
rect 15862 7050 15871 7084
rect 15871 7050 15905 7084
rect 15905 7050 15914 7084
rect 15862 7041 15914 7050
rect 17302 7084 17354 7093
rect 17302 7050 17311 7084
rect 17311 7050 17345 7084
rect 17345 7050 17354 7084
rect 17302 7041 17354 7050
rect 18262 7041 18314 7093
rect 18934 7041 18986 7093
rect 20374 7084 20426 7093
rect 20374 7050 20383 7084
rect 20383 7050 20417 7084
rect 20417 7050 20426 7084
rect 20374 7041 20426 7050
rect 23926 7124 23935 7158
rect 23935 7124 23969 7158
rect 23969 7124 23978 7158
rect 26806 7158 26858 7167
rect 23926 7115 23978 7124
rect 21430 7041 21482 7093
rect 22678 7084 22730 7093
rect 22678 7050 22687 7084
rect 22687 7050 22721 7084
rect 22721 7050 22730 7084
rect 22678 7041 22730 7050
rect 26806 7124 26815 7158
rect 26815 7124 26849 7158
rect 26849 7124 26858 7158
rect 29110 7158 29162 7167
rect 26806 7115 26858 7124
rect 25750 7041 25802 7093
rect 26422 7084 26474 7093
rect 26422 7050 26431 7084
rect 26431 7050 26465 7084
rect 26465 7050 26474 7084
rect 26422 7041 26474 7050
rect 29110 7124 29119 7158
rect 29119 7124 29153 7158
rect 29153 7124 29162 7158
rect 36598 7158 36650 7167
rect 29110 7115 29162 7124
rect 28342 7041 28394 7093
rect 28726 7084 28778 7093
rect 28726 7050 28735 7084
rect 28735 7050 28769 7084
rect 28769 7050 28778 7084
rect 28726 7041 28778 7050
rect 36598 7124 36607 7158
rect 36607 7124 36641 7158
rect 36641 7124 36650 7158
rect 36598 7115 36650 7124
rect 30934 7084 30986 7093
rect 30934 7050 30943 7084
rect 30943 7050 30977 7084
rect 30977 7050 30986 7084
rect 30934 7041 30986 7050
rect 31702 7084 31754 7093
rect 31702 7050 31711 7084
rect 31711 7050 31745 7084
rect 31745 7050 31754 7084
rect 31702 7041 31754 7050
rect 32374 7084 32426 7093
rect 32374 7050 32383 7084
rect 32383 7050 32417 7084
rect 32417 7050 32426 7084
rect 32374 7041 32426 7050
rect 33238 7084 33290 7093
rect 33238 7050 33247 7084
rect 33247 7050 33281 7084
rect 33281 7050 33290 7084
rect 33238 7041 33290 7050
rect 33814 7041 33866 7093
rect 36022 7041 36074 7093
rect 37462 7158 37514 7167
rect 37462 7124 37471 7158
rect 37471 7124 37505 7158
rect 37505 7124 37514 7158
rect 39670 7158 39722 7167
rect 37462 7115 37514 7124
rect 39670 7124 39679 7158
rect 39679 7124 39713 7158
rect 39713 7124 39722 7158
rect 41110 7158 41162 7167
rect 39670 7115 39722 7124
rect 38518 7084 38570 7093
rect 38518 7050 38527 7084
rect 38527 7050 38561 7084
rect 38561 7050 38570 7084
rect 38518 7041 38570 7050
rect 39286 7084 39338 7093
rect 39286 7050 39295 7084
rect 39295 7050 39329 7084
rect 39329 7050 39338 7084
rect 39286 7041 39338 7050
rect 41110 7124 41119 7158
rect 41119 7124 41153 7158
rect 41153 7124 41162 7158
rect 41110 7115 41162 7124
rect 41782 7115 41834 7167
rect 43414 7158 43466 7167
rect 43414 7124 43423 7158
rect 43423 7124 43457 7158
rect 43457 7124 43466 7158
rect 43414 7115 43466 7124
rect 42934 7084 42986 7093
rect 42934 7050 42943 7084
rect 42943 7050 42977 7084
rect 42977 7050 42986 7084
rect 42934 7041 42986 7050
rect 45142 7115 45194 7167
rect 48886 7115 48938 7167
rect 46678 7084 46730 7093
rect 46678 7050 46687 7084
rect 46687 7050 46721 7084
rect 46721 7050 46730 7084
rect 46678 7041 46730 7050
rect 47638 7041 47690 7093
rect 48310 7084 48362 7093
rect 48310 7050 48319 7084
rect 48319 7050 48353 7084
rect 48353 7050 48362 7084
rect 48310 7041 48362 7050
rect 49846 7115 49898 7167
rect 50230 7084 50282 7093
rect 50230 7050 50239 7084
rect 50239 7050 50273 7084
rect 50273 7050 50282 7084
rect 50230 7041 50282 7050
rect 52054 7084 52106 7093
rect 52054 7050 52063 7084
rect 52063 7050 52097 7084
rect 52097 7050 52106 7084
rect 52054 7041 52106 7050
rect 11254 7010 11306 7019
rect 11254 6976 11263 7010
rect 11263 6976 11297 7010
rect 11297 6976 11306 7010
rect 11254 6967 11306 6976
rect 12694 7010 12746 7019
rect 12694 6976 12703 7010
rect 12703 6976 12737 7010
rect 12737 6976 12746 7010
rect 12694 6967 12746 6976
rect 12310 6893 12362 6945
rect 12886 6893 12938 6945
rect 13462 6893 13514 6945
rect 13750 6893 13802 6945
rect 14614 6893 14666 6945
rect 15382 6893 15434 6945
rect 17110 6893 17162 6945
rect 17878 6893 17930 6945
rect 18550 6893 18602 6945
rect 20374 6893 20426 6945
rect 20950 6893 21002 6945
rect 21238 6893 21290 6945
rect 22006 6893 22058 6945
rect 16246 6745 16298 6797
rect 25174 6967 25226 7019
rect 25942 6967 25994 7019
rect 23350 6936 23402 6945
rect 23350 6902 23359 6936
rect 23359 6902 23393 6936
rect 23393 6902 23402 6936
rect 23350 6893 23402 6902
rect 23926 6893 23978 6945
rect 24598 6893 24650 6945
rect 31414 6967 31466 7019
rect 25174 6819 25226 6871
rect 26998 6819 27050 6871
rect 29494 6936 29546 6945
rect 27766 6819 27818 6871
rect 29494 6902 29503 6936
rect 29503 6902 29537 6936
rect 29537 6902 29546 6936
rect 29494 6893 29546 6902
rect 29974 6893 30026 6945
rect 32566 6967 32618 7019
rect 30742 6819 30794 6871
rect 32182 6819 32234 6871
rect 26614 6745 26666 6797
rect 32950 6745 33002 6797
rect 35542 6893 35594 6945
rect 36406 6893 36458 6945
rect 37078 6893 37130 6945
rect 34006 6819 34058 6871
rect 37366 6819 37418 6871
rect 38518 6893 38570 6945
rect 41206 6967 41258 7019
rect 47830 6967 47882 7019
rect 54742 7010 54794 7019
rect 37654 6745 37706 6797
rect 39862 6819 39914 6871
rect 41302 6819 41354 6871
rect 42838 6819 42890 6871
rect 43606 6745 43658 6797
rect 44566 6819 44618 6871
rect 45430 6893 45482 6945
rect 47062 6893 47114 6945
rect 46870 6819 46922 6871
rect 48886 6893 48938 6945
rect 50134 6893 50186 6945
rect 51382 6893 51434 6945
rect 52822 6936 52874 6945
rect 52822 6902 52831 6936
rect 52831 6902 52865 6936
rect 52865 6902 52874 6936
rect 52822 6893 52874 6902
rect 54742 6976 54751 7010
rect 54751 6976 54785 7010
rect 54785 6976 54794 7010
rect 54742 6967 54794 6976
rect 55414 6967 55466 7019
rect 58486 6967 58538 7019
rect 56374 6893 56426 6945
rect 4294 6634 4346 6686
rect 4358 6634 4410 6686
rect 4422 6634 4474 6686
rect 4486 6634 4538 6686
rect 35014 6634 35066 6686
rect 35078 6634 35130 6686
rect 35142 6634 35194 6686
rect 35206 6634 35258 6686
rect 5398 6566 5450 6575
rect 5398 6532 5407 6566
rect 5407 6532 5441 6566
rect 5441 6532 5450 6566
rect 5398 6523 5450 6532
rect 8470 6523 8522 6575
rect 9334 6523 9386 6575
rect 15958 6566 16010 6575
rect 15958 6532 15967 6566
rect 15967 6532 16001 6566
rect 16001 6532 16010 6566
rect 30262 6566 30314 6575
rect 15958 6523 16010 6532
rect 9046 6449 9098 6501
rect 7126 6418 7178 6427
rect 7126 6384 7135 6418
rect 7135 6384 7169 6418
rect 7169 6384 7178 6418
rect 7126 6375 7178 6384
rect 7222 6375 7274 6427
rect 8374 6375 8426 6427
rect 13078 6375 13130 6427
rect 13942 6418 13994 6427
rect 13942 6384 13951 6418
rect 13951 6384 13985 6418
rect 13985 6384 13994 6418
rect 15478 6418 15530 6427
rect 13942 6375 13994 6384
rect 15478 6384 15487 6418
rect 15487 6384 15521 6418
rect 15521 6384 15530 6418
rect 15478 6375 15530 6384
rect 30262 6532 30271 6566
rect 30271 6532 30305 6566
rect 30305 6532 30314 6566
rect 31798 6566 31850 6575
rect 30262 6523 30314 6532
rect 17686 6418 17738 6427
rect 17686 6384 17695 6418
rect 17695 6384 17729 6418
rect 17729 6384 17738 6418
rect 17686 6375 17738 6384
rect 18454 6418 18506 6427
rect 18454 6384 18463 6418
rect 18463 6384 18497 6418
rect 18497 6384 18506 6418
rect 18454 6375 18506 6384
rect 19126 6418 19178 6427
rect 19126 6384 19135 6418
rect 19135 6384 19169 6418
rect 19169 6384 19178 6418
rect 19126 6375 19178 6384
rect 19990 6418 20042 6427
rect 19990 6384 19999 6418
rect 19999 6384 20033 6418
rect 20033 6384 20042 6418
rect 19990 6375 20042 6384
rect 20854 6375 20906 6427
rect 21526 6418 21578 6427
rect 21526 6384 21535 6418
rect 21535 6384 21569 6418
rect 21569 6384 21578 6418
rect 21526 6375 21578 6384
rect 23734 6418 23786 6427
rect 23734 6384 23743 6418
rect 23743 6384 23777 6418
rect 23777 6384 23786 6418
rect 23734 6375 23786 6384
rect 24502 6418 24554 6427
rect 24502 6384 24511 6418
rect 24511 6384 24545 6418
rect 24545 6384 24554 6418
rect 24502 6375 24554 6384
rect 28246 6418 28298 6427
rect 28246 6384 28255 6418
rect 28255 6384 28289 6418
rect 28289 6384 28298 6418
rect 28246 6375 28298 6384
rect 29014 6418 29066 6427
rect 29014 6384 29023 6418
rect 29023 6384 29057 6418
rect 29057 6384 29066 6418
rect 29014 6375 29066 6384
rect 31798 6532 31807 6566
rect 31807 6532 31841 6566
rect 31841 6532 31850 6566
rect 31798 6523 31850 6532
rect 30646 6375 30698 6427
rect 34870 6523 34922 6575
rect 36886 6566 36938 6575
rect 33526 6418 33578 6427
rect 33526 6384 33535 6418
rect 33535 6384 33569 6418
rect 33569 6384 33578 6418
rect 33526 6375 33578 6384
rect 34198 6418 34250 6427
rect 34198 6384 34207 6418
rect 34207 6384 34241 6418
rect 34241 6384 34250 6418
rect 34198 6375 34250 6384
rect 36886 6532 36895 6566
rect 36895 6532 36929 6566
rect 36929 6532 36938 6566
rect 51286 6566 51338 6575
rect 36886 6523 36938 6532
rect 51286 6532 51295 6566
rect 51295 6532 51329 6566
rect 51329 6532 51338 6566
rect 51286 6523 51338 6532
rect 47734 6449 47786 6501
rect 42742 6418 42794 6427
rect 42742 6384 42751 6418
rect 42751 6384 42785 6418
rect 42785 6384 42794 6418
rect 42742 6375 42794 6384
rect 44758 6375 44810 6427
rect 50902 6418 50954 6427
rect 50902 6384 50911 6418
rect 50911 6384 50945 6418
rect 50945 6384 50954 6418
rect 50902 6375 50954 6384
rect 52438 6418 52490 6427
rect 52438 6384 52447 6418
rect 52447 6384 52481 6418
rect 52481 6384 52490 6418
rect 52438 6375 52490 6384
rect 1558 6344 1610 6353
rect 1558 6310 1567 6344
rect 1567 6310 1601 6344
rect 1601 6310 1610 6344
rect 1558 6301 1610 6310
rect 2038 6301 2090 6353
rect 3190 6344 3242 6353
rect 3190 6310 3199 6344
rect 3199 6310 3233 6344
rect 3233 6310 3242 6344
rect 3190 6301 3242 6310
rect 3862 6301 3914 6353
rect 4630 6301 4682 6353
rect 9430 6344 9482 6353
rect 9430 6310 9439 6344
rect 9439 6310 9473 6344
rect 9473 6310 9482 6344
rect 9430 6301 9482 6310
rect 10102 6301 10154 6353
rect 10870 6301 10922 6353
rect 11638 6301 11690 6353
rect 12406 6301 12458 6353
rect 18742 6301 18794 6353
rect 25654 6344 25706 6353
rect 25654 6310 25663 6344
rect 25663 6310 25697 6344
rect 25697 6310 25706 6344
rect 25654 6301 25706 6310
rect 26806 6344 26858 6353
rect 26806 6310 26815 6344
rect 26815 6310 26849 6344
rect 26849 6310 26858 6344
rect 26806 6301 26858 6310
rect 29686 6344 29738 6353
rect 29686 6310 29695 6344
rect 29695 6310 29729 6344
rect 29729 6310 29738 6344
rect 29686 6301 29738 6310
rect 31222 6344 31274 6353
rect 31222 6310 31231 6344
rect 31231 6310 31265 6344
rect 31265 6310 31274 6344
rect 31222 6301 31274 6310
rect 36310 6344 36362 6353
rect 36310 6310 36319 6344
rect 36319 6310 36353 6344
rect 36353 6310 36362 6344
rect 36310 6301 36362 6310
rect 38902 6344 38954 6353
rect 38902 6310 38911 6344
rect 38911 6310 38945 6344
rect 38945 6310 38954 6344
rect 38902 6301 38954 6310
rect 40342 6344 40394 6353
rect 40342 6310 40351 6344
rect 40351 6310 40385 6344
rect 40385 6310 40394 6344
rect 40342 6301 40394 6310
rect 41878 6344 41930 6353
rect 41878 6310 41887 6344
rect 41887 6310 41921 6344
rect 41921 6310 41930 6344
rect 41878 6301 41930 6310
rect 45526 6344 45578 6353
rect 45526 6310 45535 6344
rect 45535 6310 45569 6344
rect 45569 6310 45578 6344
rect 45526 6301 45578 6310
rect 46966 6344 47018 6353
rect 46966 6310 46975 6344
rect 46975 6310 47009 6344
rect 47009 6310 47018 6344
rect 46966 6301 47018 6310
rect 47734 6344 47786 6353
rect 47734 6310 47743 6344
rect 47743 6310 47777 6344
rect 47777 6310 47786 6344
rect 47734 6301 47786 6310
rect 48790 6301 48842 6353
rect 49558 6301 49610 6353
rect 56854 6375 56906 6427
rect 53974 6301 54026 6353
rect 15766 6227 15818 6279
rect 43798 6227 43850 6279
rect 44086 6270 44138 6279
rect 44086 6236 44095 6270
rect 44095 6236 44129 6270
rect 44129 6236 44138 6270
rect 44086 6227 44138 6236
rect 54358 6227 54410 6279
rect 14230 6153 14282 6205
rect 5494 6079 5546 6131
rect 6262 6079 6314 6131
rect 14518 6079 14570 6131
rect 18934 6153 18986 6205
rect 16534 6079 16586 6131
rect 17590 6122 17642 6131
rect 17590 6088 17599 6122
rect 17599 6088 17633 6122
rect 17633 6088 17642 6122
rect 17590 6079 17642 6088
rect 18262 6079 18314 6131
rect 19318 6079 19370 6131
rect 20086 6153 20138 6205
rect 20662 6122 20714 6131
rect 20662 6088 20671 6122
rect 20671 6088 20705 6122
rect 20705 6088 20714 6122
rect 20662 6079 20714 6088
rect 22294 6153 22346 6205
rect 21526 6079 21578 6131
rect 31798 6153 31850 6205
rect 24022 6079 24074 6131
rect 26326 6079 26378 6131
rect 29014 6079 29066 6131
rect 29782 6079 29834 6131
rect 33718 6153 33770 6205
rect 34294 6122 34346 6131
rect 34294 6088 34303 6122
rect 34303 6088 34337 6122
rect 34337 6088 34346 6122
rect 34294 6079 34346 6088
rect 40630 6153 40682 6205
rect 37270 6079 37322 6131
rect 39190 6079 39242 6131
rect 42166 6153 42218 6205
rect 51574 6153 51626 6205
rect 44182 6079 44234 6131
rect 49750 6079 49802 6131
rect 51094 6079 51146 6131
rect 55030 6153 55082 6205
rect 58102 6301 58154 6353
rect 58870 6227 58922 6279
rect 19654 5968 19706 6020
rect 19718 5968 19770 6020
rect 19782 5968 19834 6020
rect 19846 5968 19898 6020
rect 50374 5968 50426 6020
rect 50438 5968 50490 6020
rect 50502 5968 50554 6020
rect 50566 5968 50618 6020
rect 3574 5857 3626 5909
rect 7798 5857 7850 5909
rect 44086 5857 44138 5909
rect 49270 5857 49322 5909
rect 49654 5857 49706 5909
rect 7030 5709 7082 5761
rect 44950 5709 45002 5761
rect 1078 5635 1130 5687
rect 2902 5678 2954 5687
rect 2902 5644 2911 5678
rect 2911 5644 2945 5678
rect 2945 5644 2954 5678
rect 2902 5635 2954 5644
rect 4918 5635 4970 5687
rect 5110 5678 5162 5687
rect 5110 5644 5119 5678
rect 5119 5644 5153 5678
rect 5153 5644 5162 5678
rect 5110 5635 5162 5644
rect 5782 5635 5834 5687
rect 6838 5678 6890 5687
rect 6838 5644 6847 5678
rect 6847 5644 6881 5678
rect 6881 5644 6890 5678
rect 6838 5635 6890 5644
rect 7222 5635 7274 5687
rect 8758 5635 8810 5687
rect 10198 5635 10250 5687
rect 10486 5635 10538 5687
rect 12598 5678 12650 5687
rect 12598 5644 12607 5678
rect 12607 5644 12641 5678
rect 12641 5644 12650 5678
rect 12598 5635 12650 5644
rect 13366 5678 13418 5687
rect 13366 5644 13375 5678
rect 13375 5644 13409 5678
rect 13409 5644 13418 5678
rect 13366 5635 13418 5644
rect 14998 5678 15050 5687
rect 14998 5644 15007 5678
rect 15007 5644 15041 5678
rect 15041 5644 15050 5678
rect 14998 5635 15050 5644
rect 15862 5678 15914 5687
rect 15862 5644 15871 5678
rect 15871 5644 15905 5678
rect 15905 5644 15914 5678
rect 15862 5635 15914 5644
rect 16150 5635 16202 5687
rect 17302 5678 17354 5687
rect 17302 5644 17311 5678
rect 17311 5644 17345 5678
rect 17345 5644 17354 5678
rect 18742 5678 18794 5687
rect 17302 5635 17354 5644
rect 18742 5644 18751 5678
rect 18751 5644 18785 5678
rect 18785 5644 18794 5678
rect 18742 5635 18794 5644
rect 20182 5678 20234 5687
rect 20182 5644 20191 5678
rect 20191 5644 20225 5678
rect 20225 5644 20234 5678
rect 20182 5635 20234 5644
rect 20566 5635 20618 5687
rect 21814 5635 21866 5687
rect 23062 5635 23114 5687
rect 23446 5635 23498 5687
rect 24598 5635 24650 5687
rect 26230 5678 26282 5687
rect 26230 5644 26239 5678
rect 26239 5644 26273 5678
rect 26273 5644 26282 5678
rect 26230 5635 26282 5644
rect 27382 5635 27434 5687
rect 27862 5635 27914 5687
rect 28822 5635 28874 5687
rect 30262 5635 30314 5687
rect 30838 5635 30890 5687
rect 31702 5635 31754 5687
rect 33142 5678 33194 5687
rect 33142 5644 33151 5678
rect 33151 5644 33185 5678
rect 33185 5644 33194 5678
rect 33142 5635 33194 5644
rect 33238 5635 33290 5687
rect 34678 5678 34730 5687
rect 34678 5644 34687 5678
rect 34687 5644 34721 5678
rect 34721 5644 34730 5678
rect 34678 5635 34730 5644
rect 36022 5678 36074 5687
rect 36022 5644 36031 5678
rect 36031 5644 36065 5678
rect 36065 5644 36074 5678
rect 36022 5635 36074 5644
rect 36214 5635 36266 5687
rect 37558 5678 37610 5687
rect 37558 5644 37567 5678
rect 37567 5644 37601 5678
rect 37601 5644 37610 5678
rect 37558 5635 37610 5644
rect 39094 5678 39146 5687
rect 39094 5644 39103 5678
rect 39103 5644 39137 5678
rect 39137 5644 39146 5678
rect 39094 5635 39146 5644
rect 39286 5635 39338 5687
rect 40726 5635 40778 5687
rect 41782 5635 41834 5687
rect 42262 5635 42314 5687
rect 43222 5635 43274 5687
rect 43702 5635 43754 5687
rect 45142 5678 45194 5687
rect 45142 5644 45151 5678
rect 45151 5644 45185 5678
rect 45185 5644 45194 5678
rect 45142 5635 45194 5644
rect 46102 5635 46154 5687
rect 46678 5635 46730 5687
rect 47542 5635 47594 5687
rect 48982 5678 49034 5687
rect 48982 5644 48991 5678
rect 48991 5644 49025 5678
rect 49025 5644 49034 5678
rect 48982 5635 49034 5644
rect 49654 5678 49706 5687
rect 49654 5644 49663 5678
rect 49663 5644 49697 5678
rect 49697 5644 49706 5678
rect 49654 5635 49706 5644
rect 50710 5635 50762 5687
rect 52150 5678 52202 5687
rect 52150 5644 52159 5678
rect 52159 5644 52193 5678
rect 52193 5644 52202 5678
rect 52150 5635 52202 5644
rect 52534 5635 52586 5687
rect 53686 5678 53738 5687
rect 53686 5644 53695 5678
rect 53695 5644 53729 5678
rect 53729 5644 53738 5678
rect 53686 5635 53738 5644
rect 57430 5678 57482 5687
rect 46294 5561 46346 5613
rect 53590 5561 53642 5613
rect 57430 5644 57439 5678
rect 57439 5644 57473 5678
rect 57473 5644 57482 5678
rect 57430 5635 57482 5644
rect 59638 5561 59690 5613
rect 7606 5487 7658 5539
rect 21718 5487 21770 5539
rect 26038 5487 26090 5539
rect 37462 5487 37514 5539
rect 3766 5413 3818 5465
rect 8374 5413 8426 5465
rect 4294 5302 4346 5354
rect 4358 5302 4410 5354
rect 4422 5302 4474 5354
rect 4486 5302 4538 5354
rect 35014 5302 35066 5354
rect 35078 5302 35130 5354
rect 35142 5302 35194 5354
rect 35206 5302 35258 5354
rect 5014 5191 5066 5243
rect 310 4969 362 5021
rect 1846 4969 1898 5021
rect 3094 5012 3146 5021
rect 3094 4978 3103 5012
rect 3103 4978 3137 5012
rect 3137 4978 3146 5012
rect 3094 4969 3146 4978
rect 4150 5012 4202 5021
rect 4150 4978 4159 5012
rect 4159 4978 4193 5012
rect 4193 4978 4202 5012
rect 4150 4969 4202 4978
rect 5398 5012 5450 5021
rect 5398 4978 5407 5012
rect 5407 4978 5441 5012
rect 5441 4978 5450 5012
rect 5398 4969 5450 4978
rect 6070 4969 6122 5021
rect 9238 5012 9290 5021
rect 9238 4978 9247 5012
rect 9247 4978 9281 5012
rect 9281 4978 9290 5012
rect 9238 4969 9290 4978
rect 10006 5012 10058 5021
rect 10006 4978 10015 5012
rect 10015 4978 10049 5012
rect 10049 4978 10058 5012
rect 10006 4969 10058 4978
rect 10582 4969 10634 5021
rect 11830 4969 11882 5021
rect 12982 5012 13034 5021
rect 12982 4978 12991 5012
rect 12991 4978 13025 5012
rect 13025 4978 13034 5012
rect 12982 4969 13034 4978
rect 13942 5012 13994 5021
rect 13942 4978 13951 5012
rect 13951 4978 13985 5012
rect 13985 4978 13994 5012
rect 13942 4969 13994 4978
rect 14422 4969 14474 5021
rect 14806 4969 14858 5021
rect 16438 4969 16490 5021
rect 17494 5012 17546 5021
rect 17494 4978 17503 5012
rect 17503 4978 17537 5012
rect 17537 4978 17546 5012
rect 17494 4969 17546 4978
rect 17974 4969 18026 5021
rect 19030 5012 19082 5021
rect 19030 4978 19039 5012
rect 19039 4978 19073 5012
rect 19073 4978 19082 5012
rect 19030 4969 19082 4978
rect 19126 4969 19178 5021
rect 20470 4969 20522 5021
rect 21238 4969 21290 5021
rect 22774 5012 22826 5021
rect 22774 4978 22783 5012
rect 22783 4978 22817 5012
rect 22817 4978 22826 5012
rect 22774 4969 22826 4978
rect 23542 5012 23594 5021
rect 23542 4978 23551 5012
rect 23551 4978 23585 5012
rect 23585 4978 23594 5012
rect 23542 4969 23594 4978
rect 25078 5012 25130 5021
rect 7942 4895 7994 4947
rect 23158 4895 23210 4947
rect 25078 4978 25087 5012
rect 25087 4978 25121 5012
rect 25121 4978 25130 5012
rect 25078 4969 25130 4978
rect 25846 5012 25898 5021
rect 25846 4978 25855 5012
rect 25855 4978 25889 5012
rect 25889 4978 25898 5012
rect 25846 4969 25898 4978
rect 26614 5012 26666 5021
rect 26614 4978 26623 5012
rect 26623 4978 26657 5012
rect 26657 4978 26666 5012
rect 26614 4969 26666 4978
rect 28054 5012 28106 5021
rect 28054 4978 28063 5012
rect 28063 4978 28097 5012
rect 28097 4978 28106 5012
rect 28054 4969 28106 4978
rect 28918 5012 28970 5021
rect 28918 4978 28927 5012
rect 28927 4978 28961 5012
rect 28961 4978 28970 5012
rect 28918 4969 28970 4978
rect 29302 4969 29354 5021
rect 30358 5012 30410 5021
rect 30358 4978 30367 5012
rect 30367 4978 30401 5012
rect 30401 4978 30410 5012
rect 30358 4969 30410 4978
rect 31126 5012 31178 5021
rect 31126 4978 31135 5012
rect 31135 4978 31169 5012
rect 31169 4978 31178 5012
rect 31126 4969 31178 4978
rect 31894 5012 31946 5021
rect 31894 4978 31903 5012
rect 31903 4978 31937 5012
rect 31937 4978 31946 5012
rect 31894 4969 31946 4978
rect 33334 5012 33386 5021
rect 33334 4978 33343 5012
rect 33343 4978 33377 5012
rect 33377 4978 33386 5012
rect 33334 4969 33386 4978
rect 34102 5012 34154 5021
rect 34102 4978 34111 5012
rect 34111 4978 34145 5012
rect 34145 4978 34154 5012
rect 34102 4969 34154 4978
rect 34870 5012 34922 5021
rect 34870 4978 34879 5012
rect 34879 4978 34913 5012
rect 34913 4978 34922 5012
rect 34870 4969 34922 4978
rect 34582 4895 34634 4947
rect 36118 4969 36170 5021
rect 36886 4969 36938 5021
rect 38614 5012 38666 5021
rect 38614 4978 38623 5012
rect 38623 4978 38657 5012
rect 38657 4978 38666 5012
rect 38614 4969 38666 4978
rect 39382 5012 39434 5021
rect 39382 4978 39391 5012
rect 39391 4978 39425 5012
rect 39425 4978 39434 5012
rect 39382 4969 39434 4978
rect 40150 5012 40202 5021
rect 40150 4978 40159 5012
rect 40159 4978 40193 5012
rect 40193 4978 40202 5012
rect 40150 4969 40202 4978
rect 40918 5012 40970 5021
rect 40918 4978 40927 5012
rect 40927 4978 40961 5012
rect 40961 4978 40970 5012
rect 40918 4969 40970 4978
rect 41686 5012 41738 5021
rect 41686 4978 41695 5012
rect 41695 4978 41729 5012
rect 41729 4978 41738 5012
rect 41686 4969 41738 4978
rect 42070 4969 42122 5021
rect 43318 4969 43370 5021
rect 44758 5012 44810 5021
rect 44758 4978 44767 5012
rect 44767 4978 44801 5012
rect 44801 4978 44810 5012
rect 44758 4969 44810 4978
rect 45430 5012 45482 5021
rect 45430 4978 45439 5012
rect 45439 4978 45473 5012
rect 45473 4978 45482 5012
rect 45430 4969 45482 4978
rect 46198 5012 46250 5021
rect 46198 4978 46207 5012
rect 46207 4978 46241 5012
rect 46241 4978 46250 5012
rect 46198 4969 46250 4978
rect 46294 4969 46346 5021
rect 47638 4969 47690 5021
rect 49366 5012 49418 5021
rect 49366 4978 49375 5012
rect 49375 4978 49409 5012
rect 49409 4978 49418 5012
rect 49366 4969 49418 4978
rect 50422 5012 50474 5021
rect 50422 4978 50431 5012
rect 50431 4978 50465 5012
rect 50465 4978 50474 5012
rect 50422 4969 50474 4978
rect 50902 4969 50954 5021
rect 51862 5012 51914 5021
rect 51862 4978 51871 5012
rect 51871 4978 51905 5012
rect 51905 4978 51914 5012
rect 51862 4969 51914 4978
rect 52246 4969 52298 5021
rect 53302 4969 53354 5021
rect 57046 5012 57098 5021
rect 8374 4821 8426 4873
rect 57046 4978 57055 5012
rect 57055 4978 57089 5012
rect 57089 4978 57098 5012
rect 57046 4969 57098 4978
rect 57814 4895 57866 4947
rect 59254 4821 59306 4873
rect 19654 4636 19706 4688
rect 19718 4636 19770 4688
rect 19782 4636 19834 4688
rect 19846 4636 19898 4688
rect 50374 4636 50426 4688
rect 50438 4636 50490 4688
rect 50502 4636 50554 4688
rect 50566 4636 50618 4688
rect 7894 4525 7946 4577
rect 9238 4525 9290 4577
rect 11158 4525 11210 4577
rect 12118 4451 12170 4503
rect 33910 4451 33962 4503
rect 35350 4451 35402 4503
rect 790 4377 842 4429
rect 1174 4303 1226 4355
rect 11062 4377 11114 4429
rect 15094 4377 15146 4429
rect 1366 4229 1418 4281
rect 3766 4229 3818 4281
rect 4726 4303 4778 4355
rect 5014 4229 5066 4281
rect 7414 4346 7466 4355
rect 5686 4229 5738 4281
rect 7414 4312 7423 4346
rect 7423 4312 7457 4346
rect 7457 4312 7466 4346
rect 7414 4303 7466 4312
rect 9622 4346 9674 4355
rect 3478 4155 3530 4207
rect 4918 4155 4970 4207
rect 6454 4155 6506 4207
rect 9622 4312 9631 4346
rect 9631 4312 9665 4346
rect 9665 4312 9674 4346
rect 9622 4303 9674 4312
rect 10390 4346 10442 4355
rect 10390 4312 10399 4346
rect 10399 4312 10433 4346
rect 10433 4312 10442 4346
rect 10390 4303 10442 4312
rect 10774 4303 10826 4355
rect 9814 4229 9866 4281
rect 10198 4229 10250 4281
rect 11158 4155 11210 4207
rect 13558 4346 13610 4355
rect 11446 4229 11498 4281
rect 13558 4312 13567 4346
rect 13567 4312 13601 4346
rect 13601 4312 13610 4346
rect 13558 4303 13610 4312
rect 15478 4346 15530 4355
rect 15478 4312 15487 4346
rect 15487 4312 15521 4346
rect 15521 4312 15530 4346
rect 15478 4303 15530 4312
rect 15958 4303 16010 4355
rect 14902 4229 14954 4281
rect 16534 4229 16586 4281
rect 16246 4155 16298 4207
rect 20278 4346 20330 4355
rect 16918 4081 16970 4133
rect 17686 4229 17738 4281
rect 20278 4312 20287 4346
rect 20287 4312 20321 4346
rect 20321 4312 20330 4346
rect 20278 4303 20330 4312
rect 21046 4346 21098 4355
rect 21046 4312 21055 4346
rect 21055 4312 21089 4346
rect 21089 4312 21098 4346
rect 21046 4303 21098 4312
rect 21814 4346 21866 4355
rect 21814 4312 21823 4346
rect 21823 4312 21857 4346
rect 21857 4312 21866 4346
rect 21814 4303 21866 4312
rect 23254 4346 23306 4355
rect 23254 4312 23263 4346
rect 23263 4312 23297 4346
rect 23297 4312 23306 4346
rect 23254 4303 23306 4312
rect 25462 4346 25514 4355
rect 22006 4229 22058 4281
rect 25462 4312 25471 4346
rect 25471 4312 25505 4346
rect 25505 4312 25514 4346
rect 25462 4303 25514 4312
rect 26134 4303 26186 4355
rect 26518 4303 26570 4355
rect 28342 4346 28394 4355
rect 28342 4312 28351 4346
rect 28351 4312 28385 4346
rect 28385 4312 28394 4346
rect 28342 4303 28394 4312
rect 29110 4346 29162 4355
rect 29110 4312 29119 4346
rect 29119 4312 29153 4346
rect 29153 4312 29162 4346
rect 29110 4303 29162 4312
rect 30934 4346 30986 4355
rect 30934 4312 30943 4346
rect 30943 4312 30977 4346
rect 30977 4312 30986 4346
rect 30934 4303 30986 4312
rect 31702 4346 31754 4355
rect 31702 4312 31711 4346
rect 31711 4312 31745 4346
rect 31745 4312 31754 4346
rect 31702 4303 31754 4312
rect 32758 4346 32810 4355
rect 32758 4312 32767 4346
rect 32767 4312 32801 4346
rect 32801 4312 32810 4346
rect 32758 4303 32810 4312
rect 33910 4346 33962 4355
rect 33910 4312 33919 4346
rect 33919 4312 33953 4346
rect 33953 4312 33962 4346
rect 33910 4303 33962 4312
rect 34582 4303 34634 4355
rect 34198 4229 34250 4281
rect 36790 4346 36842 4355
rect 36790 4312 36799 4346
rect 36799 4312 36833 4346
rect 36833 4312 36842 4346
rect 36790 4303 36842 4312
rect 37174 4229 37226 4281
rect 38998 4346 39050 4355
rect 38998 4312 39007 4346
rect 39007 4312 39041 4346
rect 39041 4312 39050 4346
rect 38998 4303 39050 4312
rect 39766 4346 39818 4355
rect 39766 4312 39775 4346
rect 39775 4312 39809 4346
rect 39809 4312 39818 4346
rect 39766 4303 39818 4312
rect 41974 4346 42026 4355
rect 41974 4312 41983 4346
rect 41983 4312 42017 4346
rect 42017 4312 42026 4346
rect 41974 4303 42026 4312
rect 42358 4303 42410 4355
rect 43414 4303 43466 4355
rect 44950 4346 45002 4355
rect 44950 4312 44959 4346
rect 44959 4312 44993 4346
rect 44993 4312 45002 4346
rect 44950 4303 45002 4312
rect 46774 4346 46826 4355
rect 46774 4312 46783 4346
rect 46783 4312 46817 4346
rect 46817 4312 46826 4346
rect 46774 4303 46826 4312
rect 43798 4229 43850 4281
rect 47446 4229 47498 4281
rect 47830 4303 47882 4355
rect 49846 4346 49898 4355
rect 48598 4229 48650 4281
rect 49846 4312 49855 4346
rect 49855 4312 49889 4346
rect 49889 4312 49898 4346
rect 49846 4303 49898 4312
rect 52630 4346 52682 4355
rect 49942 4229 49994 4281
rect 50998 4229 51050 4281
rect 52630 4312 52639 4346
rect 52639 4312 52673 4346
rect 52673 4312 52682 4346
rect 52630 4303 52682 4312
rect 53014 4229 53066 4281
rect 54070 4303 54122 4355
rect 55606 4346 55658 4355
rect 55606 4312 55615 4346
rect 55615 4312 55649 4346
rect 55649 4312 55658 4346
rect 55606 4303 55658 4312
rect 56662 4303 56714 4355
rect 57334 4229 57386 4281
rect 59158 4229 59210 4281
rect 27478 4155 27530 4207
rect 29014 4155 29066 4207
rect 38518 4155 38570 4207
rect 40150 4155 40202 4207
rect 55222 4155 55274 4207
rect 57910 4155 57962 4207
rect 17206 4081 17258 4133
rect 4294 3970 4346 4022
rect 4358 3970 4410 4022
rect 4422 3970 4474 4022
rect 4486 3970 4538 4022
rect 35014 3970 35066 4022
rect 35078 3970 35130 4022
rect 35142 3970 35194 4022
rect 35206 3970 35258 4022
rect 1942 3859 1994 3911
rect 2998 3859 3050 3911
rect 9046 3859 9098 3911
rect 10582 3859 10634 3911
rect 12310 3859 12362 3911
rect 13174 3859 13226 3911
rect 14134 3859 14186 3911
rect 15766 3859 15818 3911
rect 17206 3859 17258 3911
rect 17782 3859 17834 3911
rect 21334 3859 21386 3911
rect 22774 3859 22826 3911
rect 28534 3859 28586 3911
rect 29494 3859 29546 3911
rect 32566 3859 32618 3911
rect 34294 3859 34346 3911
rect 502 3785 554 3837
rect 1654 3785 1706 3837
rect 2326 3785 2378 3837
rect 3094 3785 3146 3837
rect 8278 3785 8330 3837
rect 10006 3785 10058 3837
rect 16534 3785 16586 3837
rect 17302 3785 17354 3837
rect 19414 3785 19466 3837
rect 20662 3785 20714 3837
rect 24214 3785 24266 3837
rect 25846 3785 25898 3837
rect 26422 3785 26474 3837
rect 28054 3785 28106 3837
rect 29014 3785 29066 3837
rect 30358 3785 30410 3837
rect 33430 3785 33482 3837
rect 34870 3785 34922 3837
rect 982 3711 1034 3763
rect 2422 3711 2474 3763
rect 2998 3711 3050 3763
rect 3286 3711 3338 3763
rect 3382 3711 3434 3763
rect 598 3637 650 3689
rect 1462 3637 1514 3689
rect 118 3563 170 3615
rect 1654 3637 1706 3689
rect 2710 3637 2762 3689
rect 3574 3637 3626 3689
rect 8758 3711 8810 3763
rect 38710 3859 38762 3911
rect 40054 3859 40106 3911
rect 41686 3859 41738 3911
rect 37846 3785 37898 3837
rect 39382 3785 39434 3837
rect 49174 3785 49226 3837
rect 50710 3785 50762 3837
rect 44566 3711 44618 3763
rect 5590 3680 5642 3689
rect 5590 3646 5599 3680
rect 5599 3646 5633 3680
rect 5633 3646 5642 3680
rect 5590 3637 5642 3646
rect 6358 3637 6410 3689
rect 7030 3637 7082 3689
rect 7798 3637 7850 3689
rect 8566 3637 8618 3689
rect 9334 3637 9386 3689
rect 1462 3489 1514 3541
rect 2134 3489 2186 3541
rect 2422 3415 2474 3467
rect 5206 3563 5258 3615
rect 10006 3489 10058 3541
rect 13174 3637 13226 3689
rect 13654 3680 13706 3689
rect 13654 3646 13663 3680
rect 13663 3646 13697 3680
rect 13697 3646 13706 3680
rect 13654 3637 13706 3646
rect 14134 3637 14186 3689
rect 14806 3637 14858 3689
rect 15286 3637 15338 3689
rect 17398 3637 17450 3689
rect 18166 3637 18218 3689
rect 18454 3637 18506 3689
rect 19222 3637 19274 3689
rect 19990 3637 20042 3689
rect 20662 3637 20714 3689
rect 22102 3637 22154 3689
rect 22870 3637 22922 3689
rect 23638 3637 23690 3689
rect 24406 3637 24458 3689
rect 24694 3563 24746 3615
rect 17302 3489 17354 3541
rect 17494 3489 17546 3541
rect 22582 3489 22634 3541
rect 23350 3489 23402 3541
rect 25846 3489 25898 3541
rect 27286 3637 27338 3689
rect 28054 3489 28106 3541
rect 3286 3415 3338 3467
rect 3958 3415 4010 3467
rect 12022 3415 12074 3467
rect 13366 3415 13418 3467
rect 22966 3415 23018 3467
rect 24022 3415 24074 3467
rect 28726 3415 28778 3467
rect 29878 3637 29930 3689
rect 30454 3637 30506 3689
rect 31318 3637 31370 3689
rect 32470 3637 32522 3689
rect 33526 3637 33578 3689
rect 34294 3637 34346 3689
rect 34966 3637 35018 3689
rect 35734 3637 35786 3689
rect 36502 3637 36554 3689
rect 37942 3637 37994 3689
rect 38710 3637 38762 3689
rect 39382 3489 39434 3541
rect 40150 3489 40202 3541
rect 41014 3637 41066 3689
rect 41590 3563 41642 3615
rect 42742 3637 42794 3689
rect 55894 3711 55946 3763
rect 43798 3563 43850 3615
rect 45238 3563 45290 3615
rect 41206 3489 41258 3541
rect 41686 3489 41738 3541
rect 46006 3489 46058 3541
rect 47158 3637 47210 3689
rect 48214 3637 48266 3689
rect 50710 3637 50762 3689
rect 50806 3637 50858 3689
rect 51286 3637 51338 3689
rect 52054 3637 52106 3689
rect 53398 3637 53450 3689
rect 52054 3489 52106 3541
rect 52822 3489 52874 3541
rect 54454 3489 54506 3541
rect 33046 3415 33098 3467
rect 33814 3415 33866 3467
rect 43510 3415 43562 3467
rect 44758 3415 44810 3467
rect 55222 3415 55274 3467
rect 56278 3563 56330 3615
rect 58198 3637 58250 3689
rect 59734 3637 59786 3689
rect 56374 3415 56426 3467
rect 59446 3415 59498 3467
rect 19654 3304 19706 3356
rect 19718 3304 19770 3356
rect 19782 3304 19834 3356
rect 19846 3304 19898 3356
rect 50374 3304 50426 3356
rect 50438 3304 50490 3356
rect 50502 3304 50554 3356
rect 50566 3304 50618 3356
rect 3958 3193 4010 3245
rect 5110 3193 5162 3245
rect 13270 3236 13322 3245
rect 13270 3202 13279 3236
rect 13279 3202 13313 3236
rect 13313 3202 13322 3236
rect 13270 3193 13322 3202
rect 14038 3236 14090 3245
rect 14038 3202 14047 3236
rect 14047 3202 14081 3236
rect 14081 3202 14090 3236
rect 14038 3193 14090 3202
rect 15094 3193 15146 3245
rect 16822 3236 16874 3245
rect 16822 3202 16831 3236
rect 16831 3202 16865 3236
rect 16865 3202 16874 3236
rect 16822 3193 16874 3202
rect 18070 3236 18122 3245
rect 18070 3202 18079 3236
rect 18079 3202 18113 3236
rect 18113 3202 18122 3236
rect 18070 3193 18122 3202
rect 18838 3236 18890 3245
rect 18838 3202 18847 3236
rect 18847 3202 18881 3236
rect 18881 3202 18890 3236
rect 18838 3193 18890 3202
rect 19702 3193 19754 3245
rect 20374 3193 20426 3245
rect 23350 3193 23402 3245
rect 23926 3193 23978 3245
rect 24982 3193 25034 3245
rect 26614 3193 26666 3245
rect 28822 3193 28874 3245
rect 29782 3193 29834 3245
rect 30454 3193 30506 3245
rect 31894 3193 31946 3245
rect 32662 3193 32714 3245
rect 34102 3193 34154 3245
rect 44758 3193 44810 3245
rect 46198 3193 46250 3245
rect 48502 3193 48554 3245
rect 49654 3193 49706 3245
rect 56854 3193 56906 3245
rect 58006 3193 58058 3245
rect 214 3119 266 3171
rect 1750 3119 1802 3171
rect 3094 3119 3146 3171
rect 3574 3119 3626 3171
rect 12310 3119 12362 3171
rect 12982 3119 13034 3171
rect 13846 3119 13898 3171
rect 14518 3119 14570 3171
rect 17494 3119 17546 3171
rect 18262 3119 18314 3171
rect 19894 3119 19946 3171
rect 20470 3119 20522 3171
rect 21430 3119 21482 3171
rect 23830 3119 23882 3171
rect 25078 3119 25130 3171
rect 28246 3119 28298 3171
rect 29302 3119 29354 3171
rect 29494 3119 29546 3171
rect 29878 3119 29930 3171
rect 33814 3119 33866 3171
rect 34678 3119 34730 3171
rect 35926 3119 35978 3171
rect 36886 3119 36938 3171
rect 37078 3119 37130 3171
rect 38614 3119 38666 3171
rect 44086 3119 44138 3171
rect 45430 3119 45482 3171
rect 16726 3045 16778 3097
rect 17590 3045 17642 3097
rect 18358 3045 18410 3097
rect 19030 3045 19082 3097
rect 22 2971 74 3023
rect 694 2897 746 2949
rect 2134 2897 2186 2949
rect 4918 3014 4970 3023
rect 4918 2980 4927 3014
rect 4927 2980 4961 3014
rect 4961 2980 4970 3014
rect 4918 2971 4970 2980
rect 5206 2971 5258 3023
rect 5974 2971 6026 3023
rect 5110 2749 5162 2801
rect 5782 2897 5834 2949
rect 6742 2897 6794 2949
rect 8182 2971 8234 3023
rect 12982 3014 13034 3023
rect 8950 2897 9002 2949
rect 12982 2980 12991 3014
rect 12991 2980 13025 3014
rect 13025 2980 13034 3014
rect 12982 2971 13034 2980
rect 13366 2971 13418 3023
rect 14518 2971 14570 3023
rect 16630 3014 16682 3023
rect 16630 2980 16639 3014
rect 16639 2980 16673 3014
rect 16673 2980 16682 3014
rect 16630 2971 16682 2980
rect 17014 2971 17066 3023
rect 15382 2897 15434 2949
rect 16438 2897 16490 2949
rect 17686 2897 17738 2949
rect 18838 2971 18890 3023
rect 19318 2971 19370 3023
rect 19606 2971 19658 3023
rect 22390 3045 22442 3097
rect 23542 3045 23594 3097
rect 24886 3088 24938 3097
rect 24886 3054 24895 3088
rect 24895 3054 24929 3088
rect 24929 3054 24938 3088
rect 24886 3045 24938 3054
rect 25366 3045 25418 3097
rect 26230 3045 26282 3097
rect 27478 3045 27530 3097
rect 28918 3045 28970 3097
rect 29398 3045 29450 3097
rect 31126 3045 31178 3097
rect 31894 3045 31946 3097
rect 33334 3045 33386 3097
rect 35638 3045 35690 3097
rect 36118 3045 36170 3097
rect 36694 3045 36746 3097
rect 37558 3045 37610 3097
rect 38326 3045 38378 3097
rect 8758 2866 8810 2875
rect 8758 2832 8767 2866
rect 8767 2832 8801 2866
rect 8801 2832 8810 2866
rect 8758 2823 8810 2832
rect 18262 2823 18314 2875
rect 19798 2897 19850 2949
rect 20182 2897 20234 2949
rect 21430 2971 21482 3023
rect 20470 2823 20522 2875
rect 20854 2897 20906 2949
rect 20950 2897 21002 2949
rect 21718 2897 21770 2949
rect 22486 2897 22538 2949
rect 24022 2971 24074 3023
rect 25078 2897 25130 2949
rect 26902 2971 26954 3023
rect 27670 2897 27722 2949
rect 29878 2971 29930 3023
rect 30550 2897 30602 2949
rect 32086 2971 32138 3023
rect 32278 2897 32330 2949
rect 33142 2897 33194 2949
rect 33334 2897 33386 2949
rect 35446 2971 35498 3023
rect 35350 2897 35402 2949
rect 36022 2897 36074 2949
rect 36118 2897 36170 2949
rect 39670 3045 39722 3097
rect 40918 3045 40970 3097
rect 41110 3045 41162 3097
rect 42070 3045 42122 3097
rect 42550 3045 42602 3097
rect 43318 3045 43370 3097
rect 44470 3045 44522 3097
rect 45142 3045 45194 3097
rect 40534 2971 40586 3023
rect 37558 2897 37610 2949
rect 38134 2897 38186 2949
rect 39094 2897 39146 2949
rect 41206 2897 41258 2949
rect 27958 2823 28010 2875
rect 33046 2823 33098 2875
rect 35254 2823 35306 2875
rect 43318 2897 43370 2949
rect 43510 2897 43562 2949
rect 41014 2792 41066 2801
rect 41014 2758 41023 2792
rect 41023 2758 41057 2792
rect 41057 2758 41066 2792
rect 41014 2749 41066 2758
rect 43030 2749 43082 2801
rect 43222 2749 43274 2801
rect 43990 2897 44042 2949
rect 44182 2897 44234 2949
rect 45142 2823 45194 2875
rect 46294 3119 46346 3171
rect 48118 3119 48170 3171
rect 48982 3119 49034 3171
rect 46198 3045 46250 3097
rect 47638 3045 47690 3097
rect 51766 3045 51818 3097
rect 52246 3045 52298 3097
rect 45622 2971 45674 3023
rect 46294 2897 46346 2949
rect 49654 2971 49706 3023
rect 47638 2897 47690 2949
rect 48886 2897 48938 2949
rect 48982 2897 49034 2949
rect 49846 2897 49898 2949
rect 51478 2971 51530 3023
rect 51382 2897 51434 2949
rect 51862 2897 51914 2949
rect 52246 2897 52298 2949
rect 53782 2971 53834 3023
rect 52918 2897 52970 2949
rect 53686 2897 53738 2949
rect 54838 2897 54890 2949
rect 50038 2823 50090 2875
rect 46390 2792 46442 2801
rect 46390 2758 46399 2792
rect 46399 2758 46433 2792
rect 46433 2758 46442 2792
rect 46390 2749 46442 2758
rect 52438 2749 52490 2801
rect 4294 2638 4346 2690
rect 4358 2638 4410 2690
rect 4422 2638 4474 2690
rect 4486 2638 4538 2690
rect 35014 2638 35066 2690
rect 35078 2638 35130 2690
rect 35142 2638 35194 2690
rect 35206 2638 35258 2690
rect 3958 2527 4010 2579
rect 4246 2527 4298 2579
rect 4342 2527 4394 2579
rect 4822 2527 4874 2579
rect 13750 2527 13802 2579
rect 46390 2527 46442 2579
rect 19414 2453 19466 2505
rect 19894 2453 19946 2505
rect 46102 2453 46154 2505
rect 47062 2453 47114 2505
rect 41014 2379 41066 2431
rect 49270 2379 49322 2431
rect 4726 2009 4778 2061
rect 5302 2009 5354 2061
rect 4534 1861 4586 1913
rect 4822 1861 4874 1913
rect 20182 1787 20234 1839
rect 21238 1787 21290 1839
rect 30358 1713 30410 1765
rect 30646 1713 30698 1765
rect 50518 1713 50570 1765
rect 51094 1713 51146 1765
rect 36118 1639 36170 1691
rect 35638 1565 35690 1617
rect 35158 1417 35210 1469
rect 35542 1417 35594 1469
rect 35638 1417 35690 1469
rect 35926 1417 35978 1469
rect 50710 1565 50762 1617
rect 50902 1565 50954 1617
rect 36310 1491 36362 1543
rect 33238 1269 33290 1321
rect 33718 1269 33770 1321
rect 34870 1269 34922 1321
rect 36118 1269 36170 1321
rect 41014 1417 41066 1469
rect 41302 1417 41354 1469
rect 50902 1417 50954 1469
rect 51574 1417 51626 1469
rect 36310 1121 36362 1173
rect 35446 1047 35498 1099
rect 37270 1047 37322 1099
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 226 56975 254 59200
rect 214 56969 266 56975
rect 214 56911 266 56917
rect 706 56531 734 59200
rect 694 56525 746 56531
rect 694 56467 746 56473
rect 1186 55717 1214 59200
rect 1762 57049 1790 59200
rect 1750 57043 1802 57049
rect 1750 56985 1802 56991
rect 2242 56531 2270 59200
rect 2818 56531 2846 59200
rect 3298 57049 3326 59200
rect 3286 57043 3338 57049
rect 3286 56985 3338 56991
rect 3670 56895 3722 56901
rect 3670 56837 3722 56843
rect 3574 56821 3626 56827
rect 3574 56763 3626 56769
rect 2230 56525 2282 56531
rect 2230 56467 2282 56473
rect 2806 56525 2858 56531
rect 2806 56467 2858 56473
rect 2710 56303 2762 56309
rect 2710 56245 2762 56251
rect 2806 56303 2858 56309
rect 2806 56245 2858 56251
rect 2614 56229 2666 56235
rect 2614 56171 2666 56177
rect 1174 55711 1226 55717
rect 1174 55653 1226 55659
rect 1750 55563 1802 55569
rect 1750 55505 1802 55511
rect 1762 11909 1790 55505
rect 1942 51567 1994 51573
rect 1942 51509 1994 51515
rect 1954 51203 1982 51509
rect 1942 51197 1994 51203
rect 1942 51139 1994 51145
rect 2626 47207 2654 56171
rect 2614 47201 2666 47207
rect 2614 47143 2666 47149
rect 1846 42761 1898 42767
rect 1846 42703 1898 42709
rect 1750 11903 1802 11909
rect 1750 11845 1802 11851
rect 1858 8579 1886 42703
rect 2722 33073 2750 56245
rect 2818 36551 2846 56245
rect 3286 56229 3338 56235
rect 3286 56171 3338 56177
rect 2806 36545 2858 36551
rect 2806 36487 2858 36493
rect 2710 33067 2762 33073
rect 2710 33009 2762 33015
rect 3298 28263 3326 56171
rect 3286 28257 3338 28263
rect 3286 28199 3338 28205
rect 1942 26925 1994 26931
rect 1942 26867 1994 26873
rect 1954 26561 1982 26867
rect 1942 26555 1994 26561
rect 1942 26497 1994 26503
rect 2518 19155 2570 19161
rect 2518 19097 2570 19103
rect 1846 8573 1898 8579
rect 1846 8515 1898 8521
rect 2530 8431 2558 19097
rect 2518 8425 2570 8431
rect 2518 8367 2570 8373
rect 1654 8277 1706 8283
rect 1654 8219 1706 8225
rect 2134 8277 2186 8283
rect 2134 8219 2186 8225
rect 3190 8277 3242 8283
rect 3190 8219 3242 8225
rect 1462 7685 1514 7691
rect 1462 7627 1514 7633
rect 1078 5687 1130 5693
rect 1078 5629 1130 5635
rect 310 5021 362 5027
rect 310 4963 362 4969
rect 118 3615 170 3621
rect 118 3557 170 3563
rect 22 3023 74 3029
rect 22 2965 74 2971
rect 34 800 62 2965
rect 130 800 158 3557
rect 214 3171 266 3177
rect 214 3113 266 3119
rect 226 800 254 3113
rect 322 800 350 4963
rect 790 4429 842 4435
rect 790 4371 842 4377
rect 502 3837 554 3843
rect 502 3779 554 3785
rect 514 800 542 3779
rect 598 3689 650 3695
rect 598 3631 650 3637
rect 610 800 638 3631
rect 694 2949 746 2955
rect 694 2891 746 2897
rect 706 800 734 2891
rect 802 800 830 4371
rect 982 3763 1034 3769
rect 982 3705 1034 3711
rect 994 800 1022 3705
rect 1090 800 1118 5629
rect 1174 4355 1226 4361
rect 1174 4297 1226 4303
rect 1186 800 1214 4297
rect 1366 4281 1418 4287
rect 1366 4223 1418 4229
rect 1378 800 1406 4223
rect 1474 3695 1502 7627
rect 1666 7214 1694 8219
rect 1666 7186 1790 7214
rect 1654 7019 1706 7025
rect 1654 6961 1706 6967
rect 1558 6353 1610 6359
rect 1558 6295 1610 6301
rect 1462 3689 1514 3695
rect 1462 3631 1514 3637
rect 1462 3541 1514 3547
rect 1462 3483 1514 3489
rect 1474 800 1502 3483
rect 1570 800 1598 6295
rect 1666 3843 1694 6961
rect 1654 3837 1706 3843
rect 1654 3779 1706 3785
rect 1654 3689 1706 3695
rect 1654 3631 1706 3637
rect 1666 800 1694 3631
rect 1762 3177 1790 7186
rect 2038 6353 2090 6359
rect 2038 6295 2090 6301
rect 1846 5021 1898 5027
rect 1846 4963 1898 4969
rect 1750 3171 1802 3177
rect 1750 3113 1802 3119
rect 1858 800 1886 4963
rect 1942 3911 1994 3917
rect 1942 3853 1994 3859
rect 1954 800 1982 3853
rect 2050 800 2078 6295
rect 2146 3547 2174 8219
rect 2422 7463 2474 7469
rect 2422 7405 2474 7411
rect 2998 7463 3050 7469
rect 2998 7405 3050 7411
rect 2326 3837 2378 3843
rect 2326 3779 2378 3785
rect 2134 3541 2186 3547
rect 2134 3483 2186 3489
rect 2134 2949 2186 2955
rect 2134 2891 2186 2897
rect 2146 800 2174 2891
rect 2338 800 2366 3779
rect 2434 3769 2462 7405
rect 2518 7019 2570 7025
rect 2518 6961 2570 6967
rect 2422 3763 2474 3769
rect 2422 3705 2474 3711
rect 2422 3467 2474 3473
rect 2422 3409 2474 3415
rect 2434 800 2462 3409
rect 2530 800 2558 6961
rect 2902 5687 2954 5693
rect 2902 5629 2954 5635
rect 2710 3689 2762 3695
rect 2710 3631 2762 3637
rect 2722 800 2750 3631
rect 2914 2900 2942 5629
rect 3010 3917 3038 7405
rect 3202 6452 3230 8219
rect 3202 6424 3326 6452
rect 3190 6353 3242 6359
rect 3190 6295 3242 6301
rect 3094 5021 3146 5027
rect 3094 4963 3146 4969
rect 2998 3911 3050 3917
rect 2998 3853 3050 3859
rect 3106 3843 3134 4963
rect 3094 3837 3146 3843
rect 3094 3779 3146 3785
rect 2998 3763 3050 3769
rect 2998 3705 3050 3711
rect 2818 2872 2942 2900
rect 2818 800 2846 2872
rect 3010 2752 3038 3705
rect 3094 3171 3146 3177
rect 3094 3113 3146 3119
rect 2914 2724 3038 2752
rect 2914 800 2942 2724
rect 3106 1864 3134 3113
rect 3010 1836 3134 1864
rect 3010 800 3038 1836
rect 3202 800 3230 6295
rect 3298 3769 3326 6424
rect 3586 5915 3614 56763
rect 3682 7081 3710 56837
rect 3874 56531 3902 59200
rect 4354 57614 4382 59200
rect 4354 57586 4670 57614
rect 4268 57304 4564 57324
rect 4324 57302 4348 57304
rect 4404 57302 4428 57304
rect 4484 57302 4508 57304
rect 4346 57250 4348 57302
rect 4410 57250 4422 57302
rect 4484 57250 4486 57302
rect 4324 57248 4348 57250
rect 4404 57248 4428 57250
rect 4484 57248 4508 57250
rect 4268 57228 4564 57248
rect 3862 56525 3914 56531
rect 3862 56467 3914 56473
rect 4268 55972 4564 55992
rect 4324 55970 4348 55972
rect 4404 55970 4428 55972
rect 4484 55970 4508 55972
rect 4346 55918 4348 55970
rect 4410 55918 4422 55970
rect 4484 55918 4486 55970
rect 4324 55916 4348 55918
rect 4404 55916 4428 55918
rect 4484 55916 4508 55918
rect 4268 55896 4564 55916
rect 3766 55785 3818 55791
rect 3766 55727 3818 55733
rect 3778 7839 3806 55727
rect 4642 55717 4670 57586
rect 4930 56975 4958 59200
rect 4918 56969 4970 56975
rect 4918 56911 4970 56917
rect 5110 56895 5162 56901
rect 5110 56837 5162 56843
rect 4630 55711 4682 55717
rect 4630 55653 4682 55659
rect 5014 55637 5066 55643
rect 5014 55579 5066 55585
rect 4630 55563 4682 55569
rect 4630 55505 4682 55511
rect 4268 54640 4564 54660
rect 4324 54638 4348 54640
rect 4404 54638 4428 54640
rect 4484 54638 4508 54640
rect 4346 54586 4348 54638
rect 4410 54586 4422 54638
rect 4484 54586 4486 54638
rect 4324 54584 4348 54586
rect 4404 54584 4428 54586
rect 4484 54584 4508 54586
rect 4268 54564 4564 54584
rect 4268 53308 4564 53328
rect 4324 53306 4348 53308
rect 4404 53306 4428 53308
rect 4484 53306 4508 53308
rect 4346 53254 4348 53306
rect 4410 53254 4422 53306
rect 4484 53254 4486 53306
rect 4324 53252 4348 53254
rect 4404 53252 4428 53254
rect 4484 53252 4508 53254
rect 4268 53232 4564 53252
rect 4268 51976 4564 51996
rect 4324 51974 4348 51976
rect 4404 51974 4428 51976
rect 4484 51974 4508 51976
rect 4346 51922 4348 51974
rect 4410 51922 4422 51974
rect 4484 51922 4486 51974
rect 4324 51920 4348 51922
rect 4404 51920 4428 51922
rect 4484 51920 4508 51922
rect 4268 51900 4564 51920
rect 4268 50644 4564 50664
rect 4324 50642 4348 50644
rect 4404 50642 4428 50644
rect 4484 50642 4508 50644
rect 4346 50590 4348 50642
rect 4410 50590 4422 50642
rect 4484 50590 4486 50642
rect 4324 50588 4348 50590
rect 4404 50588 4428 50590
rect 4484 50588 4508 50590
rect 4268 50568 4564 50588
rect 4268 49312 4564 49332
rect 4324 49310 4348 49312
rect 4404 49310 4428 49312
rect 4484 49310 4508 49312
rect 4346 49258 4348 49310
rect 4410 49258 4422 49310
rect 4484 49258 4486 49310
rect 4324 49256 4348 49258
rect 4404 49256 4428 49258
rect 4484 49256 4508 49258
rect 4268 49236 4564 49256
rect 4268 47980 4564 48000
rect 4324 47978 4348 47980
rect 4404 47978 4428 47980
rect 4484 47978 4508 47980
rect 4346 47926 4348 47978
rect 4410 47926 4422 47978
rect 4484 47926 4486 47978
rect 4324 47924 4348 47926
rect 4404 47924 4428 47926
rect 4484 47924 4508 47926
rect 4268 47904 4564 47924
rect 4268 46648 4564 46668
rect 4324 46646 4348 46648
rect 4404 46646 4428 46648
rect 4484 46646 4508 46648
rect 4346 46594 4348 46646
rect 4410 46594 4422 46646
rect 4484 46594 4486 46646
rect 4324 46592 4348 46594
rect 4404 46592 4428 46594
rect 4484 46592 4508 46594
rect 4268 46572 4564 46592
rect 4268 45316 4564 45336
rect 4324 45314 4348 45316
rect 4404 45314 4428 45316
rect 4484 45314 4508 45316
rect 4346 45262 4348 45314
rect 4410 45262 4422 45314
rect 4484 45262 4486 45314
rect 4324 45260 4348 45262
rect 4404 45260 4428 45262
rect 4484 45260 4508 45262
rect 4268 45240 4564 45260
rect 4268 43984 4564 44004
rect 4324 43982 4348 43984
rect 4404 43982 4428 43984
rect 4484 43982 4508 43984
rect 4346 43930 4348 43982
rect 4410 43930 4422 43982
rect 4484 43930 4486 43982
rect 4324 43928 4348 43930
rect 4404 43928 4428 43930
rect 4484 43928 4508 43930
rect 4268 43908 4564 43928
rect 4268 42652 4564 42672
rect 4324 42650 4348 42652
rect 4404 42650 4428 42652
rect 4484 42650 4508 42652
rect 4346 42598 4348 42650
rect 4410 42598 4422 42650
rect 4484 42598 4486 42650
rect 4324 42596 4348 42598
rect 4404 42596 4428 42598
rect 4484 42596 4508 42598
rect 4268 42576 4564 42596
rect 4268 41320 4564 41340
rect 4324 41318 4348 41320
rect 4404 41318 4428 41320
rect 4484 41318 4508 41320
rect 4346 41266 4348 41318
rect 4410 41266 4422 41318
rect 4484 41266 4486 41318
rect 4324 41264 4348 41266
rect 4404 41264 4428 41266
rect 4484 41264 4508 41266
rect 4268 41244 4564 41264
rect 4268 39988 4564 40008
rect 4324 39986 4348 39988
rect 4404 39986 4428 39988
rect 4484 39986 4508 39988
rect 4346 39934 4348 39986
rect 4410 39934 4422 39986
rect 4484 39934 4486 39986
rect 4324 39932 4348 39934
rect 4404 39932 4428 39934
rect 4484 39932 4508 39934
rect 4268 39912 4564 39932
rect 4268 38656 4564 38676
rect 4324 38654 4348 38656
rect 4404 38654 4428 38656
rect 4484 38654 4508 38656
rect 4346 38602 4348 38654
rect 4410 38602 4422 38654
rect 4484 38602 4486 38654
rect 4324 38600 4348 38602
rect 4404 38600 4428 38602
rect 4484 38600 4508 38602
rect 4268 38580 4564 38600
rect 4054 38099 4106 38105
rect 4054 38041 4106 38047
rect 3766 7833 3818 7839
rect 3766 7775 3818 7781
rect 4066 7691 4094 38041
rect 4268 37324 4564 37344
rect 4324 37322 4348 37324
rect 4404 37322 4428 37324
rect 4484 37322 4508 37324
rect 4346 37270 4348 37322
rect 4410 37270 4422 37322
rect 4484 37270 4486 37322
rect 4324 37268 4348 37270
rect 4404 37268 4428 37270
rect 4484 37268 4508 37270
rect 4268 37248 4564 37268
rect 4268 35992 4564 36012
rect 4324 35990 4348 35992
rect 4404 35990 4428 35992
rect 4484 35990 4508 35992
rect 4346 35938 4348 35990
rect 4410 35938 4422 35990
rect 4484 35938 4486 35990
rect 4324 35936 4348 35938
rect 4404 35936 4428 35938
rect 4484 35936 4508 35938
rect 4268 35916 4564 35936
rect 4268 34660 4564 34680
rect 4324 34658 4348 34660
rect 4404 34658 4428 34660
rect 4484 34658 4508 34660
rect 4346 34606 4348 34658
rect 4410 34606 4422 34658
rect 4484 34606 4486 34658
rect 4324 34604 4348 34606
rect 4404 34604 4428 34606
rect 4484 34604 4508 34606
rect 4268 34584 4564 34604
rect 4268 33328 4564 33348
rect 4324 33326 4348 33328
rect 4404 33326 4428 33328
rect 4484 33326 4508 33328
rect 4346 33274 4348 33326
rect 4410 33274 4422 33326
rect 4484 33274 4486 33326
rect 4324 33272 4348 33274
rect 4404 33272 4428 33274
rect 4484 33272 4508 33274
rect 4268 33252 4564 33272
rect 4642 33134 4670 55505
rect 5026 37217 5054 55579
rect 5014 37211 5066 37217
rect 5014 37153 5066 37159
rect 4642 33106 4862 33134
rect 4268 31996 4564 32016
rect 4324 31994 4348 31996
rect 4404 31994 4428 31996
rect 4484 31994 4508 31996
rect 4346 31942 4348 31994
rect 4410 31942 4422 31994
rect 4484 31942 4486 31994
rect 4324 31940 4348 31942
rect 4404 31940 4428 31942
rect 4484 31940 4508 31942
rect 4268 31920 4564 31940
rect 4268 30664 4564 30684
rect 4324 30662 4348 30664
rect 4404 30662 4428 30664
rect 4484 30662 4508 30664
rect 4346 30610 4348 30662
rect 4410 30610 4422 30662
rect 4484 30610 4486 30662
rect 4324 30608 4348 30610
rect 4404 30608 4428 30610
rect 4484 30608 4508 30610
rect 4268 30588 4564 30608
rect 4268 29332 4564 29352
rect 4324 29330 4348 29332
rect 4404 29330 4428 29332
rect 4484 29330 4508 29332
rect 4346 29278 4348 29330
rect 4410 29278 4422 29330
rect 4484 29278 4486 29330
rect 4324 29276 4348 29278
rect 4404 29276 4428 29278
rect 4484 29276 4508 29278
rect 4268 29256 4564 29276
rect 4268 28000 4564 28020
rect 4324 27998 4348 28000
rect 4404 27998 4428 28000
rect 4484 27998 4508 28000
rect 4346 27946 4348 27998
rect 4410 27946 4422 27998
rect 4484 27946 4486 27998
rect 4324 27944 4348 27946
rect 4404 27944 4428 27946
rect 4484 27944 4508 27946
rect 4268 27924 4564 27944
rect 4268 26668 4564 26688
rect 4324 26666 4348 26668
rect 4404 26666 4428 26668
rect 4484 26666 4508 26668
rect 4346 26614 4348 26666
rect 4410 26614 4422 26666
rect 4484 26614 4486 26666
rect 4324 26612 4348 26614
rect 4404 26612 4428 26614
rect 4484 26612 4508 26614
rect 4268 26592 4564 26612
rect 4268 25336 4564 25356
rect 4324 25334 4348 25336
rect 4404 25334 4428 25336
rect 4484 25334 4508 25336
rect 4346 25282 4348 25334
rect 4410 25282 4422 25334
rect 4484 25282 4486 25334
rect 4324 25280 4348 25282
rect 4404 25280 4428 25282
rect 4484 25280 4508 25282
rect 4268 25260 4564 25280
rect 4268 24004 4564 24024
rect 4324 24002 4348 24004
rect 4404 24002 4428 24004
rect 4484 24002 4508 24004
rect 4346 23950 4348 24002
rect 4410 23950 4422 24002
rect 4484 23950 4486 24002
rect 4324 23948 4348 23950
rect 4404 23948 4428 23950
rect 4484 23948 4508 23950
rect 4268 23928 4564 23948
rect 4268 22672 4564 22692
rect 4324 22670 4348 22672
rect 4404 22670 4428 22672
rect 4484 22670 4508 22672
rect 4346 22618 4348 22670
rect 4410 22618 4422 22670
rect 4484 22618 4486 22670
rect 4324 22616 4348 22618
rect 4404 22616 4428 22618
rect 4484 22616 4508 22618
rect 4268 22596 4564 22616
rect 4268 21340 4564 21360
rect 4324 21338 4348 21340
rect 4404 21338 4428 21340
rect 4484 21338 4508 21340
rect 4346 21286 4348 21338
rect 4410 21286 4422 21338
rect 4484 21286 4486 21338
rect 4324 21284 4348 21286
rect 4404 21284 4428 21286
rect 4484 21284 4508 21286
rect 4268 21264 4564 21284
rect 4268 20008 4564 20028
rect 4324 20006 4348 20008
rect 4404 20006 4428 20008
rect 4484 20006 4508 20008
rect 4346 19954 4348 20006
rect 4410 19954 4422 20006
rect 4484 19954 4486 20006
rect 4324 19952 4348 19954
rect 4404 19952 4428 19954
rect 4484 19952 4508 19954
rect 4268 19932 4564 19952
rect 4268 18676 4564 18696
rect 4324 18674 4348 18676
rect 4404 18674 4428 18676
rect 4484 18674 4508 18676
rect 4346 18622 4348 18674
rect 4410 18622 4422 18674
rect 4484 18622 4486 18674
rect 4324 18620 4348 18622
rect 4404 18620 4428 18622
rect 4484 18620 4508 18622
rect 4268 18600 4564 18620
rect 4268 17344 4564 17364
rect 4324 17342 4348 17344
rect 4404 17342 4428 17344
rect 4484 17342 4508 17344
rect 4346 17290 4348 17342
rect 4410 17290 4422 17342
rect 4484 17290 4486 17342
rect 4324 17288 4348 17290
rect 4404 17288 4428 17290
rect 4484 17288 4508 17290
rect 4268 17268 4564 17288
rect 4268 16012 4564 16032
rect 4324 16010 4348 16012
rect 4404 16010 4428 16012
rect 4484 16010 4508 16012
rect 4346 15958 4348 16010
rect 4410 15958 4422 16010
rect 4484 15958 4486 16010
rect 4324 15956 4348 15958
rect 4404 15956 4428 15958
rect 4484 15956 4508 15958
rect 4268 15936 4564 15956
rect 4268 14680 4564 14700
rect 4324 14678 4348 14680
rect 4404 14678 4428 14680
rect 4484 14678 4508 14680
rect 4346 14626 4348 14678
rect 4410 14626 4422 14678
rect 4484 14626 4486 14678
rect 4324 14624 4348 14626
rect 4404 14624 4428 14626
rect 4484 14624 4508 14626
rect 4268 14604 4564 14624
rect 4726 14123 4778 14129
rect 4726 14065 4778 14071
rect 4738 13907 4766 14065
rect 4726 13901 4778 13907
rect 4726 13843 4778 13849
rect 4268 13348 4564 13368
rect 4324 13346 4348 13348
rect 4404 13346 4428 13348
rect 4484 13346 4508 13348
rect 4346 13294 4348 13346
rect 4410 13294 4422 13346
rect 4484 13294 4486 13346
rect 4324 13292 4348 13294
rect 4404 13292 4428 13294
rect 4484 13292 4508 13294
rect 4268 13272 4564 13292
rect 4834 12974 4862 33106
rect 4834 12946 5054 12974
rect 4268 12016 4564 12036
rect 4324 12014 4348 12016
rect 4404 12014 4428 12016
rect 4484 12014 4508 12016
rect 4346 11962 4348 12014
rect 4410 11962 4422 12014
rect 4484 11962 4486 12014
rect 4324 11960 4348 11962
rect 4404 11960 4428 11962
rect 4484 11960 4508 11962
rect 4268 11940 4564 11960
rect 4268 10684 4564 10704
rect 4324 10682 4348 10684
rect 4404 10682 4428 10684
rect 4484 10682 4508 10684
rect 4346 10630 4348 10682
rect 4410 10630 4422 10682
rect 4484 10630 4486 10682
rect 4324 10628 4348 10630
rect 4404 10628 4428 10630
rect 4484 10628 4508 10630
rect 4268 10608 4564 10628
rect 4268 9352 4564 9372
rect 4324 9350 4348 9352
rect 4404 9350 4428 9352
rect 4484 9350 4508 9352
rect 4346 9298 4348 9350
rect 4410 9298 4422 9350
rect 4484 9298 4486 9350
rect 4324 9296 4348 9298
rect 4404 9296 4428 9298
rect 4484 9296 4508 9298
rect 4268 9276 4564 9296
rect 4918 8499 4970 8505
rect 4918 8441 4970 8447
rect 4822 8203 4874 8209
rect 4822 8145 4874 8151
rect 4268 8020 4564 8040
rect 4324 8018 4348 8020
rect 4404 8018 4428 8020
rect 4484 8018 4508 8020
rect 4346 7966 4348 8018
rect 4410 7966 4422 8018
rect 4484 7966 4486 8018
rect 4324 7964 4348 7966
rect 4404 7964 4428 7966
rect 4484 7964 4508 7966
rect 4268 7944 4564 7964
rect 4054 7685 4106 7691
rect 4054 7627 4106 7633
rect 3958 7463 4010 7469
rect 3958 7405 4010 7411
rect 4054 7463 4106 7469
rect 4054 7405 4106 7411
rect 3682 7053 3806 7081
rect 3670 7019 3722 7025
rect 3670 6961 3722 6967
rect 3574 5909 3626 5915
rect 3574 5851 3626 5857
rect 3478 4207 3530 4213
rect 3478 4149 3530 4155
rect 3286 3763 3338 3769
rect 3286 3705 3338 3711
rect 3382 3763 3434 3769
rect 3382 3705 3434 3711
rect 3286 3467 3338 3473
rect 3286 3409 3338 3415
rect 3298 800 3326 3409
rect 3394 800 3422 3705
rect 3490 800 3518 4149
rect 3574 3689 3626 3695
rect 3574 3631 3626 3637
rect 3586 3177 3614 3631
rect 3574 3171 3626 3177
rect 3574 3113 3626 3119
rect 3682 800 3710 6961
rect 3778 5471 3806 7053
rect 3862 6353 3914 6359
rect 3862 6295 3914 6301
rect 3766 5465 3818 5471
rect 3766 5407 3818 5413
rect 3766 4281 3818 4287
rect 3766 4223 3818 4229
rect 3778 800 3806 4223
rect 3874 800 3902 6295
rect 3970 3473 3998 7405
rect 3958 3467 4010 3473
rect 3958 3409 4010 3415
rect 3958 3245 4010 3251
rect 3958 3187 4010 3193
rect 3970 2585 3998 3187
rect 3958 2579 4010 2585
rect 3958 2521 4010 2527
rect 4066 800 4094 7405
rect 4268 6688 4564 6708
rect 4324 6686 4348 6688
rect 4404 6686 4428 6688
rect 4484 6686 4508 6688
rect 4346 6634 4348 6686
rect 4410 6634 4422 6686
rect 4484 6634 4486 6686
rect 4324 6632 4348 6634
rect 4404 6632 4428 6634
rect 4484 6632 4508 6634
rect 4268 6612 4564 6632
rect 4630 6353 4682 6359
rect 4630 6295 4682 6301
rect 4268 5356 4564 5376
rect 4324 5354 4348 5356
rect 4404 5354 4428 5356
rect 4484 5354 4508 5356
rect 4346 5302 4348 5354
rect 4410 5302 4422 5354
rect 4484 5302 4486 5354
rect 4324 5300 4348 5302
rect 4404 5300 4428 5302
rect 4484 5300 4508 5302
rect 4268 5280 4564 5300
rect 4150 5021 4202 5027
rect 4150 4963 4202 4969
rect 4162 800 4190 4963
rect 4268 4024 4564 4044
rect 4324 4022 4348 4024
rect 4404 4022 4428 4024
rect 4484 4022 4508 4024
rect 4346 3970 4348 4022
rect 4410 3970 4422 4022
rect 4484 3970 4486 4022
rect 4324 3968 4348 3970
rect 4404 3968 4428 3970
rect 4484 3968 4508 3970
rect 4268 3948 4564 3968
rect 4268 2692 4564 2712
rect 4324 2690 4348 2692
rect 4404 2690 4428 2692
rect 4484 2690 4508 2692
rect 4346 2638 4348 2690
rect 4410 2638 4422 2690
rect 4484 2638 4486 2690
rect 4324 2636 4348 2638
rect 4404 2636 4428 2638
rect 4484 2636 4508 2638
rect 4268 2616 4564 2636
rect 4246 2579 4298 2585
rect 4246 2521 4298 2527
rect 4342 2579 4394 2585
rect 4342 2521 4394 2527
rect 4258 800 4286 2521
rect 4354 800 4382 2521
rect 4642 2456 4670 6295
rect 4726 4355 4778 4361
rect 4726 4297 4778 4303
rect 4450 2428 4670 2456
rect 4450 2012 4478 2428
rect 4738 2160 4766 4297
rect 4834 2585 4862 8145
rect 4930 7691 4958 8441
rect 4918 7685 4970 7691
rect 4918 7627 4970 7633
rect 4918 5687 4970 5693
rect 4918 5629 4970 5635
rect 4930 4213 4958 5629
rect 5026 5249 5054 12946
rect 5122 8431 5150 56837
rect 5410 56531 5438 59200
rect 5986 56531 6014 59200
rect 6466 56975 6494 59200
rect 6454 56969 6506 56975
rect 6454 56911 6506 56917
rect 7042 56531 7070 59200
rect 5398 56525 5450 56531
rect 5398 56467 5450 56473
rect 5974 56525 6026 56531
rect 5974 56467 6026 56473
rect 7030 56525 7082 56531
rect 7030 56467 7082 56473
rect 5590 56229 5642 56235
rect 5590 56171 5642 56177
rect 5974 56229 6026 56235
rect 5974 56171 6026 56177
rect 7222 56229 7274 56235
rect 7222 56171 7274 56177
rect 5602 42101 5630 56171
rect 5590 42095 5642 42101
rect 5590 42037 5642 42043
rect 5302 35435 5354 35441
rect 5302 35377 5354 35383
rect 5206 12199 5258 12205
rect 5206 12141 5258 12147
rect 5218 11909 5246 12141
rect 5206 11903 5258 11909
rect 5206 11845 5258 11851
rect 5110 8425 5162 8431
rect 5314 8413 5342 35377
rect 5986 28337 6014 56171
rect 6454 53417 6506 53423
rect 6454 53359 6506 53365
rect 6070 46535 6122 46541
rect 6070 46477 6122 46483
rect 5974 28331 6026 28337
rect 5974 28273 6026 28279
rect 5398 27591 5450 27597
rect 5398 27533 5450 27539
rect 5410 8579 5438 27533
rect 5974 16935 6026 16941
rect 5974 16877 6026 16883
rect 5986 16571 6014 16877
rect 5974 16565 6026 16571
rect 5974 16507 6026 16513
rect 5398 8573 5450 8579
rect 5398 8515 5450 8521
rect 5314 8385 5438 8413
rect 5110 8367 5162 8373
rect 5302 7463 5354 7469
rect 5302 7405 5354 7411
rect 5206 6797 5258 6803
rect 5206 6739 5258 6745
rect 5110 5687 5162 5693
rect 5110 5629 5162 5635
rect 5014 5243 5066 5249
rect 5014 5185 5066 5191
rect 5014 4281 5066 4287
rect 5014 4223 5066 4229
rect 4918 4207 4970 4213
rect 4918 4149 4970 4155
rect 4918 3023 4970 3029
rect 4918 2965 4970 2971
rect 4822 2579 4874 2585
rect 4822 2521 4874 2527
rect 4738 2132 4862 2160
rect 4726 2061 4778 2067
rect 4450 1984 4670 2012
rect 4726 2003 4778 2009
rect 4534 1913 4586 1919
rect 4534 1855 4586 1861
rect 4546 800 4574 1855
rect 4642 800 4670 1984
rect 4738 800 4766 2003
rect 4834 1919 4862 2132
rect 4822 1913 4874 1919
rect 4822 1855 4874 1861
rect 4930 800 4958 2965
rect 5026 800 5054 4223
rect 5122 3251 5150 5629
rect 5218 3621 5246 6739
rect 5206 3615 5258 3621
rect 5206 3557 5258 3563
rect 5110 3245 5162 3251
rect 5110 3187 5162 3193
rect 5206 3023 5258 3029
rect 5206 2965 5258 2971
rect 5110 2801 5162 2807
rect 5110 2743 5162 2749
rect 5122 800 5150 2743
rect 5218 800 5246 2965
rect 5314 2067 5342 7405
rect 5410 6581 5438 8385
rect 5494 8129 5546 8135
rect 5494 8071 5546 8077
rect 5506 7765 5534 8071
rect 5494 7759 5546 7765
rect 5494 7701 5546 7707
rect 5590 7611 5642 7617
rect 5590 7553 5642 7559
rect 5602 7247 5630 7553
rect 5590 7241 5642 7247
rect 5590 7183 5642 7189
rect 6082 7099 6110 46477
rect 6466 15854 6494 53359
rect 7234 46097 7262 56171
rect 7522 55717 7550 59200
rect 8098 56975 8126 59200
rect 8086 56969 8138 56975
rect 8086 56911 8138 56917
rect 8278 56895 8330 56901
rect 8278 56837 8330 56843
rect 8182 56229 8234 56235
rect 8182 56171 8234 56177
rect 7510 55711 7562 55717
rect 7510 55653 7562 55659
rect 7702 55563 7754 55569
rect 7702 55505 7754 55511
rect 7222 46091 7274 46097
rect 7222 46033 7274 46039
rect 6550 45425 6602 45431
rect 6550 45367 6602 45373
rect 6562 45209 6590 45367
rect 6550 45203 6602 45209
rect 6550 45145 6602 45151
rect 7714 37454 7742 55505
rect 8194 37454 8222 56171
rect 7714 37426 7838 37454
rect 7810 33134 7838 37426
rect 7714 33106 7838 33134
rect 8098 37426 8222 37454
rect 8290 37454 8318 56837
rect 8578 56531 8606 59200
rect 8566 56525 8618 56531
rect 8566 56467 8618 56473
rect 9154 55717 9182 59200
rect 9634 57049 9662 59200
rect 9622 57043 9674 57049
rect 9622 56985 9674 56991
rect 9814 56747 9866 56753
rect 9814 56689 9866 56695
rect 9142 55711 9194 55717
rect 9142 55653 9194 55659
rect 8950 55415 9002 55421
rect 8950 55357 9002 55363
rect 8290 37426 8414 37454
rect 6550 28109 6602 28115
rect 6550 28051 6602 28057
rect 6370 15826 6494 15854
rect 6070 7093 6122 7099
rect 6070 7035 6122 7041
rect 6370 7025 6398 15826
rect 6562 7173 6590 28051
rect 7714 23054 7742 33106
rect 8098 25100 8126 37426
rect 8278 29515 8330 29521
rect 8278 29457 8330 29463
rect 8290 29244 8318 29457
rect 8242 29216 8318 29244
rect 8242 28929 8270 29216
rect 8230 28923 8282 28929
rect 8230 28865 8282 28871
rect 8182 28183 8234 28189
rect 8182 28125 8234 28131
rect 8194 27523 8222 28125
rect 8182 27517 8234 27523
rect 8182 27459 8234 27465
rect 8098 25072 8222 25100
rect 8086 25001 8138 25007
rect 8086 24943 8138 24949
rect 8098 24563 8126 24943
rect 8086 24557 8138 24563
rect 8086 24499 8138 24505
rect 8086 23521 8138 23527
rect 8086 23463 8138 23469
rect 8098 23231 8126 23463
rect 8086 23225 8138 23231
rect 8086 23167 8138 23173
rect 8194 23054 8222 25072
rect 7714 23026 7838 23054
rect 7606 20783 7658 20789
rect 7606 20725 7658 20731
rect 7618 20567 7646 20725
rect 7606 20561 7658 20567
rect 7606 20503 7658 20509
rect 7606 20117 7658 20123
rect 7606 20059 7658 20065
rect 7618 19901 7646 20059
rect 7606 19895 7658 19901
rect 7606 19837 7658 19843
rect 7126 19599 7178 19605
rect 7126 19541 7178 19547
rect 7138 19235 7166 19541
rect 7126 19229 7178 19235
rect 7126 19171 7178 19177
rect 7414 18267 7466 18273
rect 7414 18209 7466 18215
rect 7426 17533 7454 18209
rect 7810 17903 7838 23026
rect 7906 23026 8222 23054
rect 7798 17897 7850 17903
rect 7798 17839 7850 17845
rect 7414 17527 7466 17533
rect 7414 17469 7466 17475
rect 7126 16935 7178 16941
rect 7126 16877 7178 16883
rect 7138 16497 7166 16877
rect 7126 16491 7178 16497
rect 7126 16433 7178 16439
rect 7702 14863 7754 14869
rect 7702 14805 7754 14811
rect 7606 13679 7658 13685
rect 7606 13621 7658 13627
rect 7618 13241 7646 13621
rect 7606 13235 7658 13241
rect 7606 13177 7658 13183
rect 6838 12421 6890 12427
rect 6838 12363 6890 12369
rect 6850 8283 6878 12363
rect 7606 8795 7658 8801
rect 7606 8737 7658 8743
rect 7618 8579 7646 8737
rect 7606 8573 7658 8579
rect 7606 8515 7658 8521
rect 7222 8425 7274 8431
rect 7714 8413 7742 14805
rect 7798 9461 7850 9467
rect 7798 9403 7850 9409
rect 7222 8367 7274 8373
rect 7618 8385 7742 8413
rect 6838 8277 6890 8283
rect 6838 8219 6890 8225
rect 6550 7167 6602 7173
rect 6550 7109 6602 7115
rect 7126 7093 7178 7099
rect 7126 7035 7178 7041
rect 6358 7019 6410 7025
rect 6358 6961 6410 6967
rect 7030 7019 7082 7025
rect 7030 6961 7082 6967
rect 5878 6945 5930 6951
rect 5878 6887 5930 6893
rect 6550 6945 6602 6951
rect 6550 6887 6602 6893
rect 6934 6945 6986 6951
rect 6934 6887 6986 6893
rect 5398 6575 5450 6581
rect 5398 6517 5450 6523
rect 5494 6131 5546 6137
rect 5494 6073 5546 6079
rect 5398 5021 5450 5027
rect 5398 4963 5450 4969
rect 5302 2061 5354 2067
rect 5302 2003 5354 2009
rect 5410 800 5438 4963
rect 5506 800 5534 6073
rect 5782 5687 5834 5693
rect 5782 5629 5834 5635
rect 5686 4281 5738 4287
rect 5686 4223 5738 4229
rect 5590 3689 5642 3695
rect 5590 3631 5642 3637
rect 5602 800 5630 3631
rect 5698 800 5726 4223
rect 5794 2955 5822 5629
rect 5782 2949 5834 2955
rect 5782 2891 5834 2897
rect 5890 800 5918 6887
rect 6262 6131 6314 6137
rect 6262 6073 6314 6079
rect 6070 5021 6122 5027
rect 6070 4963 6122 4969
rect 5974 3023 6026 3029
rect 5974 2965 6026 2971
rect 5986 800 6014 2965
rect 6082 800 6110 4963
rect 6274 800 6302 6073
rect 6454 4207 6506 4213
rect 6454 4149 6506 4155
rect 6358 3689 6410 3695
rect 6358 3631 6410 3637
rect 6370 800 6398 3631
rect 6466 800 6494 4149
rect 6562 800 6590 6887
rect 6838 5687 6890 5693
rect 6838 5629 6890 5635
rect 6742 2949 6794 2955
rect 6742 2891 6794 2897
rect 6754 800 6782 2891
rect 6850 800 6878 5629
rect 6946 800 6974 6887
rect 7042 5767 7070 6961
rect 7138 6433 7166 7035
rect 7234 6433 7262 8367
rect 7618 7025 7646 8385
rect 7702 8277 7754 8283
rect 7702 8219 7754 8225
rect 7606 7019 7658 7025
rect 7606 6961 7658 6967
rect 7318 6871 7370 6877
rect 7318 6813 7370 6819
rect 7126 6427 7178 6433
rect 7126 6369 7178 6375
rect 7222 6427 7274 6433
rect 7222 6369 7274 6375
rect 7030 5761 7082 5767
rect 7030 5703 7082 5709
rect 7222 5687 7274 5693
rect 7222 5629 7274 5635
rect 7030 3689 7082 3695
rect 7030 3631 7082 3637
rect 7042 800 7070 3631
rect 7234 800 7262 5629
rect 7330 800 7358 6813
rect 7606 5539 7658 5545
rect 7606 5481 7658 5487
rect 7414 4355 7466 4361
rect 7414 4297 7466 4303
rect 7426 800 7454 4297
rect 7618 800 7646 5481
rect 7714 800 7742 8219
rect 7810 7839 7838 9403
rect 7906 9245 7934 23026
rect 8086 22855 8138 22861
rect 8086 22797 8138 22803
rect 8098 22343 8126 22797
rect 8086 22337 8138 22343
rect 8086 22279 8138 22285
rect 8086 21597 8138 21603
rect 8086 21539 8138 21545
rect 8098 20957 8126 21539
rect 8086 20951 8138 20957
rect 8086 20893 8138 20899
rect 8278 19525 8330 19531
rect 8276 19490 8278 19499
rect 8330 19490 8332 19499
rect 8276 19425 8332 19434
rect 8086 18267 8138 18273
rect 8086 18209 8138 18215
rect 8098 17755 8126 18209
rect 8086 17749 8138 17755
rect 8086 17691 8138 17697
rect 8386 15854 8414 37426
rect 8662 29589 8714 29595
rect 8662 29531 8714 29537
rect 8674 28929 8702 29531
rect 8662 28923 8714 28929
rect 8662 28865 8714 28871
rect 8615 28775 8667 28781
rect 8615 28717 8667 28723
rect 8627 28559 8655 28717
rect 8615 28553 8667 28559
rect 8615 28495 8667 28501
rect 8758 24779 8810 24785
rect 8758 24721 8810 24727
rect 8470 23447 8522 23453
rect 8470 23389 8522 23395
rect 8482 23157 8510 23389
rect 8470 23151 8522 23157
rect 8470 23093 8522 23099
rect 8770 23054 8798 24721
rect 8674 23026 8798 23054
rect 8566 21449 8618 21455
rect 8566 21391 8618 21397
rect 8578 20789 8606 21391
rect 8566 20783 8618 20789
rect 8566 20725 8618 20731
rect 8566 17527 8618 17533
rect 8566 17469 8618 17475
rect 8194 15826 8414 15854
rect 8086 12347 8138 12353
rect 8086 12289 8138 12295
rect 8098 11761 8126 12289
rect 8086 11755 8138 11761
rect 8086 11697 8138 11703
rect 8086 11015 8138 11021
rect 8086 10957 8138 10963
rect 8098 10207 8126 10957
rect 8086 10201 8138 10207
rect 8086 10143 8138 10149
rect 8194 10004 8222 15826
rect 8374 13531 8426 13537
rect 8374 13473 8426 13479
rect 8386 13167 8414 13473
rect 8578 13463 8606 17469
rect 8566 13457 8618 13463
rect 8566 13399 8618 13405
rect 8374 13161 8426 13167
rect 8374 13103 8426 13109
rect 8566 12569 8618 12575
rect 8566 12511 8618 12517
rect 8578 11928 8606 12511
rect 8386 11909 8606 11928
rect 8374 11903 8606 11909
rect 8426 11900 8606 11903
rect 8374 11845 8426 11851
rect 8578 11835 8606 11900
rect 8566 11829 8618 11835
rect 8566 11771 8618 11777
rect 8674 11243 8702 23026
rect 8758 20783 8810 20789
rect 8758 20725 8810 20731
rect 8770 20567 8798 20725
rect 8758 20561 8810 20567
rect 8758 20503 8810 20509
rect 8758 20117 8810 20123
rect 8758 20059 8810 20065
rect 8770 19901 8798 20059
rect 8758 19895 8810 19901
rect 8758 19837 8810 19843
rect 8962 15854 8990 55357
rect 9334 27887 9386 27893
rect 9334 27829 9386 27835
rect 9346 27616 9374 27829
rect 9250 27588 9374 27616
rect 9250 27468 9278 27588
rect 9058 27449 9278 27468
rect 9334 27517 9386 27523
rect 9386 27465 9662 27468
rect 9334 27459 9662 27465
rect 9046 27443 9278 27449
rect 9098 27440 9278 27443
rect 9346 27449 9662 27459
rect 9346 27443 9674 27449
rect 9346 27440 9622 27443
rect 9046 27385 9098 27391
rect 9622 27385 9674 27391
rect 9334 20783 9386 20789
rect 9334 20725 9386 20731
rect 9346 20567 9374 20725
rect 9334 20561 9386 20567
rect 9334 20503 9386 20509
rect 9046 19525 9098 19531
rect 9044 19490 9046 19499
rect 9098 19490 9100 19499
rect 9044 19425 9100 19434
rect 9826 15854 9854 56689
rect 10210 56531 10238 59200
rect 10690 56531 10718 59200
rect 11266 57049 11294 59200
rect 11254 57043 11306 57049
rect 11254 56985 11306 56991
rect 11254 56895 11306 56901
rect 11254 56837 11306 56843
rect 10774 56821 10826 56827
rect 10774 56763 10826 56769
rect 10198 56525 10250 56531
rect 10198 56467 10250 56473
rect 10678 56525 10730 56531
rect 10678 56467 10730 56473
rect 10102 56229 10154 56235
rect 10102 56171 10154 56177
rect 10114 28855 10142 56171
rect 10678 46757 10730 46763
rect 10678 46699 10730 46705
rect 10690 46541 10718 46699
rect 10678 46535 10730 46541
rect 10678 46477 10730 46483
rect 10102 28849 10154 28855
rect 10102 28791 10154 28797
rect 10582 22929 10634 22935
rect 10582 22871 10634 22877
rect 10594 22195 10622 22871
rect 10582 22189 10634 22195
rect 10582 22131 10634 22137
rect 8962 15826 9182 15854
rect 8662 11237 8714 11243
rect 8662 11179 8714 11185
rect 8194 9976 8414 10004
rect 8086 9905 8138 9911
rect 8086 9847 8138 9853
rect 7990 9831 8042 9837
rect 7990 9773 8042 9779
rect 7894 9239 7946 9245
rect 7894 9181 7946 9187
rect 8002 8431 8030 9773
rect 8098 9023 8126 9847
rect 8278 9683 8330 9689
rect 8278 9625 8330 9631
rect 8290 9116 8318 9625
rect 8242 9088 8318 9116
rect 8242 9023 8270 9088
rect 8086 9017 8138 9023
rect 8086 8959 8138 8965
rect 8230 9017 8282 9023
rect 8230 8959 8282 8965
rect 7990 8425 8042 8431
rect 7990 8367 8042 8373
rect 8086 8425 8138 8431
rect 8086 8367 8138 8373
rect 7798 7833 7850 7839
rect 7798 7775 7850 7781
rect 7940 7798 7996 7807
rect 7940 7733 7942 7742
rect 7994 7733 7996 7742
rect 7942 7701 7994 7707
rect 8098 7617 8126 8367
rect 8086 7611 8138 7617
rect 8086 7553 8138 7559
rect 8086 6797 8138 6803
rect 8086 6739 8138 6745
rect 7798 5909 7850 5915
rect 7798 5851 7850 5857
rect 7810 4972 7838 5851
rect 7810 4953 7982 4972
rect 7810 4947 7994 4953
rect 7810 4944 7942 4947
rect 7942 4889 7994 4895
rect 7894 4577 7946 4583
rect 7894 4519 7946 4525
rect 7798 3689 7850 3695
rect 7798 3631 7850 3637
rect 7810 800 7838 3631
rect 7906 800 7934 4519
rect 8098 800 8126 6739
rect 8386 6433 8414 9976
rect 8530 9097 8990 9116
rect 8518 9091 8990 9097
rect 8570 9088 8990 9091
rect 8518 9033 8570 9039
rect 8962 9023 8990 9088
rect 8950 9017 9002 9023
rect 8950 8959 9002 8965
rect 8866 8801 9086 8820
rect 8854 8795 9098 8801
rect 8906 8792 9046 8795
rect 8854 8737 8906 8743
rect 9046 8737 9098 8743
rect 8866 8579 8894 8737
rect 8854 8573 8906 8579
rect 8854 8515 8906 8521
rect 9154 7932 9182 15826
rect 9730 15826 9854 15854
rect 9238 13753 9290 13759
rect 9238 13695 9290 13701
rect 8518 7907 8570 7913
rect 8518 7849 8570 7855
rect 9058 7904 9182 7932
rect 8530 7691 8558 7849
rect 8518 7685 8570 7691
rect 8518 7627 8570 7633
rect 8854 7019 8906 7025
rect 8854 6961 8906 6967
rect 8470 6575 8522 6581
rect 8470 6517 8522 6523
rect 8374 6427 8426 6433
rect 8374 6369 8426 6375
rect 8374 5465 8426 5471
rect 8374 5407 8426 5413
rect 8386 4879 8414 5407
rect 8374 4873 8426 4879
rect 8374 4815 8426 4821
rect 8278 3837 8330 3843
rect 8278 3779 8330 3785
rect 8182 3023 8234 3029
rect 8182 2965 8234 2971
rect 8194 800 8222 2965
rect 8290 800 8318 3779
rect 8482 800 8510 6517
rect 8758 5687 8810 5693
rect 8758 5629 8810 5635
rect 8770 4232 8798 5629
rect 8674 4204 8798 4232
rect 8566 3689 8618 3695
rect 8566 3631 8618 3637
rect 8578 800 8606 3631
rect 8674 800 8702 4204
rect 8758 3763 8810 3769
rect 8758 3705 8810 3711
rect 8770 2881 8798 3705
rect 8758 2875 8810 2881
rect 8758 2817 8810 2823
rect 8866 2752 8894 6961
rect 9058 6507 9086 7904
rect 9142 7759 9194 7765
rect 9142 7701 9194 7707
rect 9046 6501 9098 6507
rect 9046 6443 9098 6449
rect 9046 3911 9098 3917
rect 9046 3853 9098 3859
rect 8950 2949 9002 2955
rect 8950 2891 9002 2897
rect 8770 2724 8894 2752
rect 8770 800 8798 2724
rect 8962 800 8990 2891
rect 9058 800 9086 3853
rect 9154 800 9182 7701
rect 9250 6951 9278 13695
rect 9430 10127 9482 10133
rect 9430 10069 9482 10075
rect 9442 7691 9470 10069
rect 9730 8431 9758 15826
rect 9910 13679 9962 13685
rect 9910 13621 9962 13627
rect 9814 13457 9866 13463
rect 9814 13399 9866 13405
rect 9718 8425 9770 8431
rect 9718 8367 9770 8373
rect 9526 8277 9578 8283
rect 9526 8219 9578 8225
rect 9430 7685 9482 7691
rect 9430 7627 9482 7633
rect 9334 7463 9386 7469
rect 9334 7405 9386 7411
rect 9238 6945 9290 6951
rect 9238 6887 9290 6893
rect 9346 6581 9374 7405
rect 9334 6575 9386 6581
rect 9334 6517 9386 6523
rect 9430 6353 9482 6359
rect 9430 6295 9482 6301
rect 9238 5021 9290 5027
rect 9238 4963 9290 4969
rect 9250 4583 9278 4963
rect 9238 4577 9290 4583
rect 9238 4519 9290 4525
rect 9334 3689 9386 3695
rect 9334 3631 9386 3637
rect 9346 2894 9374 3631
rect 9250 2866 9374 2894
rect 9250 800 9278 2866
rect 9442 800 9470 6295
rect 9538 800 9566 8219
rect 9826 6951 9854 13399
rect 9922 12797 9950 13621
rect 9910 12791 9962 12797
rect 9910 12733 9962 12739
rect 10582 10867 10634 10873
rect 10582 10809 10634 10815
rect 10594 10503 10622 10809
rect 10582 10497 10634 10503
rect 10582 10439 10634 10445
rect 10786 9097 10814 56763
rect 11158 56229 11210 56235
rect 11158 56171 11210 56177
rect 10870 53861 10922 53867
rect 10870 53803 10922 53809
rect 10882 46541 10910 53803
rect 10966 48089 11018 48095
rect 10966 48031 11018 48037
rect 10870 46535 10922 46541
rect 10870 46477 10922 46483
rect 10870 26555 10922 26561
rect 10870 26497 10922 26503
rect 10882 10799 10910 26497
rect 10870 10793 10922 10799
rect 10870 10735 10922 10741
rect 10978 9837 11006 48031
rect 11170 38845 11198 56171
rect 11158 38839 11210 38845
rect 11158 38781 11210 38787
rect 11158 37433 11210 37439
rect 11158 37375 11210 37381
rect 11170 37217 11198 37375
rect 11158 37211 11210 37217
rect 11158 37153 11210 37159
rect 11062 25223 11114 25229
rect 11062 25165 11114 25171
rect 10966 9831 11018 9837
rect 10966 9773 11018 9779
rect 10774 9091 10826 9097
rect 10774 9033 10826 9039
rect 9910 8573 9962 8579
rect 9910 8515 9962 8521
rect 9922 8431 9950 8515
rect 9910 8425 9962 8431
rect 9910 8367 9962 8373
rect 10294 8277 10346 8283
rect 10294 8219 10346 8225
rect 10678 8277 10730 8283
rect 10678 8219 10730 8225
rect 9910 7537 9962 7543
rect 9910 7479 9962 7485
rect 9814 6945 9866 6951
rect 9814 6887 9866 6893
rect 9622 4355 9674 4361
rect 9622 4297 9674 4303
rect 9634 800 9662 4297
rect 9814 4281 9866 4287
rect 9814 4223 9866 4229
rect 9826 800 9854 4223
rect 9922 800 9950 7479
rect 10102 6353 10154 6359
rect 10102 6295 10154 6301
rect 10006 5021 10058 5027
rect 10006 4963 10058 4969
rect 10018 3843 10046 4963
rect 10006 3837 10058 3843
rect 10006 3779 10058 3785
rect 10006 3541 10058 3547
rect 10006 3483 10058 3489
rect 10018 800 10046 3483
rect 10114 800 10142 6295
rect 10198 5687 10250 5693
rect 10198 5629 10250 5635
rect 10210 4287 10238 5629
rect 10198 4281 10250 4287
rect 10198 4223 10250 4229
rect 10306 800 10334 8219
rect 10582 7167 10634 7173
rect 10582 7109 10634 7115
rect 10594 7025 10622 7109
rect 10582 7019 10634 7025
rect 10582 6961 10634 6967
rect 10486 5687 10538 5693
rect 10486 5629 10538 5635
rect 10390 4355 10442 4361
rect 10390 4297 10442 4303
rect 10402 800 10430 4297
rect 10498 800 10526 5629
rect 10582 5021 10634 5027
rect 10582 4963 10634 4969
rect 10594 3917 10622 4963
rect 10582 3911 10634 3917
rect 10582 3853 10634 3859
rect 10690 2894 10718 8219
rect 10966 7463 11018 7469
rect 10966 7405 11018 7411
rect 10870 6353 10922 6359
rect 10870 6295 10922 6301
rect 10774 4355 10826 4361
rect 10774 4297 10826 4303
rect 10594 2866 10718 2894
rect 10594 800 10622 2866
rect 10786 800 10814 4297
rect 10882 800 10910 6295
rect 10978 800 11006 7405
rect 11074 4435 11102 25165
rect 11158 10793 11210 10799
rect 11158 10735 11210 10741
rect 11170 4583 11198 10735
rect 11266 7913 11294 56837
rect 11746 56531 11774 59200
rect 12322 56531 12350 59200
rect 12802 56975 12830 59200
rect 12790 56969 12842 56975
rect 12790 56911 12842 56917
rect 12982 56895 13034 56901
rect 12982 56837 13034 56843
rect 11734 56525 11786 56531
rect 11734 56467 11786 56473
rect 12310 56525 12362 56531
rect 12310 56467 12362 56473
rect 11446 56377 11498 56383
rect 11446 56319 11498 56325
rect 12214 56377 12266 56383
rect 12214 56319 12266 56325
rect 11458 55051 11486 56319
rect 11926 56229 11978 56235
rect 11926 56171 11978 56177
rect 11938 55791 11966 56171
rect 11926 55785 11978 55791
rect 11926 55727 11978 55733
rect 11446 55045 11498 55051
rect 11446 54987 11498 54993
rect 11350 38469 11402 38475
rect 11350 38411 11402 38417
rect 11362 8431 11390 38411
rect 12118 26481 12170 26487
rect 12118 26423 12170 26429
rect 12022 25519 12074 25525
rect 12022 25461 12074 25467
rect 11350 8425 11402 8431
rect 11350 8367 11402 8373
rect 11446 8277 11498 8283
rect 11446 8219 11498 8225
rect 11254 7907 11306 7913
rect 11254 7849 11306 7855
rect 11254 7019 11306 7025
rect 11254 6961 11306 6967
rect 11158 4577 11210 4583
rect 11158 4519 11210 4525
rect 11062 4429 11114 4435
rect 11062 4371 11114 4377
rect 11158 4207 11210 4213
rect 11158 4149 11210 4155
rect 11170 800 11198 4149
rect 11266 800 11294 6961
rect 11458 5774 11486 8219
rect 11734 7759 11786 7765
rect 11734 7701 11786 7707
rect 11638 6353 11690 6359
rect 11638 6295 11690 6301
rect 11362 5746 11486 5774
rect 11362 800 11390 5746
rect 11446 4281 11498 4287
rect 11446 4223 11498 4229
rect 11458 800 11486 4223
rect 11650 800 11678 6295
rect 11746 800 11774 7701
rect 12034 7691 12062 25461
rect 12022 7685 12074 7691
rect 12022 7627 12074 7633
rect 11830 5021 11882 5027
rect 11830 4963 11882 4969
rect 11842 800 11870 4963
rect 12130 4509 12158 26423
rect 12226 9467 12254 56319
rect 12694 56229 12746 56235
rect 12694 56171 12746 56177
rect 12310 43427 12362 43433
rect 12310 43369 12362 43375
rect 12214 9461 12266 9467
rect 12214 9403 12266 9409
rect 12214 8277 12266 8283
rect 12214 8219 12266 8225
rect 12118 4503 12170 4509
rect 12118 4445 12170 4451
rect 12022 3467 12074 3473
rect 12022 3409 12074 3415
rect 12034 800 12062 3409
rect 12226 2308 12254 8219
rect 12322 7617 12350 43369
rect 12598 38765 12650 38771
rect 12598 38707 12650 38713
rect 12610 38549 12638 38707
rect 12598 38543 12650 38549
rect 12598 38485 12650 38491
rect 12706 34849 12734 56171
rect 12790 55563 12842 55569
rect 12790 55505 12842 55511
rect 12694 34843 12746 34849
rect 12694 34785 12746 34791
rect 12598 34769 12650 34775
rect 12598 34711 12650 34717
rect 12502 33585 12554 33591
rect 12502 33527 12554 33533
rect 12514 15854 12542 33527
rect 12418 15826 12542 15854
rect 12310 7611 12362 7617
rect 12310 7553 12362 7559
rect 12418 7173 12446 15826
rect 12502 12273 12554 12279
rect 12502 12215 12554 12221
rect 12514 7691 12542 12215
rect 12610 8579 12638 34711
rect 12694 27887 12746 27893
rect 12694 27829 12746 27835
rect 12706 8949 12734 27829
rect 12802 12279 12830 55505
rect 12790 12273 12842 12279
rect 12790 12215 12842 12221
rect 12886 10423 12938 10429
rect 12886 10365 12938 10371
rect 12694 8943 12746 8949
rect 12694 8885 12746 8891
rect 12598 8573 12650 8579
rect 12598 8515 12650 8521
rect 12790 8573 12842 8579
rect 12790 8515 12842 8521
rect 12502 7685 12554 7691
rect 12502 7627 12554 7633
rect 12502 7463 12554 7469
rect 12502 7405 12554 7411
rect 12406 7167 12458 7173
rect 12406 7109 12458 7115
rect 12310 6945 12362 6951
rect 12310 6887 12362 6893
rect 12322 3917 12350 6887
rect 12406 6353 12458 6359
rect 12406 6295 12458 6301
rect 12310 3911 12362 3917
rect 12310 3853 12362 3859
rect 12310 3171 12362 3177
rect 12310 3113 12362 3119
rect 12130 2280 12254 2308
rect 12130 800 12158 2280
rect 12322 2160 12350 3113
rect 12226 2132 12350 2160
rect 12226 800 12254 2132
rect 12418 2012 12446 6295
rect 12322 1984 12446 2012
rect 12322 800 12350 1984
rect 12514 800 12542 7405
rect 12694 7019 12746 7025
rect 12694 6961 12746 6967
rect 12598 5687 12650 5693
rect 12598 5629 12650 5635
rect 12610 800 12638 5629
rect 12706 800 12734 6961
rect 12802 800 12830 8515
rect 12898 6951 12926 10365
rect 12994 7807 13022 56837
rect 13378 56531 13406 59200
rect 13654 56895 13706 56901
rect 13654 56837 13706 56843
rect 13666 56753 13694 56837
rect 13654 56747 13706 56753
rect 13654 56689 13706 56695
rect 13366 56525 13418 56531
rect 13366 56467 13418 56473
rect 13270 56229 13322 56235
rect 13270 56171 13322 56177
rect 13078 35583 13130 35589
rect 13078 35525 13130 35531
rect 13090 35441 13118 35525
rect 13078 35435 13130 35441
rect 13078 35377 13130 35383
rect 13090 12427 13118 35377
rect 13282 29669 13310 56171
rect 13270 29663 13322 29669
rect 13270 29605 13322 29611
rect 13270 23521 13322 23527
rect 13270 23463 13322 23469
rect 13174 23225 13226 23231
rect 13174 23167 13226 23173
rect 13078 12421 13130 12427
rect 13078 12363 13130 12369
rect 12980 7798 13036 7807
rect 12980 7733 13036 7742
rect 12886 6945 12938 6951
rect 12886 6887 12938 6893
rect 13078 6427 13130 6433
rect 13078 6369 13130 6375
rect 12982 5021 13034 5027
rect 12982 4963 13034 4969
rect 12994 3177 13022 4963
rect 12982 3171 13034 3177
rect 12982 3113 13034 3119
rect 12982 3023 13034 3029
rect 12982 2965 13034 2971
rect 12994 800 13022 2965
rect 13090 800 13118 6369
rect 13186 3917 13214 23167
rect 13174 3911 13226 3917
rect 13174 3853 13226 3859
rect 13174 3689 13226 3695
rect 13174 3631 13226 3637
rect 13186 800 13214 3631
rect 13282 3251 13310 23463
rect 13558 16565 13610 16571
rect 13558 16507 13610 16513
rect 13570 8431 13598 16507
rect 13666 15239 13694 56689
rect 13858 55717 13886 59200
rect 14434 56975 14462 59200
rect 14422 56969 14474 56975
rect 14422 56911 14474 56917
rect 14914 56531 14942 59200
rect 14902 56525 14954 56531
rect 14902 56467 14954 56473
rect 15094 56229 15146 56235
rect 15094 56171 15146 56177
rect 13846 55711 13898 55717
rect 13846 55653 13898 55659
rect 13750 33215 13802 33221
rect 13750 33157 13802 33163
rect 13654 15233 13706 15239
rect 13654 15175 13706 15181
rect 13558 8425 13610 8431
rect 13558 8367 13610 8373
rect 13762 8357 13790 33157
rect 14422 28331 14474 28337
rect 14422 28273 14474 28279
rect 14434 27893 14462 28273
rect 14422 27887 14474 27893
rect 14422 27829 14474 27835
rect 14134 24557 14186 24563
rect 14134 24499 14186 24505
rect 14038 23151 14090 23157
rect 14038 23093 14090 23099
rect 13942 9239 13994 9245
rect 13942 9181 13994 9187
rect 13750 8351 13802 8357
rect 13750 8293 13802 8299
rect 13462 6945 13514 6951
rect 13462 6887 13514 6893
rect 13750 6945 13802 6951
rect 13750 6887 13802 6893
rect 13366 5687 13418 5693
rect 13366 5629 13418 5635
rect 13378 3473 13406 5629
rect 13366 3467 13418 3473
rect 13366 3409 13418 3415
rect 13270 3245 13322 3251
rect 13270 3187 13322 3193
rect 13366 3023 13418 3029
rect 13366 2965 13418 2971
rect 13378 800 13406 2965
rect 13474 800 13502 6887
rect 13558 4355 13610 4361
rect 13558 4297 13610 4303
rect 13570 800 13598 4297
rect 13654 3689 13706 3695
rect 13654 3631 13706 3637
rect 13666 800 13694 3631
rect 13762 2585 13790 6887
rect 13954 6433 13982 9181
rect 13942 6427 13994 6433
rect 13942 6369 13994 6375
rect 13942 5021 13994 5027
rect 13942 4963 13994 4969
rect 13846 3171 13898 3177
rect 13846 3113 13898 3119
rect 13750 2579 13802 2585
rect 13750 2521 13802 2527
rect 13858 800 13886 3113
rect 13954 800 13982 4963
rect 14050 3251 14078 23093
rect 14146 3917 14174 24499
rect 15106 17015 15134 56171
rect 15394 56161 15422 59200
rect 15970 56975 15998 59200
rect 16450 57049 16478 59200
rect 16438 57043 16490 57049
rect 16438 56985 16490 56991
rect 15958 56969 16010 56975
rect 15958 56911 16010 56917
rect 16150 56895 16202 56901
rect 16150 56837 16202 56843
rect 15382 56155 15434 56161
rect 15382 56097 15434 56103
rect 15958 33437 16010 33443
rect 15958 33379 16010 33385
rect 15478 23817 15530 23823
rect 15478 23759 15530 23765
rect 15094 17009 15146 17015
rect 15094 16951 15146 16957
rect 15094 13457 15146 13463
rect 15094 13399 15146 13405
rect 15106 13241 15134 13399
rect 15094 13235 15146 13241
rect 15094 13177 15146 13183
rect 15190 12125 15242 12131
rect 15190 12067 15242 12073
rect 15202 11909 15230 12067
rect 15190 11903 15242 11909
rect 15190 11845 15242 11851
rect 15094 9535 15146 9541
rect 15094 9477 15146 9483
rect 15106 7691 15134 9477
rect 15094 7685 15146 7691
rect 15094 7627 15146 7633
rect 14614 6945 14666 6951
rect 14614 6887 14666 6893
rect 15382 6945 15434 6951
rect 15382 6887 15434 6893
rect 14230 6205 14282 6211
rect 14230 6147 14282 6153
rect 14134 3911 14186 3917
rect 14134 3853 14186 3859
rect 14134 3689 14186 3695
rect 14134 3631 14186 3637
rect 14038 3245 14090 3251
rect 14038 3187 14090 3193
rect 14146 1272 14174 3631
rect 14050 1244 14174 1272
rect 14050 800 14078 1244
rect 14242 1124 14270 6147
rect 14518 6131 14570 6137
rect 14518 6073 14570 6079
rect 14422 5021 14474 5027
rect 14422 4963 14474 4969
rect 14434 2900 14462 4963
rect 14530 3177 14558 6073
rect 14518 3171 14570 3177
rect 14518 3113 14570 3119
rect 14518 3023 14570 3029
rect 14518 2965 14570 2971
rect 14146 1096 14270 1124
rect 14338 2872 14462 2900
rect 14146 800 14174 1096
rect 14338 800 14366 2872
rect 14530 1568 14558 2965
rect 14434 1540 14558 1568
rect 14434 800 14462 1540
rect 14626 1420 14654 6887
rect 14998 5687 15050 5693
rect 14998 5629 15050 5635
rect 14806 5021 14858 5027
rect 14530 1392 14654 1420
rect 14722 4981 14806 5009
rect 14530 800 14558 1392
rect 14722 800 14750 4981
rect 14806 4963 14858 4969
rect 14902 4281 14954 4287
rect 14902 4223 14954 4229
rect 14806 3689 14858 3695
rect 14806 3631 14858 3637
rect 14818 800 14846 3631
rect 14914 800 14942 4223
rect 15010 800 15038 5629
rect 15094 4429 15146 4435
rect 15094 4371 15146 4377
rect 15106 3251 15134 4371
rect 15286 3689 15338 3695
rect 15202 3649 15286 3677
rect 15094 3245 15146 3251
rect 15094 3187 15146 3193
rect 15202 800 15230 3649
rect 15286 3631 15338 3637
rect 15394 3492 15422 6887
rect 15490 6433 15518 23759
rect 15862 12199 15914 12205
rect 15862 12141 15914 12147
rect 15874 7691 15902 12141
rect 15862 7685 15914 7691
rect 15862 7627 15914 7633
rect 15670 7463 15722 7469
rect 15670 7405 15722 7411
rect 15862 7463 15914 7469
rect 15862 7405 15914 7411
rect 15478 6427 15530 6433
rect 15478 6369 15530 6375
rect 15478 4355 15530 4361
rect 15478 4297 15530 4303
rect 15298 3464 15422 3492
rect 15298 800 15326 3464
rect 15382 2949 15434 2955
rect 15382 2891 15434 2897
rect 15394 800 15422 2891
rect 15490 800 15518 4297
rect 15682 800 15710 7405
rect 15874 7099 15902 7405
rect 15862 7093 15914 7099
rect 15862 7035 15914 7041
rect 15970 6581 15998 33379
rect 16054 11237 16106 11243
rect 16054 11179 16106 11185
rect 16066 9560 16094 11179
rect 16162 9689 16190 56837
rect 17026 56531 17054 59200
rect 17506 56975 17534 59200
rect 17494 56969 17546 56975
rect 17494 56911 17546 56917
rect 17974 56895 18026 56901
rect 17974 56837 18026 56843
rect 17014 56525 17066 56531
rect 17014 56467 17066 56473
rect 17206 56229 17258 56235
rect 17206 56171 17258 56177
rect 16534 55563 16586 55569
rect 16534 55505 16586 55511
rect 16438 36101 16490 36107
rect 16438 36043 16490 36049
rect 16246 30329 16298 30335
rect 16246 30271 16298 30277
rect 16258 10207 16286 30271
rect 16246 10201 16298 10207
rect 16246 10143 16298 10149
rect 16150 9683 16202 9689
rect 16150 9625 16202 9631
rect 16066 9532 16190 9560
rect 16054 8277 16106 8283
rect 16054 8219 16106 8225
rect 15958 6575 16010 6581
rect 15958 6517 16010 6523
rect 15766 6279 15818 6285
rect 15766 6221 15818 6227
rect 15778 3917 15806 6221
rect 15862 5687 15914 5693
rect 15862 5629 15914 5635
rect 15766 3911 15818 3917
rect 15766 3853 15818 3859
rect 15874 2900 15902 5629
rect 15958 4355 16010 4361
rect 15958 4297 16010 4303
rect 15778 2872 15902 2900
rect 15778 800 15806 2872
rect 15970 2160 15998 4297
rect 15874 2132 15998 2160
rect 15874 800 15902 2132
rect 16066 800 16094 8219
rect 16162 7469 16190 9532
rect 16450 9171 16478 36043
rect 16546 9467 16574 55505
rect 17110 44093 17162 44099
rect 17110 44035 17162 44041
rect 16822 27443 16874 27449
rect 16822 27385 16874 27391
rect 16726 20117 16778 20123
rect 16726 20059 16778 20065
rect 16738 19827 16766 20059
rect 16726 19821 16778 19827
rect 16726 19763 16778 19769
rect 16534 9461 16586 9467
rect 16534 9403 16586 9409
rect 16438 9165 16490 9171
rect 16438 9107 16490 9113
rect 16246 8869 16298 8875
rect 16246 8811 16298 8817
rect 16258 8431 16286 8811
rect 16246 8425 16298 8431
rect 16246 8367 16298 8373
rect 16342 8277 16394 8283
rect 16342 8219 16394 8225
rect 16246 8129 16298 8135
rect 16246 8071 16298 8077
rect 16150 7463 16202 7469
rect 16150 7405 16202 7411
rect 16258 6803 16286 8071
rect 16246 6797 16298 6803
rect 16246 6739 16298 6745
rect 16150 5687 16202 5693
rect 16150 5629 16202 5635
rect 16162 800 16190 5629
rect 16246 4207 16298 4213
rect 16246 4149 16298 4155
rect 16258 800 16286 4149
rect 16354 800 16382 8219
rect 16534 6131 16586 6137
rect 16534 6073 16586 6079
rect 16438 5021 16490 5027
rect 16438 4963 16490 4969
rect 16450 2955 16478 4963
rect 16546 4287 16574 6073
rect 16534 4281 16586 4287
rect 16534 4223 16586 4229
rect 16534 3837 16586 3843
rect 16534 3779 16586 3785
rect 16438 2949 16490 2955
rect 16438 2891 16490 2897
rect 16546 800 16574 3779
rect 16834 3251 16862 27385
rect 17014 26111 17066 26117
rect 17014 26053 17066 26059
rect 17026 8431 17054 26053
rect 17122 10133 17150 44035
rect 17218 41435 17246 56171
rect 17206 41429 17258 41435
rect 17206 41371 17258 41377
rect 17878 29515 17930 29521
rect 17878 29457 17930 29463
rect 17782 14937 17834 14943
rect 17782 14879 17834 14885
rect 17794 14425 17822 14879
rect 17782 14419 17834 14425
rect 17782 14361 17834 14367
rect 17110 10127 17162 10133
rect 17110 10069 17162 10075
rect 17302 9683 17354 9689
rect 17302 9625 17354 9631
rect 17014 8425 17066 8431
rect 17014 8367 17066 8373
rect 17314 7099 17342 9625
rect 17686 9091 17738 9097
rect 17686 9033 17738 9039
rect 17302 7093 17354 7099
rect 17302 7035 17354 7041
rect 17110 6945 17162 6951
rect 17110 6887 17162 6893
rect 16918 4133 16970 4139
rect 16918 4075 16970 4081
rect 16822 3245 16874 3251
rect 16822 3187 16874 3193
rect 16726 3097 16778 3103
rect 16726 3039 16778 3045
rect 16630 3023 16682 3029
rect 16630 2965 16682 2971
rect 16642 800 16670 2965
rect 16738 800 16766 3039
rect 16930 800 16958 4075
rect 17014 3023 17066 3029
rect 17014 2965 17066 2971
rect 17026 800 17054 2965
rect 17122 800 17150 6887
rect 17698 6433 17726 9033
rect 17890 7214 17918 29457
rect 17986 9911 18014 56837
rect 18082 56531 18110 59200
rect 18562 56531 18590 59200
rect 19138 56975 19166 59200
rect 19618 57614 19646 59200
rect 19618 57586 20030 57614
rect 19126 56969 19178 56975
rect 19126 56911 19178 56917
rect 19318 56895 19370 56901
rect 19318 56837 19370 56843
rect 18070 56525 18122 56531
rect 18070 56467 18122 56473
rect 18550 56525 18602 56531
rect 18550 56467 18602 56473
rect 18262 56229 18314 56235
rect 18262 56171 18314 56177
rect 18274 42175 18302 56171
rect 19126 46831 19178 46837
rect 19126 46773 19178 46779
rect 18262 42169 18314 42175
rect 18262 42111 18314 42117
rect 18838 29589 18890 29595
rect 18838 29531 18890 29537
rect 18358 29441 18410 29447
rect 18358 29383 18410 29389
rect 18070 28183 18122 28189
rect 18070 28125 18122 28131
rect 17974 9905 18026 9911
rect 17974 9847 18026 9853
rect 17794 7186 17918 7214
rect 17686 6427 17738 6433
rect 17686 6369 17738 6375
rect 17590 6131 17642 6137
rect 17590 6073 17642 6079
rect 17302 5687 17354 5693
rect 17302 5629 17354 5635
rect 17206 4133 17258 4139
rect 17206 4075 17258 4081
rect 17218 3917 17246 4075
rect 17206 3911 17258 3917
rect 17206 3853 17258 3859
rect 17314 3843 17342 5629
rect 17494 5021 17546 5027
rect 17494 4963 17546 4969
rect 17302 3837 17354 3843
rect 17302 3779 17354 3785
rect 17398 3689 17450 3695
rect 17398 3631 17450 3637
rect 17302 3541 17354 3547
rect 17302 3483 17354 3489
rect 17314 2900 17342 3483
rect 17218 2872 17342 2900
rect 17218 800 17246 2872
rect 17410 800 17438 3631
rect 17506 3547 17534 4963
rect 17494 3541 17546 3547
rect 17494 3483 17546 3489
rect 17494 3171 17546 3177
rect 17494 3113 17546 3119
rect 17506 800 17534 3113
rect 17602 3103 17630 6073
rect 17686 4281 17738 4287
rect 17686 4223 17738 4229
rect 17590 3097 17642 3103
rect 17590 3039 17642 3045
rect 17698 3011 17726 4223
rect 17794 3917 17822 7186
rect 17878 6945 17930 6951
rect 17878 6887 17930 6893
rect 17782 3911 17834 3917
rect 17782 3853 17834 3859
rect 17602 2983 17726 3011
rect 17602 800 17630 2983
rect 17686 2949 17738 2955
rect 17686 2891 17738 2897
rect 17698 800 17726 2891
rect 17890 800 17918 6887
rect 17974 5021 18026 5027
rect 17974 4963 18026 4969
rect 17986 800 18014 4963
rect 18082 3251 18110 28125
rect 18166 26851 18218 26857
rect 18166 26793 18218 26799
rect 18178 8875 18206 26793
rect 18370 9911 18398 29383
rect 18742 12125 18794 12131
rect 18742 12067 18794 12073
rect 18358 9905 18410 9911
rect 18358 9847 18410 9853
rect 18262 9609 18314 9615
rect 18262 9551 18314 9557
rect 18166 8869 18218 8875
rect 18166 8811 18218 8817
rect 18274 7099 18302 9551
rect 18454 8943 18506 8949
rect 18454 8885 18506 8891
rect 18262 7093 18314 7099
rect 18262 7035 18314 7041
rect 18466 6433 18494 8885
rect 18550 6945 18602 6951
rect 18550 6887 18602 6893
rect 18454 6427 18506 6433
rect 18454 6369 18506 6375
rect 18262 6131 18314 6137
rect 18262 6073 18314 6079
rect 18166 3689 18218 3695
rect 18166 3631 18218 3637
rect 18070 3245 18122 3251
rect 18070 3187 18122 3193
rect 18178 1864 18206 3631
rect 18274 3177 18302 6073
rect 18454 3689 18506 3695
rect 18454 3631 18506 3637
rect 18262 3171 18314 3177
rect 18262 3113 18314 3119
rect 18358 3097 18410 3103
rect 18358 3039 18410 3045
rect 18262 2875 18314 2881
rect 18262 2817 18314 2823
rect 18082 1836 18206 1864
rect 18082 800 18110 1836
rect 18274 800 18302 2817
rect 18370 800 18398 3039
rect 18466 800 18494 3631
rect 18562 800 18590 6887
rect 18754 6359 18782 12067
rect 18742 6353 18794 6359
rect 18742 6295 18794 6301
rect 18742 5687 18794 5693
rect 18742 5629 18794 5635
rect 18754 800 18782 5629
rect 18850 3251 18878 29531
rect 18934 28553 18986 28559
rect 18934 28495 18986 28501
rect 18946 7099 18974 28495
rect 18934 7093 18986 7099
rect 18934 7035 18986 7041
rect 19138 6433 19166 46773
rect 19330 9023 19358 56837
rect 19628 56638 19924 56658
rect 19684 56636 19708 56638
rect 19764 56636 19788 56638
rect 19844 56636 19868 56638
rect 19706 56584 19708 56636
rect 19770 56584 19782 56636
rect 19844 56584 19846 56636
rect 19684 56582 19708 56584
rect 19764 56582 19788 56584
rect 19844 56582 19868 56584
rect 19628 56562 19924 56582
rect 20002 56531 20030 57586
rect 19990 56525 20042 56531
rect 19990 56467 20042 56473
rect 20194 55717 20222 59200
rect 20674 56975 20702 59200
rect 20662 56969 20714 56975
rect 20662 56911 20714 56917
rect 21250 56531 21278 59200
rect 21730 56531 21758 59200
rect 22306 56975 22334 59200
rect 22294 56969 22346 56975
rect 22294 56911 22346 56917
rect 22786 56531 22814 59200
rect 21238 56525 21290 56531
rect 21238 56467 21290 56473
rect 21718 56525 21770 56531
rect 21718 56467 21770 56473
rect 22774 56525 22826 56531
rect 22774 56467 22826 56473
rect 20374 56229 20426 56235
rect 20374 56171 20426 56177
rect 21430 56229 21482 56235
rect 21430 56171 21482 56177
rect 22198 56229 22250 56235
rect 22198 56171 22250 56177
rect 22966 56229 23018 56235
rect 22966 56171 23018 56177
rect 20182 55711 20234 55717
rect 20182 55653 20234 55659
rect 20278 55563 20330 55569
rect 20278 55505 20330 55511
rect 19628 55306 19924 55326
rect 19684 55304 19708 55306
rect 19764 55304 19788 55306
rect 19844 55304 19868 55306
rect 19706 55252 19708 55304
rect 19770 55252 19782 55304
rect 19844 55252 19846 55304
rect 19684 55250 19708 55252
rect 19764 55250 19788 55252
rect 19844 55250 19868 55252
rect 19628 55230 19924 55250
rect 19990 55193 20042 55199
rect 19990 55135 20042 55141
rect 19628 53974 19924 53994
rect 19684 53972 19708 53974
rect 19764 53972 19788 53974
rect 19844 53972 19868 53974
rect 19706 53920 19708 53972
rect 19770 53920 19782 53972
rect 19844 53920 19846 53972
rect 19684 53918 19708 53920
rect 19764 53918 19788 53920
rect 19844 53918 19868 53920
rect 19628 53898 19924 53918
rect 19628 52642 19924 52662
rect 19684 52640 19708 52642
rect 19764 52640 19788 52642
rect 19844 52640 19868 52642
rect 19706 52588 19708 52640
rect 19770 52588 19782 52640
rect 19844 52588 19846 52640
rect 19684 52586 19708 52588
rect 19764 52586 19788 52588
rect 19844 52586 19868 52588
rect 19628 52566 19924 52586
rect 19628 51310 19924 51330
rect 19684 51308 19708 51310
rect 19764 51308 19788 51310
rect 19844 51308 19868 51310
rect 19706 51256 19708 51308
rect 19770 51256 19782 51308
rect 19844 51256 19846 51308
rect 19684 51254 19708 51256
rect 19764 51254 19788 51256
rect 19844 51254 19868 51256
rect 19628 51234 19924 51254
rect 19628 49978 19924 49998
rect 19684 49976 19708 49978
rect 19764 49976 19788 49978
rect 19844 49976 19868 49978
rect 19706 49924 19708 49976
rect 19770 49924 19782 49976
rect 19844 49924 19846 49976
rect 19684 49922 19708 49924
rect 19764 49922 19788 49924
rect 19844 49922 19868 49924
rect 19628 49902 19924 49922
rect 19628 48646 19924 48666
rect 19684 48644 19708 48646
rect 19764 48644 19788 48646
rect 19844 48644 19868 48646
rect 19706 48592 19708 48644
rect 19770 48592 19782 48644
rect 19844 48592 19846 48644
rect 19684 48590 19708 48592
rect 19764 48590 19788 48592
rect 19844 48590 19868 48592
rect 19628 48570 19924 48590
rect 19628 47314 19924 47334
rect 19684 47312 19708 47314
rect 19764 47312 19788 47314
rect 19844 47312 19868 47314
rect 19706 47260 19708 47312
rect 19770 47260 19782 47312
rect 19844 47260 19846 47312
rect 19684 47258 19708 47260
rect 19764 47258 19788 47260
rect 19844 47258 19868 47260
rect 19628 47238 19924 47258
rect 19628 45982 19924 46002
rect 19684 45980 19708 45982
rect 19764 45980 19788 45982
rect 19844 45980 19868 45982
rect 19706 45928 19708 45980
rect 19770 45928 19782 45980
rect 19844 45928 19846 45980
rect 19684 45926 19708 45928
rect 19764 45926 19788 45928
rect 19844 45926 19868 45928
rect 19628 45906 19924 45926
rect 19628 44650 19924 44670
rect 19684 44648 19708 44650
rect 19764 44648 19788 44650
rect 19844 44648 19868 44650
rect 19706 44596 19708 44648
rect 19770 44596 19782 44648
rect 19844 44596 19846 44648
rect 19684 44594 19708 44596
rect 19764 44594 19788 44596
rect 19844 44594 19868 44596
rect 19628 44574 19924 44594
rect 19628 43318 19924 43338
rect 19684 43316 19708 43318
rect 19764 43316 19788 43318
rect 19844 43316 19868 43318
rect 19706 43264 19708 43316
rect 19770 43264 19782 43316
rect 19844 43264 19846 43316
rect 19684 43262 19708 43264
rect 19764 43262 19788 43264
rect 19844 43262 19868 43264
rect 19628 43242 19924 43262
rect 19628 41986 19924 42006
rect 19684 41984 19708 41986
rect 19764 41984 19788 41986
rect 19844 41984 19868 41986
rect 19706 41932 19708 41984
rect 19770 41932 19782 41984
rect 19844 41932 19846 41984
rect 19684 41930 19708 41932
rect 19764 41930 19788 41932
rect 19844 41930 19868 41932
rect 19628 41910 19924 41930
rect 19628 40654 19924 40674
rect 19684 40652 19708 40654
rect 19764 40652 19788 40654
rect 19844 40652 19868 40654
rect 19706 40600 19708 40652
rect 19770 40600 19782 40652
rect 19844 40600 19846 40652
rect 19684 40598 19708 40600
rect 19764 40598 19788 40600
rect 19844 40598 19868 40600
rect 19628 40578 19924 40598
rect 19628 39322 19924 39342
rect 19684 39320 19708 39322
rect 19764 39320 19788 39322
rect 19844 39320 19868 39322
rect 19706 39268 19708 39320
rect 19770 39268 19782 39320
rect 19844 39268 19846 39320
rect 19684 39266 19708 39268
rect 19764 39266 19788 39268
rect 19844 39266 19868 39268
rect 19628 39246 19924 39266
rect 19628 37990 19924 38010
rect 19684 37988 19708 37990
rect 19764 37988 19788 37990
rect 19844 37988 19868 37990
rect 19706 37936 19708 37988
rect 19770 37936 19782 37988
rect 19844 37936 19846 37988
rect 19684 37934 19708 37936
rect 19764 37934 19788 37936
rect 19844 37934 19868 37936
rect 19628 37914 19924 37934
rect 19628 36658 19924 36678
rect 19684 36656 19708 36658
rect 19764 36656 19788 36658
rect 19844 36656 19868 36658
rect 19706 36604 19708 36656
rect 19770 36604 19782 36656
rect 19844 36604 19846 36656
rect 19684 36602 19708 36604
rect 19764 36602 19788 36604
rect 19844 36602 19868 36604
rect 19628 36582 19924 36602
rect 19628 35326 19924 35346
rect 19684 35324 19708 35326
rect 19764 35324 19788 35326
rect 19844 35324 19868 35326
rect 19706 35272 19708 35324
rect 19770 35272 19782 35324
rect 19844 35272 19846 35324
rect 19684 35270 19708 35272
rect 19764 35270 19788 35272
rect 19844 35270 19868 35272
rect 19628 35250 19924 35270
rect 19628 33994 19924 34014
rect 19684 33992 19708 33994
rect 19764 33992 19788 33994
rect 19844 33992 19868 33994
rect 19706 33940 19708 33992
rect 19770 33940 19782 33992
rect 19844 33940 19846 33992
rect 19684 33938 19708 33940
rect 19764 33938 19788 33940
rect 19844 33938 19868 33940
rect 19628 33918 19924 33938
rect 19628 32662 19924 32682
rect 19684 32660 19708 32662
rect 19764 32660 19788 32662
rect 19844 32660 19868 32662
rect 19706 32608 19708 32660
rect 19770 32608 19782 32660
rect 19844 32608 19846 32660
rect 19684 32606 19708 32608
rect 19764 32606 19788 32608
rect 19844 32606 19868 32608
rect 19628 32586 19924 32606
rect 19628 31330 19924 31350
rect 19684 31328 19708 31330
rect 19764 31328 19788 31330
rect 19844 31328 19868 31330
rect 19706 31276 19708 31328
rect 19770 31276 19782 31328
rect 19844 31276 19846 31328
rect 19684 31274 19708 31276
rect 19764 31274 19788 31276
rect 19844 31274 19868 31276
rect 19628 31254 19924 31274
rect 19628 29998 19924 30018
rect 19684 29996 19708 29998
rect 19764 29996 19788 29998
rect 19844 29996 19868 29998
rect 19706 29944 19708 29996
rect 19770 29944 19782 29996
rect 19844 29944 19846 29996
rect 19684 29942 19708 29944
rect 19764 29942 19788 29944
rect 19844 29942 19868 29944
rect 19628 29922 19924 29942
rect 19628 28666 19924 28686
rect 19684 28664 19708 28666
rect 19764 28664 19788 28666
rect 19844 28664 19868 28666
rect 19706 28612 19708 28664
rect 19770 28612 19782 28664
rect 19844 28612 19846 28664
rect 19684 28610 19708 28612
rect 19764 28610 19788 28612
rect 19844 28610 19868 28612
rect 19628 28590 19924 28610
rect 19628 27334 19924 27354
rect 19684 27332 19708 27334
rect 19764 27332 19788 27334
rect 19844 27332 19868 27334
rect 19706 27280 19708 27332
rect 19770 27280 19782 27332
rect 19844 27280 19846 27332
rect 19684 27278 19708 27280
rect 19764 27278 19788 27280
rect 19844 27278 19868 27280
rect 19628 27258 19924 27278
rect 19628 26002 19924 26022
rect 19684 26000 19708 26002
rect 19764 26000 19788 26002
rect 19844 26000 19868 26002
rect 19706 25948 19708 26000
rect 19770 25948 19782 26000
rect 19844 25948 19846 26000
rect 19684 25946 19708 25948
rect 19764 25946 19788 25948
rect 19844 25946 19868 25948
rect 19628 25926 19924 25946
rect 19628 24670 19924 24690
rect 19684 24668 19708 24670
rect 19764 24668 19788 24670
rect 19844 24668 19868 24670
rect 19706 24616 19708 24668
rect 19770 24616 19782 24668
rect 19844 24616 19846 24668
rect 19684 24614 19708 24616
rect 19764 24614 19788 24616
rect 19844 24614 19868 24616
rect 19628 24594 19924 24614
rect 19628 23338 19924 23358
rect 19684 23336 19708 23338
rect 19764 23336 19788 23338
rect 19844 23336 19868 23338
rect 19706 23284 19708 23336
rect 19770 23284 19782 23336
rect 19844 23284 19846 23336
rect 19684 23282 19708 23284
rect 19764 23282 19788 23284
rect 19844 23282 19868 23284
rect 19628 23262 19924 23282
rect 19628 22006 19924 22026
rect 19684 22004 19708 22006
rect 19764 22004 19788 22006
rect 19844 22004 19868 22006
rect 19706 21952 19708 22004
rect 19770 21952 19782 22004
rect 19844 21952 19846 22004
rect 19684 21950 19708 21952
rect 19764 21950 19788 21952
rect 19844 21950 19868 21952
rect 19628 21930 19924 21950
rect 19628 20674 19924 20694
rect 19684 20672 19708 20674
rect 19764 20672 19788 20674
rect 19844 20672 19868 20674
rect 19706 20620 19708 20672
rect 19770 20620 19782 20672
rect 19844 20620 19846 20672
rect 19684 20618 19708 20620
rect 19764 20618 19788 20620
rect 19844 20618 19868 20620
rect 19628 20598 19924 20618
rect 19628 19342 19924 19362
rect 19684 19340 19708 19342
rect 19764 19340 19788 19342
rect 19844 19340 19868 19342
rect 19706 19288 19708 19340
rect 19770 19288 19782 19340
rect 19844 19288 19846 19340
rect 19684 19286 19708 19288
rect 19764 19286 19788 19288
rect 19844 19286 19868 19288
rect 19628 19266 19924 19286
rect 19628 18010 19924 18030
rect 19684 18008 19708 18010
rect 19764 18008 19788 18010
rect 19844 18008 19868 18010
rect 19706 17956 19708 18008
rect 19770 17956 19782 18008
rect 19844 17956 19846 18008
rect 19684 17954 19708 17956
rect 19764 17954 19788 17956
rect 19844 17954 19868 17956
rect 19628 17934 19924 17954
rect 19628 16678 19924 16698
rect 19684 16676 19708 16678
rect 19764 16676 19788 16678
rect 19844 16676 19868 16678
rect 19706 16624 19708 16676
rect 19770 16624 19782 16676
rect 19844 16624 19846 16676
rect 19684 16622 19708 16624
rect 19764 16622 19788 16624
rect 19844 16622 19868 16624
rect 19628 16602 19924 16622
rect 19628 15346 19924 15366
rect 19684 15344 19708 15346
rect 19764 15344 19788 15346
rect 19844 15344 19868 15346
rect 19706 15292 19708 15344
rect 19770 15292 19782 15344
rect 19844 15292 19846 15344
rect 19684 15290 19708 15292
rect 19764 15290 19788 15292
rect 19844 15290 19868 15292
rect 19628 15270 19924 15290
rect 19628 14014 19924 14034
rect 19684 14012 19708 14014
rect 19764 14012 19788 14014
rect 19844 14012 19868 14014
rect 19706 13960 19708 14012
rect 19770 13960 19782 14012
rect 19844 13960 19846 14012
rect 19684 13958 19708 13960
rect 19764 13958 19788 13960
rect 19844 13958 19868 13960
rect 19628 13938 19924 13958
rect 19628 12682 19924 12702
rect 19684 12680 19708 12682
rect 19764 12680 19788 12682
rect 19844 12680 19868 12682
rect 19706 12628 19708 12680
rect 19770 12628 19782 12680
rect 19844 12628 19846 12680
rect 19684 12626 19708 12628
rect 19764 12626 19788 12628
rect 19844 12626 19868 12628
rect 19628 12606 19924 12626
rect 19628 11350 19924 11370
rect 19684 11348 19708 11350
rect 19764 11348 19788 11350
rect 19844 11348 19868 11350
rect 19706 11296 19708 11348
rect 19770 11296 19782 11348
rect 19844 11296 19846 11348
rect 19684 11294 19708 11296
rect 19764 11294 19788 11296
rect 19844 11294 19868 11296
rect 19628 11274 19924 11294
rect 19628 10018 19924 10038
rect 19684 10016 19708 10018
rect 19764 10016 19788 10018
rect 19844 10016 19868 10018
rect 19706 9964 19708 10016
rect 19770 9964 19782 10016
rect 19844 9964 19846 10016
rect 19684 9962 19708 9964
rect 19764 9962 19788 9964
rect 19844 9962 19868 9964
rect 19628 9942 19924 9962
rect 19318 9017 19370 9023
rect 19318 8959 19370 8965
rect 19628 8686 19924 8706
rect 19684 8684 19708 8686
rect 19764 8684 19788 8686
rect 19844 8684 19868 8686
rect 19706 8632 19708 8684
rect 19770 8632 19782 8684
rect 19844 8632 19846 8684
rect 19684 8630 19708 8632
rect 19764 8630 19788 8632
rect 19844 8630 19868 8632
rect 19628 8610 19924 8630
rect 19628 7354 19924 7374
rect 19684 7352 19708 7354
rect 19764 7352 19788 7354
rect 19844 7352 19868 7354
rect 19706 7300 19708 7352
rect 19770 7300 19782 7352
rect 19844 7300 19846 7352
rect 19684 7298 19708 7300
rect 19764 7298 19788 7300
rect 19844 7298 19868 7300
rect 19628 7278 19924 7298
rect 20002 6433 20030 55135
rect 20290 37439 20318 55505
rect 20278 37433 20330 37439
rect 20278 37375 20330 37381
rect 20386 31667 20414 56171
rect 21238 31735 21290 31741
rect 21238 31677 21290 31683
rect 20374 31661 20426 31667
rect 20374 31603 20426 31609
rect 21250 27374 21278 31677
rect 21334 28109 21386 28115
rect 21334 28051 21386 28057
rect 21346 27893 21374 28051
rect 21334 27887 21386 27893
rect 21334 27829 21386 27835
rect 21250 27346 21374 27374
rect 21238 18785 21290 18791
rect 21238 18727 21290 18733
rect 20374 9831 20426 9837
rect 20374 9773 20426 9779
rect 20386 7099 20414 9773
rect 20854 9757 20906 9763
rect 20854 9699 20906 9705
rect 20662 9461 20714 9467
rect 20662 9403 20714 9409
rect 20674 7173 20702 9403
rect 20758 7463 20810 7469
rect 20758 7405 20810 7411
rect 20662 7167 20714 7173
rect 20662 7109 20714 7115
rect 20374 7093 20426 7099
rect 20374 7035 20426 7041
rect 20374 6945 20426 6951
rect 20374 6887 20426 6893
rect 19126 6427 19178 6433
rect 19126 6369 19178 6375
rect 19990 6427 20042 6433
rect 19990 6369 20042 6375
rect 18934 6205 18986 6211
rect 18934 6147 18986 6153
rect 20086 6205 20138 6211
rect 20086 6147 20138 6153
rect 18838 3245 18890 3251
rect 18838 3187 18890 3193
rect 18838 3023 18890 3029
rect 18838 2965 18890 2971
rect 18850 800 18878 2965
rect 18946 800 18974 6147
rect 19318 6131 19370 6137
rect 19318 6073 19370 6079
rect 19030 5021 19082 5027
rect 19030 4963 19082 4969
rect 19126 5021 19178 5027
rect 19126 4963 19178 4969
rect 19042 3103 19070 4963
rect 19030 3097 19082 3103
rect 19030 3039 19082 3045
rect 19138 2012 19166 4963
rect 19222 3689 19274 3695
rect 19222 3631 19274 3637
rect 19042 1984 19166 2012
rect 19042 800 19070 1984
rect 19234 800 19262 3631
rect 19330 3029 19358 6073
rect 19628 6022 19924 6042
rect 19684 6020 19708 6022
rect 19764 6020 19788 6022
rect 19844 6020 19868 6022
rect 19706 5968 19708 6020
rect 19770 5968 19782 6020
rect 19844 5968 19846 6020
rect 19684 5966 19708 5968
rect 19764 5966 19788 5968
rect 19844 5966 19868 5968
rect 19628 5946 19924 5966
rect 19628 4690 19924 4710
rect 19684 4688 19708 4690
rect 19764 4688 19788 4690
rect 19844 4688 19868 4690
rect 19706 4636 19708 4688
rect 19770 4636 19782 4688
rect 19844 4636 19846 4688
rect 19684 4634 19708 4636
rect 19764 4634 19788 4636
rect 19844 4634 19868 4636
rect 19628 4614 19924 4634
rect 19414 3837 19466 3843
rect 19414 3779 19466 3785
rect 19318 3023 19370 3029
rect 19318 2965 19370 2971
rect 19426 2900 19454 3779
rect 19990 3689 20042 3695
rect 19990 3631 20042 3637
rect 19628 3358 19924 3378
rect 19684 3356 19708 3358
rect 19764 3356 19788 3358
rect 19844 3356 19868 3358
rect 19706 3304 19708 3356
rect 19770 3304 19782 3356
rect 19844 3304 19846 3356
rect 19684 3302 19708 3304
rect 19764 3302 19788 3304
rect 19844 3302 19868 3304
rect 19628 3282 19924 3302
rect 19702 3245 19754 3251
rect 19702 3187 19754 3193
rect 19606 3023 19658 3029
rect 19606 2965 19658 2971
rect 19330 2872 19454 2900
rect 19330 800 19358 2872
rect 19414 2505 19466 2511
rect 19414 2447 19466 2453
rect 19426 800 19454 2447
rect 19618 800 19646 2965
rect 19714 800 19742 3187
rect 19894 3171 19946 3177
rect 19894 3113 19946 3119
rect 19798 2949 19850 2955
rect 19798 2891 19850 2897
rect 19810 800 19838 2891
rect 19906 2511 19934 3113
rect 19894 2505 19946 2511
rect 19894 2447 19946 2453
rect 20002 1864 20030 3631
rect 19906 1836 20030 1864
rect 19906 800 19934 1836
rect 20098 800 20126 6147
rect 20182 5687 20234 5693
rect 20182 5629 20234 5635
rect 20194 2955 20222 5629
rect 20278 4355 20330 4361
rect 20278 4297 20330 4303
rect 20182 2949 20234 2955
rect 20182 2891 20234 2897
rect 20182 1839 20234 1845
rect 20182 1781 20234 1787
rect 20194 800 20222 1781
rect 20290 800 20318 4297
rect 20386 3251 20414 6887
rect 20662 6131 20714 6137
rect 20662 6073 20714 6079
rect 20566 5687 20618 5693
rect 20566 5629 20618 5635
rect 20470 5021 20522 5027
rect 20470 4963 20522 4969
rect 20374 3245 20426 3251
rect 20374 3187 20426 3193
rect 20482 3177 20510 4963
rect 20470 3171 20522 3177
rect 20470 3113 20522 3119
rect 20470 2875 20522 2881
rect 20470 2817 20522 2823
rect 20482 800 20510 2817
rect 20578 800 20606 5629
rect 20674 3843 20702 6073
rect 20662 3837 20714 3843
rect 20662 3779 20714 3785
rect 20662 3689 20714 3695
rect 20662 3631 20714 3637
rect 20674 800 20702 3631
rect 20770 800 20798 7405
rect 20866 6433 20894 9699
rect 20950 8795 21002 8801
rect 20950 8737 21002 8743
rect 20962 7765 20990 8737
rect 20950 7759 21002 7765
rect 20950 7701 21002 7707
rect 21250 7617 21278 18727
rect 21346 11095 21374 27346
rect 21442 15609 21470 56171
rect 21430 15603 21482 15609
rect 21430 15545 21482 15551
rect 22210 15239 22238 56171
rect 22678 52751 22730 52757
rect 22678 52693 22730 52699
rect 22294 34917 22346 34923
rect 22294 34859 22346 34865
rect 22198 15233 22250 15239
rect 22198 15175 22250 15181
rect 21334 11089 21386 11095
rect 21334 11031 21386 11037
rect 21526 9905 21578 9911
rect 21526 9847 21578 9853
rect 21238 7611 21290 7617
rect 21238 7553 21290 7559
rect 21430 7093 21482 7099
rect 21430 7035 21482 7041
rect 20950 6945 21002 6951
rect 21238 6945 21290 6951
rect 20950 6887 21002 6893
rect 21154 6905 21238 6933
rect 20854 6427 20906 6433
rect 20854 6369 20906 6375
rect 20962 3011 20990 6887
rect 21046 4355 21098 4361
rect 21046 4297 21098 4303
rect 20866 2983 20990 3011
rect 20866 2955 20894 2983
rect 20854 2949 20906 2955
rect 20854 2891 20906 2897
rect 20950 2949 21002 2955
rect 20950 2891 21002 2897
rect 20962 800 20990 2891
rect 21058 800 21086 4297
rect 21154 800 21182 6905
rect 21238 6887 21290 6893
rect 21238 5021 21290 5027
rect 21238 4963 21290 4969
rect 21250 1845 21278 4963
rect 21334 3911 21386 3917
rect 21334 3853 21386 3859
rect 21238 1839 21290 1845
rect 21238 1781 21290 1787
rect 21346 1716 21374 3853
rect 21442 3177 21470 7035
rect 21538 6433 21566 9847
rect 21718 9831 21770 9837
rect 21718 9773 21770 9779
rect 21730 9097 21758 9773
rect 21718 9091 21770 9097
rect 21718 9033 21770 9039
rect 22306 8801 22334 34859
rect 22294 8795 22346 8801
rect 22294 8737 22346 8743
rect 22690 7099 22718 52693
rect 22978 35589 23006 56171
rect 23362 55717 23390 59200
rect 23842 56975 23870 59200
rect 23830 56969 23882 56975
rect 23830 56911 23882 56917
rect 24022 56895 24074 56901
rect 24022 56837 24074 56843
rect 23350 55711 23402 55717
rect 23350 55653 23402 55659
rect 23158 55563 23210 55569
rect 23158 55505 23210 55511
rect 23170 55421 23198 55505
rect 23158 55415 23210 55421
rect 23158 55357 23210 55363
rect 22966 35583 23018 35589
rect 22966 35525 23018 35531
rect 22966 34251 23018 34257
rect 22966 34193 23018 34199
rect 22978 7543 23006 34193
rect 23170 8875 23198 55357
rect 23830 50531 23882 50537
rect 23830 50473 23882 50479
rect 23734 17453 23786 17459
rect 23734 17395 23786 17401
rect 23158 8869 23210 8875
rect 23158 8811 23210 8817
rect 22966 7537 23018 7543
rect 22966 7479 23018 7485
rect 22678 7093 22730 7099
rect 22678 7035 22730 7041
rect 22006 6945 22058 6951
rect 21922 6905 22006 6933
rect 21526 6427 21578 6433
rect 21526 6369 21578 6375
rect 21526 6131 21578 6137
rect 21526 6073 21578 6079
rect 21430 3171 21482 3177
rect 21430 3113 21482 3119
rect 21430 3023 21482 3029
rect 21430 2965 21482 2971
rect 21250 1688 21374 1716
rect 21250 800 21278 1688
rect 21442 800 21470 2965
rect 21538 800 21566 6073
rect 21814 5687 21866 5693
rect 21634 5647 21814 5675
rect 21634 800 21662 5647
rect 21814 5629 21866 5635
rect 21718 5539 21770 5545
rect 21718 5481 21770 5487
rect 21730 2955 21758 5481
rect 21814 4355 21866 4361
rect 21814 4297 21866 4303
rect 21718 2949 21770 2955
rect 21718 2891 21770 2897
rect 21826 800 21854 4297
rect 21922 800 21950 6905
rect 22006 6887 22058 6893
rect 23350 6945 23402 6951
rect 23350 6887 23402 6893
rect 22294 6205 22346 6211
rect 22294 6147 22346 6153
rect 22006 4281 22058 4287
rect 22006 4223 22058 4229
rect 22018 800 22046 4223
rect 22102 3689 22154 3695
rect 22102 3631 22154 3637
rect 22114 800 22142 3631
rect 22306 800 22334 6147
rect 23062 5687 23114 5693
rect 23062 5629 23114 5635
rect 22774 5021 22826 5027
rect 22774 4963 22826 4969
rect 22786 3917 22814 4963
rect 22774 3911 22826 3917
rect 22774 3853 22826 3859
rect 23074 3788 23102 5629
rect 23158 4947 23210 4953
rect 23158 4889 23210 4895
rect 22786 3760 23102 3788
rect 22582 3541 22634 3547
rect 22582 3483 22634 3489
rect 22390 3097 22442 3103
rect 22390 3039 22442 3045
rect 22402 800 22430 3039
rect 22486 2949 22538 2955
rect 22486 2891 22538 2897
rect 22498 800 22526 2891
rect 22594 800 22622 3483
rect 22786 800 22814 3760
rect 22870 3689 22922 3695
rect 22870 3631 22922 3637
rect 22882 800 22910 3631
rect 22966 3467 23018 3473
rect 22966 3409 23018 3415
rect 22978 800 23006 3409
rect 23170 800 23198 4889
rect 23254 4355 23306 4361
rect 23254 4297 23306 4303
rect 23266 800 23294 4297
rect 23362 3547 23390 6887
rect 23746 6433 23774 17395
rect 23842 12224 23870 50473
rect 23926 39431 23978 39437
rect 23926 39373 23978 39379
rect 23938 12372 23966 39373
rect 24034 12668 24062 56837
rect 24418 56531 24446 59200
rect 24406 56525 24458 56531
rect 24406 56467 24458 56473
rect 24898 55717 24926 59200
rect 25474 56975 25502 59200
rect 25462 56969 25514 56975
rect 25462 56911 25514 56917
rect 25954 56531 25982 59200
rect 26530 56531 26558 59200
rect 27010 56975 27038 59200
rect 26998 56969 27050 56975
rect 26998 56911 27050 56917
rect 27190 56895 27242 56901
rect 27190 56837 27242 56843
rect 25942 56525 25994 56531
rect 25942 56467 25994 56473
rect 26518 56525 26570 56531
rect 26518 56467 26570 56473
rect 26614 56451 26666 56457
rect 26614 56393 26666 56399
rect 26134 56229 26186 56235
rect 26134 56171 26186 56177
rect 24886 55711 24938 55717
rect 24886 55653 24938 55659
rect 24886 55563 24938 55569
rect 24886 55505 24938 55511
rect 25654 55563 25706 55569
rect 25654 55505 25706 55511
rect 24898 55421 24926 55505
rect 25666 55421 25694 55505
rect 24886 55415 24938 55421
rect 24886 55357 24938 55363
rect 25654 55415 25706 55421
rect 25654 55357 25706 55363
rect 24118 38765 24170 38771
rect 24118 38707 24170 38713
rect 24130 17294 24158 38707
rect 24130 17266 24350 17294
rect 24034 12640 24254 12668
rect 23938 12344 24062 12372
rect 23842 12196 23966 12224
rect 23830 7463 23882 7469
rect 23830 7405 23882 7411
rect 23734 6427 23786 6433
rect 23734 6369 23786 6375
rect 23446 5687 23498 5693
rect 23446 5629 23498 5635
rect 23350 3541 23402 3547
rect 23350 3483 23402 3489
rect 23350 3245 23402 3251
rect 23350 3187 23402 3193
rect 23362 800 23390 3187
rect 23458 800 23486 5629
rect 23542 5021 23594 5027
rect 23542 4963 23594 4969
rect 23554 3103 23582 4963
rect 23638 3689 23690 3695
rect 23842 3640 23870 7405
rect 23938 7173 23966 12196
rect 24034 7765 24062 12344
rect 24226 11021 24254 12640
rect 24322 11761 24350 17266
rect 24310 11755 24362 11761
rect 24310 11697 24362 11703
rect 24214 11015 24266 11021
rect 24214 10957 24266 10963
rect 24502 11015 24554 11021
rect 24502 10957 24554 10963
rect 24022 7759 24074 7765
rect 24022 7701 24074 7707
rect 24118 7463 24170 7469
rect 24118 7405 24170 7411
rect 23926 7167 23978 7173
rect 23926 7109 23978 7115
rect 23926 6945 23978 6951
rect 23926 6887 23978 6893
rect 23638 3631 23690 3637
rect 23542 3097 23594 3103
rect 23542 3039 23594 3045
rect 23650 800 23678 3631
rect 23746 3612 23870 3640
rect 23746 800 23774 3612
rect 23938 3251 23966 6887
rect 24022 6131 24074 6137
rect 24022 6073 24074 6079
rect 24034 3473 24062 6073
rect 24022 3467 24074 3473
rect 24022 3409 24074 3415
rect 23926 3245 23978 3251
rect 23926 3187 23978 3193
rect 23830 3171 23882 3177
rect 23830 3113 23882 3119
rect 23842 800 23870 3113
rect 24022 3023 24074 3029
rect 24022 2965 24074 2971
rect 24034 800 24062 2965
rect 24130 800 24158 7405
rect 24514 6433 24542 10957
rect 24790 7463 24842 7469
rect 24790 7405 24842 7411
rect 24598 6945 24650 6951
rect 24598 6887 24650 6893
rect 24502 6427 24554 6433
rect 24502 6369 24554 6375
rect 24610 5860 24638 6887
rect 24514 5832 24638 5860
rect 24214 3837 24266 3843
rect 24214 3779 24266 3785
rect 24226 800 24254 3779
rect 24406 3689 24458 3695
rect 24406 3631 24458 3637
rect 24418 1864 24446 3631
rect 24322 1836 24446 1864
rect 24322 800 24350 1836
rect 24514 800 24542 5832
rect 24598 5687 24650 5693
rect 24598 5629 24650 5635
rect 24610 800 24638 5629
rect 24694 3615 24746 3621
rect 24694 3557 24746 3563
rect 24706 800 24734 3557
rect 24802 800 24830 7405
rect 24898 3103 24926 55357
rect 25462 23891 25514 23897
rect 25462 23833 25514 23839
rect 25174 10349 25226 10355
rect 25174 10291 25226 10297
rect 25186 7025 25214 10291
rect 25474 7765 25502 23833
rect 25666 13759 25694 55357
rect 26146 44173 26174 56171
rect 26134 44167 26186 44173
rect 26134 44109 26186 44115
rect 25750 41429 25802 41435
rect 25750 41371 25802 41377
rect 25762 41213 25790 41371
rect 25750 41207 25802 41213
rect 25750 41149 25802 41155
rect 26230 27591 26282 27597
rect 26230 27533 26282 27539
rect 25750 22559 25802 22565
rect 25750 22501 25802 22507
rect 25654 13753 25706 13759
rect 25654 13695 25706 13701
rect 25462 7759 25514 7765
rect 25462 7701 25514 7707
rect 25558 7463 25610 7469
rect 25558 7405 25610 7411
rect 25174 7019 25226 7025
rect 25174 6961 25226 6967
rect 25174 6871 25226 6877
rect 25174 6813 25226 6819
rect 25078 5021 25130 5027
rect 25078 4963 25130 4969
rect 24982 3245 25034 3251
rect 24982 3187 25034 3193
rect 24886 3097 24938 3103
rect 24886 3039 24938 3045
rect 24994 800 25022 3187
rect 25090 3177 25118 4963
rect 25078 3171 25130 3177
rect 25078 3113 25130 3119
rect 25078 2949 25130 2955
rect 25078 2891 25130 2897
rect 25090 800 25118 2891
rect 25186 800 25214 6813
rect 25462 4355 25514 4361
rect 25462 4297 25514 4303
rect 25366 3097 25418 3103
rect 25366 3039 25418 3045
rect 25378 800 25406 3039
rect 25474 800 25502 4297
rect 25570 800 25598 7405
rect 25762 7099 25790 22501
rect 25846 9461 25898 9467
rect 25846 9403 25898 9409
rect 25858 7247 25886 9403
rect 26242 7765 26270 27533
rect 26422 26777 26474 26783
rect 26422 26719 26474 26725
rect 26230 7759 26282 7765
rect 26230 7701 26282 7707
rect 25846 7241 25898 7247
rect 25846 7183 25898 7189
rect 26434 7099 26462 26719
rect 26626 22861 26654 56393
rect 26806 56229 26858 56235
rect 26806 56171 26858 56177
rect 26614 22855 26666 22861
rect 26614 22797 26666 22803
rect 26818 10873 26846 56171
rect 26902 24927 26954 24933
rect 26902 24869 26954 24875
rect 26806 10867 26858 10873
rect 26806 10809 26858 10815
rect 26614 10275 26666 10281
rect 26614 10217 26666 10223
rect 25750 7093 25802 7099
rect 25750 7035 25802 7041
rect 26422 7093 26474 7099
rect 26422 7035 26474 7041
rect 25942 7019 25994 7025
rect 25942 6961 25994 6967
rect 25654 6353 25706 6359
rect 25654 6295 25706 6301
rect 25666 800 25694 6295
rect 25846 5021 25898 5027
rect 25846 4963 25898 4969
rect 25858 3843 25886 4963
rect 25846 3837 25898 3843
rect 25846 3779 25898 3785
rect 25846 3541 25898 3547
rect 25846 3483 25898 3489
rect 25858 800 25886 3483
rect 25954 800 25982 6961
rect 26626 6803 26654 10217
rect 26806 9165 26858 9171
rect 26806 9107 26858 9113
rect 26710 7463 26762 7469
rect 26710 7405 26762 7411
rect 26614 6797 26666 6803
rect 26614 6739 26666 6745
rect 26326 6131 26378 6137
rect 26326 6073 26378 6079
rect 26230 5687 26282 5693
rect 26230 5629 26282 5635
rect 26038 5539 26090 5545
rect 26038 5481 26090 5487
rect 26050 800 26078 5481
rect 26134 4355 26186 4361
rect 26134 4297 26186 4303
rect 26146 800 26174 4297
rect 26242 3103 26270 5629
rect 26230 3097 26282 3103
rect 26230 3039 26282 3045
rect 26338 800 26366 6073
rect 26614 5021 26666 5027
rect 26614 4963 26666 4969
rect 26518 4355 26570 4361
rect 26518 4297 26570 4303
rect 26422 3837 26474 3843
rect 26422 3779 26474 3785
rect 26434 800 26462 3779
rect 26530 800 26558 4297
rect 26626 3251 26654 4963
rect 26614 3245 26666 3251
rect 26614 3187 26666 3193
rect 26722 800 26750 7405
rect 26818 7173 26846 9107
rect 26914 8875 26942 24869
rect 27202 12353 27230 56837
rect 27586 56531 27614 59200
rect 28066 56531 28094 59200
rect 28642 56975 28670 59200
rect 29122 57049 29150 59200
rect 29110 57043 29162 57049
rect 29110 56985 29162 56991
rect 28630 56969 28682 56975
rect 28630 56911 28682 56917
rect 29698 56531 29726 59200
rect 30178 56957 30206 59200
rect 30262 56969 30314 56975
rect 30178 56929 30262 56957
rect 30262 56911 30314 56917
rect 29974 56895 30026 56901
rect 29974 56837 30026 56843
rect 27574 56525 27626 56531
rect 27574 56467 27626 56473
rect 28054 56525 28106 56531
rect 28054 56467 28106 56473
rect 29686 56525 29738 56531
rect 29686 56467 29738 56473
rect 28726 56377 28778 56383
rect 28726 56319 28778 56325
rect 27478 56229 27530 56235
rect 27478 56171 27530 56177
rect 28150 56229 28202 56235
rect 28150 56171 28202 56177
rect 27490 13907 27518 56171
rect 28162 17294 28190 56171
rect 28738 47873 28766 56319
rect 29302 56229 29354 56235
rect 29302 56171 29354 56177
rect 28726 47867 28778 47873
rect 28726 47809 28778 47815
rect 29110 40837 29162 40843
rect 29110 40779 29162 40785
rect 28534 34769 28586 34775
rect 28534 34711 28586 34717
rect 28546 17294 28574 34711
rect 29014 28109 29066 28115
rect 29014 28051 29066 28057
rect 27970 17266 28190 17294
rect 28258 17266 28574 17294
rect 27478 13901 27530 13907
rect 27478 13843 27530 13849
rect 27190 12347 27242 12353
rect 27190 12289 27242 12295
rect 26902 8869 26954 8875
rect 26902 8811 26954 8817
rect 26998 8795 27050 8801
rect 26998 8737 27050 8743
rect 27010 7765 27038 8737
rect 26998 7759 27050 7765
rect 26998 7701 27050 7707
rect 26806 7167 26858 7173
rect 26806 7109 26858 7115
rect 26998 6871 27050 6877
rect 26998 6813 27050 6819
rect 27766 6871 27818 6877
rect 27766 6813 27818 6819
rect 26806 6353 26858 6359
rect 26806 6295 26858 6301
rect 26818 800 26846 6295
rect 26902 3023 26954 3029
rect 26902 2965 26954 2971
rect 26914 800 26942 2965
rect 27010 800 27038 6813
rect 27382 5687 27434 5693
rect 27382 5629 27434 5635
rect 27394 3788 27422 5629
rect 27478 4207 27530 4213
rect 27478 4149 27530 4155
rect 27202 3760 27422 3788
rect 27202 800 27230 3760
rect 27286 3689 27338 3695
rect 27286 3631 27338 3637
rect 27298 800 27326 3631
rect 27490 3196 27518 4149
rect 27394 3168 27518 3196
rect 27394 800 27422 3168
rect 27478 3097 27530 3103
rect 27478 3039 27530 3045
rect 27490 800 27518 3039
rect 27670 2949 27722 2955
rect 27670 2891 27722 2897
rect 27682 800 27710 2891
rect 27778 800 27806 6813
rect 27862 5687 27914 5693
rect 27862 5629 27914 5635
rect 27874 800 27902 5629
rect 27970 2881 27998 17266
rect 28150 13013 28202 13019
rect 28150 12955 28202 12961
rect 28162 9412 28190 12955
rect 28258 9615 28286 17266
rect 28438 10867 28490 10873
rect 28438 10809 28490 10815
rect 28246 9609 28298 9615
rect 28246 9551 28298 9557
rect 28342 9609 28394 9615
rect 28342 9551 28394 9557
rect 28162 9384 28286 9412
rect 28150 7463 28202 7469
rect 28150 7405 28202 7411
rect 28054 5021 28106 5027
rect 28054 4963 28106 4969
rect 28066 3843 28094 4963
rect 28054 3837 28106 3843
rect 28054 3779 28106 3785
rect 28054 3541 28106 3547
rect 28054 3483 28106 3489
rect 27958 2875 28010 2881
rect 27958 2817 28010 2823
rect 28066 800 28094 3483
rect 28162 800 28190 7405
rect 28258 6433 28286 9384
rect 28354 7099 28382 9551
rect 28450 7765 28478 10809
rect 28726 9165 28778 9171
rect 28726 9107 28778 9113
rect 28438 7759 28490 7765
rect 28438 7701 28490 7707
rect 28738 7099 28766 9107
rect 28342 7093 28394 7099
rect 28342 7035 28394 7041
rect 28726 7093 28778 7099
rect 28726 7035 28778 7041
rect 29026 6433 29054 28051
rect 29122 7173 29150 40779
rect 29314 12575 29342 56171
rect 29590 37433 29642 37439
rect 29590 37375 29642 37381
rect 29494 32993 29546 32999
rect 29494 32935 29546 32941
rect 29398 23521 29450 23527
rect 29398 23463 29450 23469
rect 29302 12569 29354 12575
rect 29302 12511 29354 12517
rect 29410 7765 29438 23463
rect 29506 9615 29534 32935
rect 29602 10873 29630 37375
rect 29986 13537 30014 56837
rect 30658 56531 30686 59200
rect 31234 56531 31262 59200
rect 31714 56975 31742 59200
rect 31702 56969 31754 56975
rect 31702 56911 31754 56917
rect 32290 56531 32318 59200
rect 30646 56525 30698 56531
rect 30646 56467 30698 56473
rect 31222 56525 31274 56531
rect 31222 56467 31274 56473
rect 32278 56525 32330 56531
rect 32278 56467 32330 56473
rect 30934 56229 30986 56235
rect 30934 56171 30986 56177
rect 31702 56229 31754 56235
rect 31702 56171 31754 56177
rect 32470 56229 32522 56235
rect 32470 56171 32522 56177
rect 30070 54749 30122 54755
rect 30070 54691 30122 54697
rect 29974 13531 30026 13537
rect 29974 13473 30026 13479
rect 29590 10867 29642 10873
rect 29590 10809 29642 10815
rect 29494 9609 29546 9615
rect 29494 9551 29546 9557
rect 29398 7759 29450 7765
rect 29398 7701 29450 7707
rect 29590 7759 29642 7765
rect 29590 7701 29642 7707
rect 29206 7463 29258 7469
rect 29206 7405 29258 7411
rect 29110 7167 29162 7173
rect 29110 7109 29162 7115
rect 28246 6427 28298 6433
rect 28246 6369 28298 6375
rect 29014 6427 29066 6433
rect 29014 6369 29066 6375
rect 29014 6131 29066 6137
rect 29014 6073 29066 6079
rect 28822 5687 28874 5693
rect 28822 5629 28874 5635
rect 28342 4355 28394 4361
rect 28342 4297 28394 4303
rect 28246 3171 28298 3177
rect 28246 3113 28298 3119
rect 28258 800 28286 3113
rect 28354 800 28382 4297
rect 28534 3911 28586 3917
rect 28534 3853 28586 3859
rect 28546 800 28574 3853
rect 28834 3640 28862 5629
rect 28918 5021 28970 5027
rect 28918 4963 28970 4969
rect 28642 3612 28862 3640
rect 28642 800 28670 3612
rect 28726 3467 28778 3473
rect 28726 3409 28778 3415
rect 28738 800 28766 3409
rect 28822 3245 28874 3251
rect 28822 3187 28874 3193
rect 28834 2937 28862 3187
rect 28930 3103 28958 4963
rect 29026 4213 29054 6073
rect 29110 4355 29162 4361
rect 29110 4297 29162 4303
rect 29014 4207 29066 4213
rect 29014 4149 29066 4155
rect 29014 3837 29066 3843
rect 29014 3779 29066 3785
rect 28918 3097 28970 3103
rect 28918 3039 28970 3045
rect 28834 2909 28958 2937
rect 28930 800 28958 2909
rect 29026 800 29054 3779
rect 29122 800 29150 4297
rect 29218 800 29246 7405
rect 29494 6945 29546 6951
rect 29494 6887 29546 6893
rect 29302 5021 29354 5027
rect 29302 4963 29354 4969
rect 29314 3177 29342 4963
rect 29506 3917 29534 6887
rect 29494 3911 29546 3917
rect 29494 3853 29546 3859
rect 29302 3171 29354 3177
rect 29302 3113 29354 3119
rect 29494 3171 29546 3177
rect 29494 3113 29546 3119
rect 29398 3097 29450 3103
rect 29398 3039 29450 3045
rect 29410 800 29438 3039
rect 29506 800 29534 3113
rect 29602 800 29630 7701
rect 30082 7691 30110 54691
rect 30946 52831 30974 56171
rect 30934 52825 30986 52831
rect 30934 52767 30986 52773
rect 31318 50753 31370 50759
rect 31318 50695 31370 50701
rect 31510 50753 31562 50759
rect 31510 50695 31562 50701
rect 31330 50463 31358 50695
rect 31522 50537 31550 50695
rect 31510 50531 31562 50537
rect 31510 50473 31562 50479
rect 31318 50457 31370 50463
rect 31318 50399 31370 50405
rect 30934 49125 30986 49131
rect 30934 49067 30986 49073
rect 30262 37211 30314 37217
rect 30262 37153 30314 37159
rect 30166 16565 30218 16571
rect 30166 16507 30218 16513
rect 30178 8801 30206 16507
rect 30166 8795 30218 8801
rect 30166 8737 30218 8743
rect 30070 7685 30122 7691
rect 30070 7627 30122 7633
rect 29974 6945 30026 6951
rect 29974 6887 30026 6893
rect 29686 6353 29738 6359
rect 29686 6295 29738 6301
rect 29698 800 29726 6295
rect 29782 6131 29834 6137
rect 29782 6073 29834 6079
rect 29794 3251 29822 6073
rect 29878 3689 29930 3695
rect 29878 3631 29930 3637
rect 29782 3245 29834 3251
rect 29782 3187 29834 3193
rect 29890 3177 29918 3631
rect 29878 3171 29930 3177
rect 29878 3113 29930 3119
rect 29878 3023 29930 3029
rect 29878 2965 29930 2971
rect 29890 800 29918 2965
rect 29986 800 30014 6887
rect 30274 6581 30302 37153
rect 30946 7099 30974 49067
rect 31714 27227 31742 56171
rect 32374 51197 32426 51203
rect 32374 51139 32426 51145
rect 31798 50161 31850 50167
rect 31798 50103 31850 50109
rect 31702 27221 31754 27227
rect 31702 27163 31754 27169
rect 31702 24927 31754 24933
rect 31702 24869 31754 24875
rect 31222 8129 31274 8135
rect 31222 8071 31274 8077
rect 31234 7765 31262 8071
rect 31222 7759 31274 7765
rect 31222 7701 31274 7707
rect 31030 7463 31082 7469
rect 31030 7405 31082 7411
rect 30934 7093 30986 7099
rect 30934 7035 30986 7041
rect 30742 6871 30794 6877
rect 30742 6813 30794 6819
rect 30262 6575 30314 6581
rect 30262 6517 30314 6523
rect 30646 6427 30698 6433
rect 30646 6369 30698 6375
rect 30262 5687 30314 5693
rect 30262 5629 30314 5635
rect 30274 2900 30302 5629
rect 30358 5021 30410 5027
rect 30358 4963 30410 4969
rect 30370 3843 30398 4963
rect 30358 3837 30410 3843
rect 30358 3779 30410 3785
rect 30454 3689 30506 3695
rect 30082 2872 30302 2900
rect 30370 3649 30454 3677
rect 30082 800 30110 2872
rect 30370 1864 30398 3649
rect 30454 3631 30506 3637
rect 30454 3245 30506 3251
rect 30454 3187 30506 3193
rect 30274 1836 30398 1864
rect 30274 800 30302 1836
rect 30358 1765 30410 1771
rect 30358 1707 30410 1713
rect 30370 800 30398 1707
rect 30466 800 30494 3187
rect 30550 2949 30602 2955
rect 30550 2891 30602 2897
rect 30562 800 30590 2891
rect 30658 1771 30686 6369
rect 30646 1765 30698 1771
rect 30646 1707 30698 1713
rect 30754 800 30782 6813
rect 30838 5687 30890 5693
rect 30838 5629 30890 5635
rect 30850 800 30878 5629
rect 30934 4355 30986 4361
rect 30934 4297 30986 4303
rect 30946 800 30974 4297
rect 31042 800 31070 7405
rect 31714 7099 31742 24869
rect 31702 7093 31754 7099
rect 31702 7035 31754 7041
rect 31414 7019 31466 7025
rect 31414 6961 31466 6967
rect 31222 6353 31274 6359
rect 31222 6295 31274 6301
rect 31126 5021 31178 5027
rect 31126 4963 31178 4969
rect 31138 3103 31166 4963
rect 31126 3097 31178 3103
rect 31126 3039 31178 3045
rect 31234 800 31262 6295
rect 31318 3689 31370 3695
rect 31318 3631 31370 3637
rect 31330 800 31358 3631
rect 31426 800 31454 6961
rect 31810 6581 31838 50103
rect 32182 32105 32234 32111
rect 32182 32047 32234 32053
rect 32194 31889 32222 32047
rect 32182 31883 32234 31889
rect 32182 31825 32234 31831
rect 31990 24113 32042 24119
rect 31990 24055 32042 24061
rect 32002 23897 32030 24055
rect 31990 23891 32042 23897
rect 31990 23833 32042 23839
rect 32386 7099 32414 51139
rect 32482 35071 32510 56171
rect 32770 56161 32798 59200
rect 33346 56975 33374 59200
rect 33334 56969 33386 56975
rect 33334 56911 33386 56917
rect 33826 56531 33854 59200
rect 34402 57614 34430 59200
rect 34402 57586 34622 57614
rect 34102 56895 34154 56901
rect 34102 56837 34154 56843
rect 33814 56525 33866 56531
rect 33814 56467 33866 56473
rect 32854 56229 32906 56235
rect 32854 56171 32906 56177
rect 34006 56229 34058 56235
rect 34006 56171 34058 56177
rect 32758 56155 32810 56161
rect 32758 56097 32810 56103
rect 32470 35065 32522 35071
rect 32470 35007 32522 35013
rect 32566 20117 32618 20123
rect 32566 20059 32618 20065
rect 32374 7093 32426 7099
rect 32374 7035 32426 7041
rect 32578 7025 32606 20059
rect 32866 13685 32894 56171
rect 33814 46313 33866 46319
rect 33814 46255 33866 46261
rect 32950 40097 33002 40103
rect 32950 40039 33002 40045
rect 32854 13679 32906 13685
rect 32854 13621 32906 13627
rect 32962 9245 32990 40039
rect 33238 32771 33290 32777
rect 33238 32713 33290 32719
rect 33046 21449 33098 21455
rect 33046 21391 33098 21397
rect 33058 9245 33086 21391
rect 32950 9239 33002 9245
rect 32950 9181 33002 9187
rect 33046 9239 33098 9245
rect 33046 9181 33098 9187
rect 33250 7099 33278 32713
rect 33526 12125 33578 12131
rect 33526 12067 33578 12073
rect 33238 7093 33290 7099
rect 33238 7035 33290 7041
rect 32566 7019 32618 7025
rect 32566 6961 32618 6967
rect 32182 6871 32234 6877
rect 32182 6813 32234 6819
rect 31798 6575 31850 6581
rect 31798 6517 31850 6523
rect 31798 6205 31850 6211
rect 31798 6147 31850 6153
rect 31702 5687 31754 5693
rect 31702 5629 31754 5635
rect 31714 4528 31742 5629
rect 31618 4500 31742 4528
rect 31618 800 31646 4500
rect 31702 4355 31754 4361
rect 31702 4297 31754 4303
rect 31714 800 31742 4297
rect 31810 800 31838 6147
rect 31894 5021 31946 5027
rect 31894 4963 31946 4969
rect 31906 3251 31934 4963
rect 31894 3245 31946 3251
rect 31894 3187 31946 3193
rect 31894 3097 31946 3103
rect 31894 3039 31946 3045
rect 31906 800 31934 3039
rect 32086 3023 32138 3029
rect 32086 2965 32138 2971
rect 32098 800 32126 2965
rect 32194 800 32222 6813
rect 32950 6797 33002 6803
rect 32950 6739 33002 6745
rect 32758 4355 32810 4361
rect 32758 4297 32810 4303
rect 32566 3911 32618 3917
rect 32566 3853 32618 3859
rect 32470 3689 32522 3695
rect 32470 3631 32522 3637
rect 32278 2949 32330 2955
rect 32278 2891 32330 2897
rect 32290 800 32318 2891
rect 32482 800 32510 3631
rect 32578 800 32606 3853
rect 32662 3245 32714 3251
rect 32662 3187 32714 3193
rect 32674 800 32702 3187
rect 32770 800 32798 4297
rect 32962 800 32990 6739
rect 33538 6433 33566 12067
rect 33826 11021 33854 46255
rect 34018 13093 34046 56171
rect 34114 14203 34142 56837
rect 34594 56531 34622 57586
rect 34882 56975 34910 59200
rect 34988 57304 35284 57324
rect 35044 57302 35068 57304
rect 35124 57302 35148 57304
rect 35204 57302 35228 57304
rect 35066 57250 35068 57302
rect 35130 57250 35142 57302
rect 35204 57250 35206 57302
rect 35044 57248 35068 57250
rect 35124 57248 35148 57250
rect 35204 57248 35228 57250
rect 34988 57228 35284 57248
rect 34870 56969 34922 56975
rect 34870 56911 34922 56917
rect 34582 56525 34634 56531
rect 34582 56467 34634 56473
rect 34390 56229 34442 56235
rect 34390 56171 34442 56177
rect 34198 47645 34250 47651
rect 34198 47587 34250 47593
rect 34102 14197 34154 14203
rect 34102 14139 34154 14145
rect 34006 13087 34058 13093
rect 34006 13029 34058 13035
rect 33814 11015 33866 11021
rect 33814 10957 33866 10963
rect 33910 7611 33962 7617
rect 33910 7553 33962 7559
rect 33622 7463 33674 7469
rect 33622 7405 33674 7411
rect 33526 6427 33578 6433
rect 33526 6369 33578 6375
rect 33142 5687 33194 5693
rect 33142 5629 33194 5635
rect 33238 5687 33290 5693
rect 33238 5629 33290 5635
rect 33046 3467 33098 3473
rect 33046 3409 33098 3415
rect 33058 2881 33086 3409
rect 33154 2955 33182 5629
rect 33142 2949 33194 2955
rect 33142 2891 33194 2897
rect 33046 2875 33098 2881
rect 33046 2817 33098 2823
rect 33250 2752 33278 5629
rect 33334 5021 33386 5027
rect 33334 4963 33386 4969
rect 33346 3103 33374 4963
rect 33430 3837 33482 3843
rect 33430 3779 33482 3785
rect 33334 3097 33386 3103
rect 33334 3039 33386 3045
rect 33334 2949 33386 2955
rect 33334 2891 33386 2897
rect 33058 2724 33278 2752
rect 33058 800 33086 2724
rect 33346 1420 33374 2891
rect 33154 1392 33374 1420
rect 33154 800 33182 1392
rect 33238 1321 33290 1327
rect 33238 1263 33290 1269
rect 33250 800 33278 1263
rect 33442 800 33470 3779
rect 33526 3689 33578 3695
rect 33526 3631 33578 3637
rect 33538 800 33566 3631
rect 33634 800 33662 7405
rect 33814 7093 33866 7099
rect 33814 7035 33866 7041
rect 33718 6205 33770 6211
rect 33718 6147 33770 6153
rect 33730 1327 33758 6147
rect 33826 3473 33854 7035
rect 33922 4509 33950 7553
rect 34006 6871 34058 6877
rect 34006 6813 34058 6819
rect 33910 4503 33962 4509
rect 33910 4445 33962 4451
rect 33910 4355 33962 4361
rect 33910 4297 33962 4303
rect 33814 3467 33866 3473
rect 33814 3409 33866 3415
rect 33814 3171 33866 3177
rect 33814 3113 33866 3119
rect 33718 1321 33770 1327
rect 33718 1263 33770 1269
rect 33826 800 33854 3113
rect 33922 800 33950 4297
rect 34018 800 34046 6813
rect 34210 6433 34238 47587
rect 34402 23675 34430 56171
rect 35458 56161 35486 59200
rect 35938 56513 35966 59200
rect 36514 56901 36542 59200
rect 36994 57614 37022 59200
rect 36994 57586 37118 57614
rect 36502 56895 36554 56901
rect 36502 56837 36554 56843
rect 36694 56747 36746 56753
rect 36694 56689 36746 56695
rect 36022 56525 36074 56531
rect 35938 56485 36022 56513
rect 36022 56467 36074 56473
rect 35830 56229 35882 56235
rect 35830 56171 35882 56177
rect 35446 56155 35498 56161
rect 35446 56097 35498 56103
rect 34988 55972 35284 55992
rect 35044 55970 35068 55972
rect 35124 55970 35148 55972
rect 35204 55970 35228 55972
rect 35066 55918 35068 55970
rect 35130 55918 35142 55970
rect 35204 55918 35206 55970
rect 35044 55916 35068 55918
rect 35124 55916 35148 55918
rect 35204 55916 35228 55918
rect 34988 55896 35284 55916
rect 34988 54640 35284 54660
rect 35044 54638 35068 54640
rect 35124 54638 35148 54640
rect 35204 54638 35228 54640
rect 35066 54586 35068 54638
rect 35130 54586 35142 54638
rect 35204 54586 35206 54638
rect 35044 54584 35068 54586
rect 35124 54584 35148 54586
rect 35204 54584 35228 54586
rect 34988 54564 35284 54584
rect 34988 53308 35284 53328
rect 35044 53306 35068 53308
rect 35124 53306 35148 53308
rect 35204 53306 35228 53308
rect 35066 53254 35068 53306
rect 35130 53254 35142 53306
rect 35204 53254 35206 53306
rect 35044 53252 35068 53254
rect 35124 53252 35148 53254
rect 35204 53252 35228 53254
rect 34988 53232 35284 53252
rect 34988 51976 35284 51996
rect 35044 51974 35068 51976
rect 35124 51974 35148 51976
rect 35204 51974 35228 51976
rect 35066 51922 35068 51974
rect 35130 51922 35142 51974
rect 35204 51922 35206 51974
rect 35044 51920 35068 51922
rect 35124 51920 35148 51922
rect 35204 51920 35228 51922
rect 34988 51900 35284 51920
rect 34988 50644 35284 50664
rect 35044 50642 35068 50644
rect 35124 50642 35148 50644
rect 35204 50642 35228 50644
rect 35066 50590 35068 50642
rect 35130 50590 35142 50642
rect 35204 50590 35206 50642
rect 35044 50588 35068 50590
rect 35124 50588 35148 50590
rect 35204 50588 35228 50590
rect 34988 50568 35284 50588
rect 34988 49312 35284 49332
rect 35044 49310 35068 49312
rect 35124 49310 35148 49312
rect 35204 49310 35228 49312
rect 35066 49258 35068 49310
rect 35130 49258 35142 49310
rect 35204 49258 35206 49310
rect 35044 49256 35068 49258
rect 35124 49256 35148 49258
rect 35204 49256 35228 49258
rect 34988 49236 35284 49256
rect 34988 47980 35284 48000
rect 35044 47978 35068 47980
rect 35124 47978 35148 47980
rect 35204 47978 35228 47980
rect 35066 47926 35068 47978
rect 35130 47926 35142 47978
rect 35204 47926 35206 47978
rect 35044 47924 35068 47926
rect 35124 47924 35148 47926
rect 35204 47924 35228 47926
rect 34988 47904 35284 47924
rect 34988 46648 35284 46668
rect 35044 46646 35068 46648
rect 35124 46646 35148 46648
rect 35204 46646 35228 46648
rect 35066 46594 35068 46646
rect 35130 46594 35142 46646
rect 35204 46594 35206 46646
rect 35044 46592 35068 46594
rect 35124 46592 35148 46594
rect 35204 46592 35228 46594
rect 34988 46572 35284 46592
rect 34988 45316 35284 45336
rect 35044 45314 35068 45316
rect 35124 45314 35148 45316
rect 35204 45314 35228 45316
rect 35066 45262 35068 45314
rect 35130 45262 35142 45314
rect 35204 45262 35206 45314
rect 35044 45260 35068 45262
rect 35124 45260 35148 45262
rect 35204 45260 35228 45262
rect 34988 45240 35284 45260
rect 34988 43984 35284 44004
rect 35044 43982 35068 43984
rect 35124 43982 35148 43984
rect 35204 43982 35228 43984
rect 35066 43930 35068 43982
rect 35130 43930 35142 43982
rect 35204 43930 35206 43982
rect 35044 43928 35068 43930
rect 35124 43928 35148 43930
rect 35204 43928 35228 43930
rect 34988 43908 35284 43928
rect 34988 42652 35284 42672
rect 35044 42650 35068 42652
rect 35124 42650 35148 42652
rect 35204 42650 35228 42652
rect 35066 42598 35068 42650
rect 35130 42598 35142 42650
rect 35204 42598 35206 42650
rect 35044 42596 35068 42598
rect 35124 42596 35148 42598
rect 35204 42596 35228 42598
rect 34988 42576 35284 42596
rect 34988 41320 35284 41340
rect 35044 41318 35068 41320
rect 35124 41318 35148 41320
rect 35204 41318 35228 41320
rect 35066 41266 35068 41318
rect 35130 41266 35142 41318
rect 35204 41266 35206 41318
rect 35044 41264 35068 41266
rect 35124 41264 35148 41266
rect 35204 41264 35228 41266
rect 34988 41244 35284 41264
rect 34988 39988 35284 40008
rect 35044 39986 35068 39988
rect 35124 39986 35148 39988
rect 35204 39986 35228 39988
rect 35066 39934 35068 39986
rect 35130 39934 35142 39986
rect 35204 39934 35206 39986
rect 35044 39932 35068 39934
rect 35124 39932 35148 39934
rect 35204 39932 35228 39934
rect 34988 39912 35284 39932
rect 34988 38656 35284 38676
rect 35044 38654 35068 38656
rect 35124 38654 35148 38656
rect 35204 38654 35228 38656
rect 35066 38602 35068 38654
rect 35130 38602 35142 38654
rect 35204 38602 35206 38654
rect 35044 38600 35068 38602
rect 35124 38600 35148 38602
rect 35204 38600 35228 38602
rect 34988 38580 35284 38600
rect 34988 37324 35284 37344
rect 35044 37322 35068 37324
rect 35124 37322 35148 37324
rect 35204 37322 35228 37324
rect 35066 37270 35068 37322
rect 35130 37270 35142 37322
rect 35204 37270 35206 37322
rect 35044 37268 35068 37270
rect 35124 37268 35148 37270
rect 35204 37268 35228 37270
rect 34988 37248 35284 37268
rect 34988 35992 35284 36012
rect 35044 35990 35068 35992
rect 35124 35990 35148 35992
rect 35204 35990 35228 35992
rect 35066 35938 35068 35990
rect 35130 35938 35142 35990
rect 35204 35938 35206 35990
rect 35044 35936 35068 35938
rect 35124 35936 35148 35938
rect 35204 35936 35228 35938
rect 34988 35916 35284 35936
rect 34988 34660 35284 34680
rect 35044 34658 35068 34660
rect 35124 34658 35148 34660
rect 35204 34658 35228 34660
rect 35066 34606 35068 34658
rect 35130 34606 35142 34658
rect 35204 34606 35206 34658
rect 35044 34604 35068 34606
rect 35124 34604 35148 34606
rect 35204 34604 35228 34606
rect 34988 34584 35284 34604
rect 34582 33659 34634 33665
rect 34582 33601 34634 33607
rect 34390 23669 34442 23675
rect 34390 23611 34442 23617
rect 34486 9461 34538 9467
rect 34486 9403 34538 9409
rect 34498 7617 34526 9403
rect 34594 7765 34622 33601
rect 34988 33328 35284 33348
rect 35044 33326 35068 33328
rect 35124 33326 35148 33328
rect 35204 33326 35228 33328
rect 35066 33274 35068 33326
rect 35130 33274 35142 33326
rect 35204 33274 35206 33326
rect 35044 33272 35068 33274
rect 35124 33272 35148 33274
rect 35204 33272 35228 33274
rect 34988 33252 35284 33272
rect 34988 31996 35284 32016
rect 35044 31994 35068 31996
rect 35124 31994 35148 31996
rect 35204 31994 35228 31996
rect 35066 31942 35068 31994
rect 35130 31942 35142 31994
rect 35204 31942 35206 31994
rect 35044 31940 35068 31942
rect 35124 31940 35148 31942
rect 35204 31940 35228 31942
rect 34988 31920 35284 31940
rect 35446 30773 35498 30779
rect 35446 30715 35498 30721
rect 34988 30664 35284 30684
rect 35044 30662 35068 30664
rect 35124 30662 35148 30664
rect 35204 30662 35228 30664
rect 35066 30610 35068 30662
rect 35130 30610 35142 30662
rect 35204 30610 35206 30662
rect 35044 30608 35068 30610
rect 35124 30608 35148 30610
rect 35204 30608 35228 30610
rect 34988 30588 35284 30608
rect 34988 29332 35284 29352
rect 35044 29330 35068 29332
rect 35124 29330 35148 29332
rect 35204 29330 35228 29332
rect 35066 29278 35068 29330
rect 35130 29278 35142 29330
rect 35204 29278 35206 29330
rect 35044 29276 35068 29278
rect 35124 29276 35148 29278
rect 35204 29276 35228 29278
rect 34988 29256 35284 29276
rect 34988 28000 35284 28020
rect 35044 27998 35068 28000
rect 35124 27998 35148 28000
rect 35204 27998 35228 28000
rect 35066 27946 35068 27998
rect 35130 27946 35142 27998
rect 35204 27946 35206 27998
rect 35044 27944 35068 27946
rect 35124 27944 35148 27946
rect 35204 27944 35228 27946
rect 34988 27924 35284 27944
rect 34870 26925 34922 26931
rect 34870 26867 34922 26873
rect 34774 19599 34826 19605
rect 34774 19541 34826 19547
rect 34786 19161 34814 19541
rect 34774 19155 34826 19161
rect 34774 19097 34826 19103
rect 34582 7759 34634 7765
rect 34582 7701 34634 7707
rect 34486 7611 34538 7617
rect 34486 7553 34538 7559
rect 34390 7463 34442 7469
rect 34390 7405 34442 7411
rect 34774 7463 34826 7469
rect 34774 7405 34826 7411
rect 34198 6427 34250 6433
rect 34198 6369 34250 6375
rect 34294 6131 34346 6137
rect 34294 6073 34346 6079
rect 34102 5021 34154 5027
rect 34102 4963 34154 4969
rect 34114 3251 34142 4963
rect 34198 4281 34250 4287
rect 34198 4223 34250 4229
rect 34102 3245 34154 3251
rect 34102 3187 34154 3193
rect 34210 2894 34238 4223
rect 34306 3917 34334 6073
rect 34294 3911 34346 3917
rect 34294 3853 34346 3859
rect 34294 3689 34346 3695
rect 34294 3631 34346 3637
rect 34114 2866 34238 2894
rect 34114 800 34142 2866
rect 34306 800 34334 3631
rect 34402 800 34430 7405
rect 34678 5687 34730 5693
rect 34678 5629 34730 5635
rect 34582 4947 34634 4953
rect 34582 4889 34634 4895
rect 34594 4528 34622 4889
rect 34498 4500 34622 4528
rect 34498 800 34526 4500
rect 34582 4355 34634 4361
rect 34582 4297 34634 4303
rect 34594 800 34622 4297
rect 34690 3177 34718 5629
rect 34678 3171 34730 3177
rect 34678 3113 34730 3119
rect 34786 800 34814 7405
rect 34882 6581 34910 26867
rect 34988 26668 35284 26688
rect 35044 26666 35068 26668
rect 35124 26666 35148 26668
rect 35204 26666 35228 26668
rect 35066 26614 35068 26666
rect 35130 26614 35142 26666
rect 35204 26614 35206 26666
rect 35044 26612 35068 26614
rect 35124 26612 35148 26614
rect 35204 26612 35228 26614
rect 34988 26592 35284 26612
rect 34988 25336 35284 25356
rect 35044 25334 35068 25336
rect 35124 25334 35148 25336
rect 35204 25334 35228 25336
rect 35066 25282 35068 25334
rect 35130 25282 35142 25334
rect 35204 25282 35206 25334
rect 35044 25280 35068 25282
rect 35124 25280 35148 25282
rect 35204 25280 35228 25282
rect 34988 25260 35284 25280
rect 35350 24187 35402 24193
rect 35350 24129 35402 24135
rect 34988 24004 35284 24024
rect 35044 24002 35068 24004
rect 35124 24002 35148 24004
rect 35204 24002 35228 24004
rect 35066 23950 35068 24002
rect 35130 23950 35142 24002
rect 35204 23950 35206 24002
rect 35044 23948 35068 23950
rect 35124 23948 35148 23950
rect 35204 23948 35228 23950
rect 34988 23928 35284 23948
rect 34988 22672 35284 22692
rect 35044 22670 35068 22672
rect 35124 22670 35148 22672
rect 35204 22670 35228 22672
rect 35066 22618 35068 22670
rect 35130 22618 35142 22670
rect 35204 22618 35206 22670
rect 35044 22616 35068 22618
rect 35124 22616 35148 22618
rect 35204 22616 35228 22618
rect 34988 22596 35284 22616
rect 34988 21340 35284 21360
rect 35044 21338 35068 21340
rect 35124 21338 35148 21340
rect 35204 21338 35228 21340
rect 35066 21286 35068 21338
rect 35130 21286 35142 21338
rect 35204 21286 35206 21338
rect 35044 21284 35068 21286
rect 35124 21284 35148 21286
rect 35204 21284 35228 21286
rect 34988 21264 35284 21284
rect 34988 20008 35284 20028
rect 35044 20006 35068 20008
rect 35124 20006 35148 20008
rect 35204 20006 35228 20008
rect 35066 19954 35068 20006
rect 35130 19954 35142 20006
rect 35204 19954 35206 20006
rect 35044 19952 35068 19954
rect 35124 19952 35148 19954
rect 35204 19952 35228 19954
rect 34988 19932 35284 19952
rect 34988 18676 35284 18696
rect 35044 18674 35068 18676
rect 35124 18674 35148 18676
rect 35204 18674 35228 18676
rect 35066 18622 35068 18674
rect 35130 18622 35142 18674
rect 35204 18622 35206 18674
rect 35044 18620 35068 18622
rect 35124 18620 35148 18622
rect 35204 18620 35228 18622
rect 34988 18600 35284 18620
rect 34988 17344 35284 17364
rect 35044 17342 35068 17344
rect 35124 17342 35148 17344
rect 35204 17342 35228 17344
rect 35066 17290 35068 17342
rect 35130 17290 35142 17342
rect 35204 17290 35206 17342
rect 35044 17288 35068 17290
rect 35124 17288 35148 17290
rect 35204 17288 35228 17290
rect 34988 17268 35284 17288
rect 34988 16012 35284 16032
rect 35044 16010 35068 16012
rect 35124 16010 35148 16012
rect 35204 16010 35228 16012
rect 35066 15958 35068 16010
rect 35130 15958 35142 16010
rect 35204 15958 35206 16010
rect 35044 15956 35068 15958
rect 35124 15956 35148 15958
rect 35204 15956 35228 15958
rect 34988 15936 35284 15956
rect 34988 14680 35284 14700
rect 35044 14678 35068 14680
rect 35124 14678 35148 14680
rect 35204 14678 35228 14680
rect 35066 14626 35068 14678
rect 35130 14626 35142 14678
rect 35204 14626 35206 14678
rect 35044 14624 35068 14626
rect 35124 14624 35148 14626
rect 35204 14624 35228 14626
rect 34988 14604 35284 14624
rect 34988 13348 35284 13368
rect 35044 13346 35068 13348
rect 35124 13346 35148 13348
rect 35204 13346 35228 13348
rect 35066 13294 35068 13346
rect 35130 13294 35142 13346
rect 35204 13294 35206 13346
rect 35044 13292 35068 13294
rect 35124 13292 35148 13294
rect 35204 13292 35228 13294
rect 34988 13272 35284 13292
rect 34988 12016 35284 12036
rect 35044 12014 35068 12016
rect 35124 12014 35148 12016
rect 35204 12014 35228 12016
rect 35066 11962 35068 12014
rect 35130 11962 35142 12014
rect 35204 11962 35206 12014
rect 35044 11960 35068 11962
rect 35124 11960 35148 11962
rect 35204 11960 35228 11962
rect 34988 11940 35284 11960
rect 34988 10684 35284 10704
rect 35044 10682 35068 10684
rect 35124 10682 35148 10684
rect 35204 10682 35228 10684
rect 35066 10630 35068 10682
rect 35130 10630 35142 10682
rect 35204 10630 35206 10682
rect 35044 10628 35068 10630
rect 35124 10628 35148 10630
rect 35204 10628 35228 10630
rect 34988 10608 35284 10628
rect 34988 9352 35284 9372
rect 35044 9350 35068 9352
rect 35124 9350 35148 9352
rect 35204 9350 35228 9352
rect 35066 9298 35068 9350
rect 35130 9298 35142 9350
rect 35204 9298 35206 9350
rect 35044 9296 35068 9298
rect 35124 9296 35148 9298
rect 35204 9296 35228 9298
rect 34988 9276 35284 9296
rect 34988 8020 35284 8040
rect 35044 8018 35068 8020
rect 35124 8018 35148 8020
rect 35204 8018 35228 8020
rect 35066 7966 35068 8018
rect 35130 7966 35142 8018
rect 35204 7966 35206 8018
rect 35044 7964 35068 7966
rect 35124 7964 35148 7966
rect 35204 7964 35228 7966
rect 34988 7944 35284 7964
rect 35362 7765 35390 24129
rect 35458 9467 35486 30715
rect 35842 17681 35870 56171
rect 36502 54157 36554 54163
rect 36502 54099 36554 54105
rect 36118 31735 36170 31741
rect 36118 31677 36170 31683
rect 35830 17675 35882 17681
rect 35830 17617 35882 17623
rect 36022 10793 36074 10799
rect 36022 10735 36074 10741
rect 35446 9461 35498 9467
rect 35446 9403 35498 9409
rect 35350 7759 35402 7765
rect 35350 7701 35402 7707
rect 35830 7463 35882 7469
rect 35830 7405 35882 7411
rect 35542 6945 35594 6951
rect 35542 6887 35594 6893
rect 34988 6688 35284 6708
rect 35044 6686 35068 6688
rect 35124 6686 35148 6688
rect 35204 6686 35228 6688
rect 35066 6634 35068 6686
rect 35130 6634 35142 6686
rect 35204 6634 35206 6686
rect 35044 6632 35068 6634
rect 35124 6632 35148 6634
rect 35204 6632 35228 6634
rect 34988 6612 35284 6632
rect 34870 6575 34922 6581
rect 34870 6517 34922 6523
rect 34988 5356 35284 5376
rect 35044 5354 35068 5356
rect 35124 5354 35148 5356
rect 35204 5354 35228 5356
rect 35066 5302 35068 5354
rect 35130 5302 35142 5354
rect 35204 5302 35206 5354
rect 35044 5300 35068 5302
rect 35124 5300 35148 5302
rect 35204 5300 35228 5302
rect 34988 5280 35284 5300
rect 34870 5021 34922 5027
rect 34870 4963 34922 4969
rect 34882 3843 34910 4963
rect 35350 4503 35402 4509
rect 35350 4445 35402 4451
rect 34988 4024 35284 4044
rect 35044 4022 35068 4024
rect 35124 4022 35148 4024
rect 35204 4022 35228 4024
rect 35066 3970 35068 4022
rect 35130 3970 35142 4022
rect 35204 3970 35206 4022
rect 35044 3968 35068 3970
rect 35124 3968 35148 3970
rect 35204 3968 35228 3970
rect 34988 3948 35284 3968
rect 34870 3837 34922 3843
rect 34870 3779 34922 3785
rect 34966 3689 35018 3695
rect 34882 3649 34966 3677
rect 34882 1420 34910 3649
rect 34966 3631 35018 3637
rect 35362 3196 35390 4445
rect 35266 3168 35390 3196
rect 35266 2881 35294 3168
rect 35446 3023 35498 3029
rect 35446 2965 35498 2971
rect 35350 2949 35402 2955
rect 35350 2891 35402 2897
rect 35254 2875 35306 2881
rect 35254 2817 35306 2823
rect 34988 2692 35284 2712
rect 35044 2690 35068 2692
rect 35124 2690 35148 2692
rect 35204 2690 35228 2692
rect 35066 2638 35068 2690
rect 35130 2638 35142 2690
rect 35204 2638 35206 2690
rect 35044 2636 35068 2638
rect 35124 2636 35148 2638
rect 35204 2636 35228 2638
rect 34988 2616 35284 2636
rect 35362 1568 35390 2891
rect 35266 1540 35390 1568
rect 35158 1469 35210 1475
rect 34882 1392 35006 1420
rect 35158 1411 35210 1417
rect 34870 1321 34922 1327
rect 34870 1263 34922 1269
rect 34882 800 34910 1263
rect 34978 800 35006 1392
rect 35170 800 35198 1411
rect 35266 800 35294 1540
rect 35458 1420 35486 2965
rect 35554 1475 35582 6887
rect 35734 3689 35786 3695
rect 35734 3631 35786 3637
rect 35638 3097 35690 3103
rect 35638 3039 35690 3045
rect 35650 1623 35678 3039
rect 35638 1617 35690 1623
rect 35638 1559 35690 1565
rect 35362 1392 35486 1420
rect 35542 1469 35594 1475
rect 35542 1411 35594 1417
rect 35638 1469 35690 1475
rect 35638 1411 35690 1417
rect 35362 800 35390 1392
rect 35446 1099 35498 1105
rect 35446 1041 35498 1047
rect 35458 800 35486 1041
rect 35650 800 35678 1411
rect 35746 800 35774 3631
rect 35842 800 35870 7405
rect 36034 7099 36062 10735
rect 36130 7765 36158 31677
rect 36214 26777 36266 26783
rect 36214 26719 36266 26725
rect 36226 17294 36254 26719
rect 36226 17266 36350 17294
rect 36214 13161 36266 13167
rect 36214 13103 36266 13109
rect 36118 7759 36170 7765
rect 36118 7701 36170 7707
rect 36226 7543 36254 13103
rect 36322 9171 36350 17266
rect 36310 9165 36362 9171
rect 36310 9107 36362 9113
rect 36514 7913 36542 54099
rect 36598 34843 36650 34849
rect 36598 34785 36650 34791
rect 36502 7907 36554 7913
rect 36502 7849 36554 7855
rect 36514 7765 36542 7849
rect 36502 7759 36554 7765
rect 36502 7701 36554 7707
rect 36214 7537 36266 7543
rect 36214 7479 36266 7485
rect 36610 7173 36638 34785
rect 36706 15535 36734 56689
rect 36790 56229 36842 56235
rect 36790 56171 36842 56177
rect 36694 15529 36746 15535
rect 36694 15471 36746 15477
rect 36802 14129 36830 56171
rect 37090 56161 37118 57586
rect 37570 56531 37598 59200
rect 38050 56975 38078 59200
rect 38038 56969 38090 56975
rect 38038 56911 38090 56917
rect 38626 56531 38654 59200
rect 37558 56525 37610 56531
rect 37558 56467 37610 56473
rect 38614 56525 38666 56531
rect 38614 56467 38666 56473
rect 37750 56229 37802 56235
rect 37750 56171 37802 56177
rect 38710 56229 38762 56235
rect 38710 56171 38762 56177
rect 37078 56155 37130 56161
rect 37078 56097 37130 56103
rect 36886 54157 36938 54163
rect 36886 54099 36938 54105
rect 36790 14123 36842 14129
rect 36790 14065 36842 14071
rect 36694 7463 36746 7469
rect 36694 7405 36746 7411
rect 36598 7167 36650 7173
rect 36598 7109 36650 7115
rect 36022 7093 36074 7099
rect 36022 7035 36074 7041
rect 36406 6945 36458 6951
rect 36406 6887 36458 6893
rect 36310 6353 36362 6359
rect 36310 6295 36362 6301
rect 36022 5687 36074 5693
rect 36022 5629 36074 5635
rect 36214 5687 36266 5693
rect 36214 5629 36266 5635
rect 35926 3171 35978 3177
rect 35926 3113 35978 3119
rect 35938 1475 35966 3113
rect 36034 2955 36062 5629
rect 36118 5021 36170 5027
rect 36118 4963 36170 4969
rect 36130 3103 36158 4963
rect 36118 3097 36170 3103
rect 36118 3039 36170 3045
rect 36022 2949 36074 2955
rect 36022 2891 36074 2897
rect 36118 2949 36170 2955
rect 36118 2891 36170 2897
rect 36130 1697 36158 2891
rect 36118 1691 36170 1697
rect 36118 1633 36170 1639
rect 35926 1469 35978 1475
rect 36226 1420 36254 5629
rect 36322 1549 36350 6295
rect 36310 1543 36362 1549
rect 36310 1485 36362 1491
rect 35926 1411 35978 1417
rect 36034 1392 36254 1420
rect 36034 800 36062 1392
rect 36118 1321 36170 1327
rect 36418 1272 36446 6887
rect 36502 3689 36554 3695
rect 36706 3640 36734 7405
rect 36898 6581 36926 54099
rect 37462 44759 37514 44765
rect 37462 44701 37514 44707
rect 37474 7173 37502 44701
rect 37762 26265 37790 56171
rect 38422 49421 38474 49427
rect 38422 49363 38474 49369
rect 38434 49057 38462 49363
rect 38422 49051 38474 49057
rect 38422 48993 38474 48999
rect 37750 26259 37802 26265
rect 37750 26201 37802 26207
rect 37558 22781 37610 22787
rect 37558 22723 37610 22729
rect 37570 22565 37598 22723
rect 37558 22559 37610 22565
rect 37558 22501 37610 22507
rect 38518 11607 38570 11613
rect 38518 11549 38570 11555
rect 38038 7463 38090 7469
rect 38038 7405 38090 7411
rect 37462 7167 37514 7173
rect 37462 7109 37514 7115
rect 37078 6945 37130 6951
rect 37078 6887 37130 6893
rect 36886 6575 36938 6581
rect 36886 6517 36938 6523
rect 36886 5021 36938 5027
rect 36886 4963 36938 4969
rect 36790 4355 36842 4361
rect 36790 4297 36842 4303
rect 36502 3631 36554 3637
rect 36118 1263 36170 1269
rect 36130 800 36158 1263
rect 36226 1244 36446 1272
rect 36226 800 36254 1244
rect 36310 1173 36362 1179
rect 36310 1115 36362 1121
rect 36322 800 36350 1115
rect 36514 800 36542 3631
rect 36610 3612 36734 3640
rect 36610 800 36638 3612
rect 36694 3097 36746 3103
rect 36694 3039 36746 3045
rect 36706 800 36734 3039
rect 36802 800 36830 4297
rect 36898 3177 36926 4963
rect 37090 3492 37118 6887
rect 37366 6871 37418 6877
rect 37366 6813 37418 6819
rect 37270 6131 37322 6137
rect 37270 6073 37322 6079
rect 37174 4281 37226 4287
rect 37174 4223 37226 4229
rect 36994 3464 37118 3492
rect 36886 3171 36938 3177
rect 36886 3113 36938 3119
rect 36994 800 37022 3464
rect 37078 3171 37130 3177
rect 37078 3113 37130 3119
rect 37090 800 37118 3113
rect 37186 800 37214 4223
rect 37282 1105 37310 6073
rect 37270 1099 37322 1105
rect 37270 1041 37322 1047
rect 37378 800 37406 6813
rect 37654 6797 37706 6803
rect 37654 6739 37706 6745
rect 37558 5687 37610 5693
rect 37558 5629 37610 5635
rect 37462 5539 37514 5545
rect 37462 5481 37514 5487
rect 37474 800 37502 5481
rect 37570 3103 37598 5629
rect 37558 3097 37610 3103
rect 37558 3039 37610 3045
rect 37558 2949 37610 2955
rect 37558 2891 37610 2897
rect 37570 800 37598 2891
rect 37666 800 37694 6739
rect 37846 3837 37898 3843
rect 37846 3779 37898 3785
rect 37858 800 37886 3779
rect 37942 3689 37994 3695
rect 37942 3631 37994 3637
rect 37954 800 37982 3631
rect 38050 800 38078 7405
rect 38530 7099 38558 11549
rect 38518 7093 38570 7099
rect 38518 7035 38570 7041
rect 38518 6945 38570 6951
rect 38434 6905 38518 6933
rect 38326 3097 38378 3103
rect 38326 3039 38378 3045
rect 38134 2949 38186 2955
rect 38134 2891 38186 2897
rect 38146 800 38174 2891
rect 38338 800 38366 3039
rect 38434 800 38462 6905
rect 38518 6887 38570 6893
rect 38614 5021 38666 5027
rect 38614 4963 38666 4969
rect 38518 4207 38570 4213
rect 38518 4149 38570 4155
rect 38530 800 38558 4149
rect 38626 3177 38654 4963
rect 38722 3917 38750 56171
rect 38806 56081 38858 56087
rect 38806 56023 38858 56029
rect 38818 55495 38846 56023
rect 39106 55717 39134 59200
rect 39682 56901 39710 59200
rect 39670 56895 39722 56901
rect 39670 56837 39722 56843
rect 39766 56747 39818 56753
rect 39766 56689 39818 56695
rect 39094 55711 39146 55717
rect 39094 55653 39146 55659
rect 38806 55489 38858 55495
rect 38806 55431 38858 55437
rect 38902 55415 38954 55421
rect 38902 55357 38954 55363
rect 38914 15461 38942 55357
rect 39670 42243 39722 42249
rect 39670 42185 39722 42191
rect 39286 32105 39338 32111
rect 39286 32047 39338 32053
rect 38902 15455 38954 15461
rect 38902 15397 38954 15403
rect 38806 7463 38858 7469
rect 38806 7405 38858 7411
rect 38710 3911 38762 3917
rect 38710 3853 38762 3859
rect 38710 3689 38762 3695
rect 38710 3631 38762 3637
rect 38614 3171 38666 3177
rect 38614 3113 38666 3119
rect 38722 800 38750 3631
rect 38818 800 38846 7405
rect 39298 7099 39326 32047
rect 39574 7463 39626 7469
rect 39574 7405 39626 7411
rect 39586 7214 39614 7405
rect 39490 7186 39614 7214
rect 39286 7093 39338 7099
rect 39286 7035 39338 7041
rect 38902 6353 38954 6359
rect 38902 6295 38954 6301
rect 38914 800 38942 6295
rect 39190 6131 39242 6137
rect 39190 6073 39242 6079
rect 39094 5687 39146 5693
rect 39094 5629 39146 5635
rect 38998 4355 39050 4361
rect 38998 4297 39050 4303
rect 39010 800 39038 4297
rect 39106 2955 39134 5629
rect 39094 2949 39146 2955
rect 39094 2891 39146 2897
rect 39202 800 39230 6073
rect 39286 5687 39338 5693
rect 39286 5629 39338 5635
rect 39298 800 39326 5629
rect 39382 5021 39434 5027
rect 39382 4963 39434 4969
rect 39394 3843 39422 4963
rect 39382 3837 39434 3843
rect 39382 3779 39434 3785
rect 39382 3541 39434 3547
rect 39382 3483 39434 3489
rect 39394 800 39422 3483
rect 39490 800 39518 7186
rect 39682 7173 39710 42185
rect 39778 16867 39806 56689
rect 40162 56531 40190 59200
rect 40630 56895 40682 56901
rect 40630 56837 40682 56843
rect 40342 56821 40394 56827
rect 40342 56763 40394 56769
rect 40150 56525 40202 56531
rect 40150 56467 40202 56473
rect 39862 56229 39914 56235
rect 39862 56171 39914 56177
rect 39874 18939 39902 56171
rect 40354 49205 40382 56763
rect 40438 55415 40490 55421
rect 40438 55357 40490 55363
rect 40342 49199 40394 49205
rect 40342 49141 40394 49147
rect 40342 19821 40394 19827
rect 40342 19763 40394 19769
rect 39862 18933 39914 18939
rect 39862 18875 39914 18881
rect 39766 16861 39818 16867
rect 39766 16803 39818 16809
rect 40354 7765 40382 19763
rect 40450 11687 40478 55357
rect 40642 47534 40670 56837
rect 40738 55717 40766 59200
rect 41218 56975 41246 59200
rect 41206 56969 41258 56975
rect 41206 56911 41258 56917
rect 40822 56747 40874 56753
rect 40822 56689 40874 56695
rect 40834 56161 40862 56689
rect 41794 56531 41822 59200
rect 42274 56531 42302 59200
rect 42850 56901 42878 59200
rect 42838 56895 42890 56901
rect 42838 56837 42890 56843
rect 42934 56747 42986 56753
rect 42934 56689 42986 56695
rect 41782 56525 41834 56531
rect 41782 56467 41834 56473
rect 42262 56525 42314 56531
rect 42262 56467 42314 56473
rect 42550 56303 42602 56309
rect 42550 56245 42602 56251
rect 41974 56229 42026 56235
rect 41974 56171 42026 56177
rect 40822 56155 40874 56161
rect 40822 56097 40874 56103
rect 40726 55711 40778 55717
rect 40726 55653 40778 55659
rect 40642 47506 40766 47534
rect 40738 25599 40766 47506
rect 41986 46245 42014 56171
rect 42166 55415 42218 55421
rect 42166 55357 42218 55363
rect 41974 46239 42026 46245
rect 41974 46181 42026 46187
rect 41110 46165 41162 46171
rect 41110 46107 41162 46113
rect 41014 45425 41066 45431
rect 41014 45367 41066 45373
rect 40726 25593 40778 25599
rect 40726 25535 40778 25541
rect 40726 18267 40778 18273
rect 40726 18209 40778 18215
rect 40438 11681 40490 11687
rect 40438 11623 40490 11629
rect 40738 10799 40766 18209
rect 40726 10793 40778 10799
rect 40726 10735 40778 10741
rect 41026 7913 41054 45367
rect 41014 7907 41066 7913
rect 41014 7849 41066 7855
rect 40342 7759 40394 7765
rect 40342 7701 40394 7707
rect 40246 7685 40298 7691
rect 40246 7627 40298 7633
rect 39670 7167 39722 7173
rect 39670 7109 39722 7115
rect 39862 6871 39914 6877
rect 39862 6813 39914 6819
rect 39766 4355 39818 4361
rect 39766 4297 39818 4303
rect 39670 3097 39722 3103
rect 39670 3039 39722 3045
rect 39682 800 39710 3039
rect 39778 800 39806 4297
rect 39874 800 39902 6813
rect 40150 5021 40202 5027
rect 40150 4963 40202 4969
rect 40162 4213 40190 4963
rect 40150 4207 40202 4213
rect 40150 4149 40202 4155
rect 40054 3911 40106 3917
rect 40054 3853 40106 3859
rect 40066 800 40094 3853
rect 40150 3541 40202 3547
rect 40150 3483 40202 3489
rect 40162 800 40190 3483
rect 40258 800 40286 7627
rect 41026 7617 41054 7849
rect 41014 7611 41066 7617
rect 41014 7553 41066 7559
rect 41122 7173 41150 46107
rect 41878 23595 41930 23601
rect 41878 23537 41930 23543
rect 41782 9461 41834 9467
rect 41782 9403 41834 9409
rect 41398 7463 41450 7469
rect 41398 7405 41450 7411
rect 41110 7167 41162 7173
rect 41110 7109 41162 7115
rect 41206 7019 41258 7025
rect 41206 6961 41258 6967
rect 40342 6353 40394 6359
rect 40342 6295 40394 6301
rect 40354 800 40382 6295
rect 40630 6205 40682 6211
rect 40630 6147 40682 6153
rect 40534 3023 40586 3029
rect 40534 2965 40586 2971
rect 40546 800 40574 2965
rect 40642 800 40670 6147
rect 40726 5687 40778 5693
rect 40726 5629 40778 5635
rect 40738 800 40766 5629
rect 40918 5021 40970 5027
rect 40918 4963 40970 4969
rect 40930 3103 40958 4963
rect 41014 3689 41066 3695
rect 41014 3631 41066 3637
rect 40918 3097 40970 3103
rect 40918 3039 40970 3045
rect 41026 2900 41054 3631
rect 41218 3547 41246 6961
rect 41302 6871 41354 6877
rect 41302 6813 41354 6819
rect 41206 3541 41258 3547
rect 41206 3483 41258 3489
rect 41110 3097 41162 3103
rect 41110 3039 41162 3045
rect 40930 2872 41054 2900
rect 40930 800 40958 2872
rect 41014 2801 41066 2807
rect 41014 2743 41066 2749
rect 41026 2437 41054 2743
rect 41014 2431 41066 2437
rect 41014 2373 41066 2379
rect 41014 1469 41066 1475
rect 41014 1411 41066 1417
rect 41026 800 41054 1411
rect 41122 800 41150 3039
rect 41206 2949 41258 2955
rect 41206 2891 41258 2897
rect 41218 800 41246 2891
rect 41314 1475 41342 6813
rect 41302 1469 41354 1475
rect 41302 1411 41354 1417
rect 41410 800 41438 7405
rect 41794 7173 41822 9403
rect 41890 7765 41918 23537
rect 41878 7759 41930 7765
rect 41878 7701 41930 7707
rect 42178 7691 42206 55357
rect 42262 50457 42314 50463
rect 42262 50399 42314 50405
rect 42274 7913 42302 50399
rect 42562 47534 42590 56245
rect 42646 56229 42698 56235
rect 42646 56171 42698 56177
rect 42466 47506 42590 47534
rect 42466 12205 42494 47506
rect 42658 16793 42686 56171
rect 42838 52085 42890 52091
rect 42838 52027 42890 52033
rect 42742 40911 42794 40917
rect 42742 40853 42794 40859
rect 42646 16787 42698 16793
rect 42646 16729 42698 16735
rect 42454 12199 42506 12205
rect 42454 12141 42506 12147
rect 42262 7907 42314 7913
rect 42262 7849 42314 7855
rect 42274 7765 42302 7849
rect 42262 7759 42314 7765
rect 42262 7701 42314 7707
rect 42166 7685 42218 7691
rect 42166 7627 42218 7633
rect 42454 7463 42506 7469
rect 42454 7405 42506 7411
rect 41782 7167 41834 7173
rect 41782 7109 41834 7115
rect 41878 6353 41930 6359
rect 41878 6295 41930 6301
rect 41782 5687 41834 5693
rect 41782 5629 41834 5635
rect 41686 5021 41738 5027
rect 41686 4963 41738 4969
rect 41698 3917 41726 4963
rect 41686 3911 41738 3917
rect 41686 3853 41738 3859
rect 41794 3788 41822 5629
rect 41506 3760 41822 3788
rect 41506 800 41534 3760
rect 41590 3615 41642 3621
rect 41590 3557 41642 3563
rect 41602 800 41630 3557
rect 41686 3541 41738 3547
rect 41686 3483 41738 3489
rect 41698 800 41726 3483
rect 41890 800 41918 6295
rect 42166 6205 42218 6211
rect 42166 6147 42218 6153
rect 42070 5021 42122 5027
rect 42070 4963 42122 4969
rect 41974 4355 42026 4361
rect 41974 4297 42026 4303
rect 41986 800 42014 4297
rect 42082 3103 42110 4963
rect 42070 3097 42122 3103
rect 42070 3039 42122 3045
rect 42178 2900 42206 6147
rect 42262 5687 42314 5693
rect 42262 5629 42314 5635
rect 42082 2872 42206 2900
rect 42082 800 42110 2872
rect 42274 800 42302 5629
rect 42358 4355 42410 4361
rect 42358 4297 42410 4303
rect 42370 800 42398 4297
rect 42466 800 42494 7405
rect 42754 6433 42782 40853
rect 42850 9911 42878 52027
rect 42946 17755 42974 56689
rect 43330 56531 43358 59200
rect 43906 56531 43934 59200
rect 44386 56975 44414 59200
rect 44374 56969 44426 56975
rect 44374 56911 44426 56917
rect 44962 56531 44990 59200
rect 43318 56525 43370 56531
rect 43318 56467 43370 56473
rect 43894 56525 43946 56531
rect 43894 56467 43946 56473
rect 44950 56525 45002 56531
rect 44950 56467 45002 56473
rect 43894 56377 43946 56383
rect 43894 56319 43946 56325
rect 43606 56229 43658 56235
rect 43606 56171 43658 56177
rect 43414 34843 43466 34849
rect 43414 34785 43466 34791
rect 43126 33437 43178 33443
rect 43126 33379 43178 33385
rect 43138 33221 43166 33379
rect 43126 33215 43178 33221
rect 43126 33157 43178 33163
rect 42934 17749 42986 17755
rect 42934 17691 42986 17697
rect 42934 11903 42986 11909
rect 42934 11845 42986 11851
rect 42838 9905 42890 9911
rect 42838 9847 42890 9853
rect 42946 7099 42974 11845
rect 43426 7173 43454 34785
rect 43618 9541 43646 56171
rect 43906 21677 43934 56319
rect 44182 56229 44234 56235
rect 44182 56171 44234 56177
rect 45046 56229 45098 56235
rect 45046 56171 45098 56177
rect 43894 21671 43946 21677
rect 43894 21613 43946 21619
rect 44194 20197 44222 56171
rect 44662 54749 44714 54755
rect 44662 54691 44714 54697
rect 44182 20191 44234 20197
rect 44182 20133 44234 20139
rect 44674 9689 44702 54691
rect 44854 44759 44906 44765
rect 44854 44701 44906 44707
rect 44758 24113 44810 24119
rect 44758 24055 44810 24061
rect 44662 9683 44714 9689
rect 44662 9625 44714 9631
rect 43606 9535 43658 9541
rect 43606 9477 43658 9483
rect 44086 8943 44138 8949
rect 44086 8885 44138 8891
rect 44098 7765 44126 8885
rect 44086 7759 44138 7765
rect 44086 7701 44138 7707
rect 43894 7463 43946 7469
rect 43894 7405 43946 7411
rect 44662 7463 44714 7469
rect 44662 7405 44714 7411
rect 43414 7167 43466 7173
rect 43414 7109 43466 7115
rect 42934 7093 42986 7099
rect 42934 7035 42986 7041
rect 42838 6871 42890 6877
rect 42838 6813 42890 6819
rect 42742 6427 42794 6433
rect 42742 6369 42794 6375
rect 42742 3689 42794 3695
rect 42742 3631 42794 3637
rect 42550 3097 42602 3103
rect 42550 3039 42602 3045
rect 42562 800 42590 3039
rect 42754 800 42782 3631
rect 42850 800 42878 6813
rect 43606 6797 43658 6803
rect 43606 6739 43658 6745
rect 43222 5687 43274 5693
rect 43222 5629 43274 5635
rect 43234 2900 43262 5629
rect 43318 5021 43370 5027
rect 43318 4963 43370 4969
rect 43330 3103 43358 4963
rect 43414 4355 43466 4361
rect 43414 4297 43466 4303
rect 43318 3097 43370 3103
rect 43318 3039 43370 3045
rect 42946 2872 43262 2900
rect 43318 2949 43370 2955
rect 43318 2891 43370 2897
rect 42946 800 42974 2872
rect 43030 2801 43082 2807
rect 43030 2743 43082 2749
rect 43222 2801 43274 2807
rect 43222 2743 43274 2749
rect 43042 800 43070 2743
rect 43234 800 43262 2743
rect 43330 800 43358 2891
rect 43426 800 43454 4297
rect 43510 3467 43562 3473
rect 43510 3409 43562 3415
rect 43522 2955 43550 3409
rect 43510 2949 43562 2955
rect 43510 2891 43562 2897
rect 43618 800 43646 6739
rect 43798 6279 43850 6285
rect 43798 6221 43850 6227
rect 43702 5687 43754 5693
rect 43702 5629 43754 5635
rect 43714 800 43742 5629
rect 43810 4287 43838 6221
rect 43798 4281 43850 4287
rect 43798 4223 43850 4229
rect 43798 3615 43850 3621
rect 43798 3557 43850 3563
rect 43810 800 43838 3557
rect 43906 800 43934 7405
rect 44566 6871 44618 6877
rect 44290 6831 44566 6859
rect 44086 6279 44138 6285
rect 44086 6221 44138 6227
rect 44098 5915 44126 6221
rect 44182 6131 44234 6137
rect 44182 6073 44234 6079
rect 44086 5909 44138 5915
rect 44086 5851 44138 5857
rect 44194 3344 44222 6073
rect 44002 3316 44222 3344
rect 44002 2955 44030 3316
rect 44086 3171 44138 3177
rect 44086 3113 44138 3119
rect 43990 2949 44042 2955
rect 43990 2891 44042 2897
rect 44098 800 44126 3113
rect 44182 2949 44234 2955
rect 44182 2891 44234 2897
rect 44194 800 44222 2891
rect 44290 800 44318 6831
rect 44566 6813 44618 6819
rect 44566 3763 44618 3769
rect 44566 3705 44618 3711
rect 44470 3097 44522 3103
rect 44470 3039 44522 3045
rect 44482 800 44510 3039
rect 44578 800 44606 3705
rect 44674 800 44702 7405
rect 44770 6433 44798 24055
rect 44866 7765 44894 44701
rect 45058 14573 45086 56171
rect 45442 55717 45470 59200
rect 45922 56883 45950 59200
rect 46102 56895 46154 56901
rect 45922 56855 46102 56883
rect 46102 56837 46154 56843
rect 46102 56747 46154 56753
rect 46102 56689 46154 56695
rect 45430 55711 45482 55717
rect 45430 55653 45482 55659
rect 45238 55415 45290 55421
rect 45238 55357 45290 55363
rect 45142 40763 45194 40769
rect 45142 40705 45194 40711
rect 45046 14567 45098 14573
rect 45046 14509 45098 14515
rect 44950 8129 45002 8135
rect 44950 8071 45002 8077
rect 44854 7759 44906 7765
rect 44854 7701 44906 7707
rect 44758 6427 44810 6433
rect 44758 6369 44810 6375
rect 44962 5767 44990 8071
rect 45046 7759 45098 7765
rect 45046 7701 45098 7707
rect 44950 5761 45002 5767
rect 44950 5703 45002 5709
rect 44758 5021 44810 5027
rect 44758 4963 44810 4969
rect 44770 3473 44798 4963
rect 44950 4355 45002 4361
rect 44950 4297 45002 4303
rect 44758 3467 44810 3473
rect 44758 3409 44810 3415
rect 44758 3245 44810 3251
rect 44758 3187 44810 3193
rect 44770 800 44798 3187
rect 44962 800 44990 4297
rect 45058 800 45086 7701
rect 45154 7173 45182 40705
rect 45250 18495 45278 55357
rect 46114 19531 46142 56689
rect 46498 56531 46526 59200
rect 46486 56525 46538 56531
rect 46486 56467 46538 56473
rect 46774 56229 46826 56235
rect 46774 56171 46826 56177
rect 46582 55415 46634 55421
rect 46582 55357 46634 55363
rect 46294 42095 46346 42101
rect 46294 42037 46346 42043
rect 46198 41207 46250 41213
rect 46198 41149 46250 41155
rect 46102 19525 46154 19531
rect 46102 19467 46154 19473
rect 45238 18489 45290 18495
rect 45238 18431 45290 18437
rect 45238 14493 45290 14499
rect 45238 14435 45290 14441
rect 45250 7913 45278 14435
rect 46210 7913 46238 41149
rect 45238 7907 45290 7913
rect 45238 7849 45290 7855
rect 46198 7907 46250 7913
rect 46198 7849 46250 7855
rect 45250 7617 45278 7849
rect 45814 7759 45866 7765
rect 45814 7701 45866 7707
rect 45238 7611 45290 7617
rect 45238 7553 45290 7559
rect 45142 7167 45194 7173
rect 45142 7109 45194 7115
rect 45430 6945 45482 6951
rect 45346 6905 45430 6933
rect 45142 5687 45194 5693
rect 45142 5629 45194 5635
rect 45154 3103 45182 5629
rect 45238 3615 45290 3621
rect 45238 3557 45290 3563
rect 45142 3097 45194 3103
rect 45142 3039 45194 3045
rect 45142 2875 45194 2881
rect 45142 2817 45194 2823
rect 45154 800 45182 2817
rect 45250 800 45278 3557
rect 45346 3085 45374 6905
rect 45430 6887 45482 6893
rect 45526 6353 45578 6359
rect 45526 6295 45578 6301
rect 45430 5021 45482 5027
rect 45430 4963 45482 4969
rect 45442 3177 45470 4963
rect 45430 3171 45482 3177
rect 45430 3113 45482 3119
rect 45346 3057 45470 3085
rect 45442 800 45470 3057
rect 45538 800 45566 6295
rect 45622 3023 45674 3029
rect 45622 2965 45674 2971
rect 45634 800 45662 2965
rect 45826 800 45854 7701
rect 46210 7691 46238 7849
rect 46198 7685 46250 7691
rect 46198 7627 46250 7633
rect 46102 5687 46154 5693
rect 46102 5629 46154 5635
rect 46114 3640 46142 5629
rect 46306 5619 46334 42037
rect 46594 14943 46622 55357
rect 46786 52239 46814 56171
rect 46978 55717 47006 59200
rect 47554 56975 47582 59200
rect 47542 56969 47594 56975
rect 47542 56911 47594 56917
rect 48034 56531 48062 59200
rect 48022 56525 48074 56531
rect 48022 56467 48074 56473
rect 48214 56229 48266 56235
rect 48214 56171 48266 56177
rect 46966 55711 47018 55717
rect 46966 55653 47018 55659
rect 46774 52233 46826 52239
rect 46774 52175 46826 52181
rect 47830 48755 47882 48761
rect 47830 48697 47882 48703
rect 46966 23595 47018 23601
rect 46966 23537 47018 23543
rect 46678 22855 46730 22861
rect 46678 22797 46730 22803
rect 46582 14937 46634 14943
rect 46582 14879 46634 14885
rect 46486 7463 46538 7469
rect 46486 7405 46538 7411
rect 46294 5613 46346 5619
rect 46294 5555 46346 5561
rect 46198 5021 46250 5027
rect 46198 4963 46250 4969
rect 46294 5021 46346 5027
rect 46294 4963 46346 4969
rect 45922 3612 46142 3640
rect 45922 800 45950 3612
rect 46006 3541 46058 3547
rect 46006 3483 46058 3489
rect 46018 800 46046 3483
rect 46210 3251 46238 4963
rect 46198 3245 46250 3251
rect 46198 3187 46250 3193
rect 46306 3177 46334 4963
rect 46294 3171 46346 3177
rect 46294 3113 46346 3119
rect 46198 3097 46250 3103
rect 46198 3039 46250 3045
rect 46102 2505 46154 2511
rect 46102 2447 46154 2453
rect 46114 800 46142 2447
rect 46210 1420 46238 3039
rect 46294 2949 46346 2955
rect 46294 2891 46346 2897
rect 46306 1568 46334 2891
rect 46390 2801 46442 2807
rect 46390 2743 46442 2749
rect 46402 2585 46430 2743
rect 46390 2579 46442 2585
rect 46390 2521 46442 2527
rect 46306 1540 46430 1568
rect 46210 1392 46334 1420
rect 46306 800 46334 1392
rect 46402 800 46430 1540
rect 46498 800 46526 7405
rect 46690 7099 46718 22797
rect 46870 16935 46922 16941
rect 46870 16877 46922 16883
rect 46882 16571 46910 16877
rect 46870 16565 46922 16571
rect 46870 16507 46922 16513
rect 46978 9689 47006 23537
rect 47638 18785 47690 18791
rect 47638 18727 47690 18733
rect 47158 18341 47210 18347
rect 47158 18283 47210 18289
rect 46966 9683 47018 9689
rect 46966 9625 47018 9631
rect 47170 7765 47198 18283
rect 47542 12273 47594 12279
rect 47542 12215 47594 12221
rect 47554 7913 47582 12215
rect 47542 7907 47594 7913
rect 47542 7849 47594 7855
rect 47554 7765 47582 7849
rect 47158 7759 47210 7765
rect 47158 7701 47210 7707
rect 47542 7759 47594 7765
rect 47542 7701 47594 7707
rect 47254 7463 47306 7469
rect 47254 7405 47306 7411
rect 46678 7093 46730 7099
rect 46678 7035 46730 7041
rect 47062 6945 47114 6951
rect 47062 6887 47114 6893
rect 46870 6871 46922 6877
rect 46870 6813 46922 6819
rect 46678 5687 46730 5693
rect 46594 5647 46678 5675
rect 46594 800 46622 5647
rect 46678 5629 46730 5635
rect 46774 4355 46826 4361
rect 46774 4297 46826 4303
rect 46786 800 46814 4297
rect 46882 800 46910 6813
rect 46966 6353 47018 6359
rect 46966 6295 47018 6301
rect 46978 800 47006 6295
rect 47074 2511 47102 6887
rect 47158 3689 47210 3695
rect 47158 3631 47210 3637
rect 47062 2505 47114 2511
rect 47062 2447 47114 2453
rect 47170 800 47198 3631
rect 47266 800 47294 7405
rect 47650 7099 47678 18727
rect 47734 9461 47786 9467
rect 47734 9403 47786 9409
rect 47638 7093 47690 7099
rect 47638 7035 47690 7041
rect 47746 6507 47774 9403
rect 47842 7025 47870 48697
rect 48226 33591 48254 56171
rect 48610 56161 48638 59200
rect 49090 56901 49118 59200
rect 49078 56895 49130 56901
rect 49078 56837 49130 56843
rect 48694 56747 48746 56753
rect 48694 56689 48746 56695
rect 48598 56155 48650 56161
rect 48598 56097 48650 56103
rect 48598 51493 48650 51499
rect 48598 51435 48650 51441
rect 48214 33585 48266 33591
rect 48214 33527 48266 33533
rect 48118 27887 48170 27893
rect 48118 27829 48170 27835
rect 48130 8431 48158 27829
rect 48310 13235 48362 13241
rect 48310 13177 48362 13183
rect 48118 8425 48170 8431
rect 48118 8367 48170 8373
rect 48022 8203 48074 8209
rect 48022 8145 48074 8151
rect 47830 7019 47882 7025
rect 47830 6961 47882 6967
rect 47734 6501 47786 6507
rect 47734 6443 47786 6449
rect 47734 6353 47786 6359
rect 47734 6295 47786 6301
rect 47542 5687 47594 5693
rect 47542 5629 47594 5635
rect 47554 4380 47582 5629
rect 47638 5021 47690 5027
rect 47638 4963 47690 4969
rect 47362 4352 47582 4380
rect 47362 800 47390 4352
rect 47446 4281 47498 4287
rect 47446 4223 47498 4229
rect 47458 800 47486 4223
rect 47650 3103 47678 4963
rect 47638 3097 47690 3103
rect 47638 3039 47690 3045
rect 47638 2949 47690 2955
rect 47638 2891 47690 2897
rect 47650 800 47678 2891
rect 47746 800 47774 6295
rect 47830 4355 47882 4361
rect 47830 4297 47882 4303
rect 47842 800 47870 4297
rect 48034 800 48062 8145
rect 48322 7099 48350 13177
rect 48610 8579 48638 51435
rect 48706 21603 48734 56689
rect 49666 56531 49694 59200
rect 50146 56531 50174 59200
rect 50722 56901 50750 59200
rect 50710 56895 50762 56901
rect 50710 56837 50762 56843
rect 50806 56747 50858 56753
rect 50806 56689 50858 56695
rect 50348 56638 50644 56658
rect 50404 56636 50428 56638
rect 50484 56636 50508 56638
rect 50564 56636 50588 56638
rect 50426 56584 50428 56636
rect 50490 56584 50502 56636
rect 50564 56584 50566 56636
rect 50404 56582 50428 56584
rect 50484 56582 50508 56584
rect 50564 56582 50588 56584
rect 50348 56562 50644 56582
rect 49654 56525 49706 56531
rect 49654 56467 49706 56473
rect 50134 56525 50186 56531
rect 50134 56467 50186 56473
rect 48790 56229 48842 56235
rect 48790 56171 48842 56177
rect 49942 56229 49994 56235
rect 49942 56171 49994 56177
rect 48694 21597 48746 21603
rect 48694 21539 48746 21545
rect 48802 19901 48830 56171
rect 48886 52899 48938 52905
rect 48886 52841 48938 52847
rect 48790 19895 48842 19901
rect 48790 19837 48842 19843
rect 48598 8573 48650 8579
rect 48598 8515 48650 8521
rect 48694 8277 48746 8283
rect 48694 8219 48746 8225
rect 48406 7759 48458 7765
rect 48406 7701 48458 7707
rect 48310 7093 48362 7099
rect 48310 7035 48362 7041
rect 48214 3689 48266 3695
rect 48418 3640 48446 7701
rect 48598 4281 48650 4287
rect 48598 4223 48650 4229
rect 48214 3631 48266 3637
rect 48118 3171 48170 3177
rect 48118 3113 48170 3119
rect 48130 800 48158 3113
rect 48226 800 48254 3631
rect 48322 3612 48446 3640
rect 48322 800 48350 3612
rect 48502 3245 48554 3251
rect 48502 3187 48554 3193
rect 48514 800 48542 3187
rect 48610 800 48638 4223
rect 48706 800 48734 8219
rect 48898 7173 48926 52841
rect 49174 50235 49226 50241
rect 49174 50177 49226 50183
rect 49186 50093 49214 50177
rect 49174 50087 49226 50093
rect 49174 50029 49226 50035
rect 48982 49051 49034 49057
rect 48982 48993 49034 48999
rect 48994 7913 49022 48993
rect 49186 9837 49214 50029
rect 49954 47534 49982 56171
rect 50348 55306 50644 55326
rect 50404 55304 50428 55306
rect 50484 55304 50508 55306
rect 50564 55304 50588 55306
rect 50426 55252 50428 55304
rect 50490 55252 50502 55304
rect 50564 55252 50566 55304
rect 50404 55250 50428 55252
rect 50484 55250 50508 55252
rect 50564 55250 50588 55252
rect 50348 55230 50644 55250
rect 50348 53974 50644 53994
rect 50404 53972 50428 53974
rect 50484 53972 50508 53974
rect 50564 53972 50588 53974
rect 50426 53920 50428 53972
rect 50490 53920 50502 53972
rect 50564 53920 50566 53972
rect 50404 53918 50428 53920
rect 50484 53918 50508 53920
rect 50564 53918 50588 53920
rect 50348 53898 50644 53918
rect 50348 52642 50644 52662
rect 50404 52640 50428 52642
rect 50484 52640 50508 52642
rect 50564 52640 50588 52642
rect 50426 52588 50428 52640
rect 50490 52588 50502 52640
rect 50564 52588 50566 52640
rect 50404 52586 50428 52588
rect 50484 52586 50508 52588
rect 50564 52586 50588 52588
rect 50348 52566 50644 52586
rect 50348 51310 50644 51330
rect 50404 51308 50428 51310
rect 50484 51308 50508 51310
rect 50564 51308 50588 51310
rect 50426 51256 50428 51308
rect 50490 51256 50502 51308
rect 50564 51256 50566 51308
rect 50404 51254 50428 51256
rect 50484 51254 50508 51256
rect 50564 51254 50588 51256
rect 50348 51234 50644 51254
rect 50348 49978 50644 49998
rect 50404 49976 50428 49978
rect 50484 49976 50508 49978
rect 50564 49976 50588 49978
rect 50426 49924 50428 49976
rect 50490 49924 50502 49976
rect 50564 49924 50566 49976
rect 50404 49922 50428 49924
rect 50484 49922 50508 49924
rect 50564 49922 50588 49924
rect 50348 49902 50644 49922
rect 50348 48646 50644 48666
rect 50404 48644 50428 48646
rect 50484 48644 50508 48646
rect 50564 48644 50588 48646
rect 50426 48592 50428 48644
rect 50490 48592 50502 48644
rect 50564 48592 50566 48644
rect 50404 48590 50428 48592
rect 50484 48590 50508 48592
rect 50564 48590 50588 48592
rect 50348 48570 50644 48590
rect 49666 47506 49982 47534
rect 49666 33221 49694 47506
rect 50348 47314 50644 47334
rect 50404 47312 50428 47314
rect 50484 47312 50508 47314
rect 50564 47312 50588 47314
rect 50426 47260 50428 47312
rect 50490 47260 50502 47312
rect 50564 47260 50566 47312
rect 50404 47258 50428 47260
rect 50484 47258 50508 47260
rect 50564 47258 50588 47260
rect 50348 47238 50644 47258
rect 50348 45982 50644 46002
rect 50404 45980 50428 45982
rect 50484 45980 50508 45982
rect 50564 45980 50588 45982
rect 50426 45928 50428 45980
rect 50490 45928 50502 45980
rect 50564 45928 50566 45980
rect 50404 45926 50428 45928
rect 50484 45926 50508 45928
rect 50564 45926 50588 45928
rect 50348 45906 50644 45926
rect 50348 44650 50644 44670
rect 50404 44648 50428 44650
rect 50484 44648 50508 44650
rect 50564 44648 50588 44650
rect 50426 44596 50428 44648
rect 50490 44596 50502 44648
rect 50564 44596 50566 44648
rect 50404 44594 50428 44596
rect 50484 44594 50508 44596
rect 50564 44594 50588 44596
rect 50348 44574 50644 44594
rect 50348 43318 50644 43338
rect 50404 43316 50428 43318
rect 50484 43316 50508 43318
rect 50564 43316 50588 43318
rect 50426 43264 50428 43316
rect 50490 43264 50502 43316
rect 50564 43264 50566 43316
rect 50404 43262 50428 43264
rect 50484 43262 50508 43264
rect 50564 43262 50588 43264
rect 50348 43242 50644 43262
rect 50348 41986 50644 42006
rect 50404 41984 50428 41986
rect 50484 41984 50508 41986
rect 50564 41984 50588 41986
rect 50426 41932 50428 41984
rect 50490 41932 50502 41984
rect 50564 41932 50566 41984
rect 50404 41930 50428 41932
rect 50484 41930 50508 41932
rect 50564 41930 50588 41932
rect 50348 41910 50644 41930
rect 50348 40654 50644 40674
rect 50404 40652 50428 40654
rect 50484 40652 50508 40654
rect 50564 40652 50588 40654
rect 50426 40600 50428 40652
rect 50490 40600 50502 40652
rect 50564 40600 50566 40652
rect 50404 40598 50428 40600
rect 50484 40598 50508 40600
rect 50564 40598 50588 40600
rect 50348 40578 50644 40598
rect 50348 39322 50644 39342
rect 50404 39320 50428 39322
rect 50484 39320 50508 39322
rect 50564 39320 50588 39322
rect 50426 39268 50428 39320
rect 50490 39268 50502 39320
rect 50564 39268 50566 39320
rect 50404 39266 50428 39268
rect 50484 39266 50508 39268
rect 50564 39266 50588 39268
rect 50348 39246 50644 39266
rect 50230 38247 50282 38253
rect 50230 38189 50282 38195
rect 49654 33215 49706 33221
rect 49654 33157 49706 33163
rect 49750 23447 49802 23453
rect 49750 23389 49802 23395
rect 49174 9831 49226 9837
rect 49174 9773 49226 9779
rect 49762 8431 49790 23389
rect 49846 19229 49898 19235
rect 49846 19171 49898 19177
rect 49750 8425 49802 8431
rect 49750 8367 49802 8373
rect 49462 8277 49514 8283
rect 49462 8219 49514 8225
rect 48982 7907 49034 7913
rect 48982 7849 49034 7855
rect 48994 7691 49022 7849
rect 48982 7685 49034 7691
rect 48982 7627 49034 7633
rect 49078 7537 49130 7543
rect 49078 7479 49130 7485
rect 48886 7167 48938 7173
rect 48886 7109 48938 7115
rect 48886 6945 48938 6951
rect 48886 6887 48938 6893
rect 48790 6353 48842 6359
rect 48790 6295 48842 6301
rect 48802 800 48830 6295
rect 48898 2955 48926 6887
rect 48982 5687 49034 5693
rect 48982 5629 49034 5635
rect 48994 3177 49022 5629
rect 48982 3171 49034 3177
rect 48982 3113 49034 3119
rect 48886 2949 48938 2955
rect 48886 2891 48938 2897
rect 48982 2949 49034 2955
rect 48982 2891 49034 2897
rect 48994 800 49022 2891
rect 49090 800 49118 7479
rect 49270 5909 49322 5915
rect 49270 5851 49322 5857
rect 49174 3837 49226 3843
rect 49174 3779 49226 3785
rect 49186 800 49214 3779
rect 49282 2437 49310 5851
rect 49366 5021 49418 5027
rect 49366 4963 49418 4969
rect 49270 2431 49322 2437
rect 49270 2373 49322 2379
rect 49378 800 49406 4963
rect 49474 800 49502 8219
rect 49654 7685 49706 7691
rect 49654 7627 49706 7633
rect 49558 6353 49610 6359
rect 49558 6295 49610 6301
rect 49570 800 49598 6295
rect 49666 5915 49694 7627
rect 49858 7173 49886 19171
rect 49846 7167 49898 7173
rect 49846 7109 49898 7115
rect 50242 7099 50270 38189
rect 50348 37990 50644 38010
rect 50404 37988 50428 37990
rect 50484 37988 50508 37990
rect 50564 37988 50588 37990
rect 50426 37936 50428 37988
rect 50490 37936 50502 37988
rect 50564 37936 50566 37988
rect 50404 37934 50428 37936
rect 50484 37934 50508 37936
rect 50564 37934 50588 37936
rect 50348 37914 50644 37934
rect 50348 36658 50644 36678
rect 50404 36656 50428 36658
rect 50484 36656 50508 36658
rect 50564 36656 50588 36658
rect 50426 36604 50428 36656
rect 50490 36604 50502 36656
rect 50564 36604 50566 36656
rect 50404 36602 50428 36604
rect 50484 36602 50508 36604
rect 50564 36602 50588 36604
rect 50348 36582 50644 36602
rect 50348 35326 50644 35346
rect 50404 35324 50428 35326
rect 50484 35324 50508 35326
rect 50564 35324 50588 35326
rect 50426 35272 50428 35324
rect 50490 35272 50502 35324
rect 50564 35272 50566 35324
rect 50404 35270 50428 35272
rect 50484 35270 50508 35272
rect 50564 35270 50588 35272
rect 50348 35250 50644 35270
rect 50348 33994 50644 34014
rect 50404 33992 50428 33994
rect 50484 33992 50508 33994
rect 50564 33992 50588 33994
rect 50426 33940 50428 33992
rect 50490 33940 50502 33992
rect 50564 33940 50566 33992
rect 50404 33938 50428 33940
rect 50484 33938 50508 33940
rect 50564 33938 50588 33940
rect 50348 33918 50644 33938
rect 50348 32662 50644 32682
rect 50404 32660 50428 32662
rect 50484 32660 50508 32662
rect 50564 32660 50588 32662
rect 50426 32608 50428 32660
rect 50490 32608 50502 32660
rect 50564 32608 50566 32660
rect 50404 32606 50428 32608
rect 50484 32606 50508 32608
rect 50564 32606 50588 32608
rect 50348 32586 50644 32606
rect 50348 31330 50644 31350
rect 50404 31328 50428 31330
rect 50484 31328 50508 31330
rect 50564 31328 50588 31330
rect 50426 31276 50428 31328
rect 50490 31276 50502 31328
rect 50564 31276 50566 31328
rect 50404 31274 50428 31276
rect 50484 31274 50508 31276
rect 50564 31274 50588 31276
rect 50348 31254 50644 31274
rect 50348 29998 50644 30018
rect 50404 29996 50428 29998
rect 50484 29996 50508 29998
rect 50564 29996 50588 29998
rect 50426 29944 50428 29996
rect 50490 29944 50502 29996
rect 50564 29944 50566 29996
rect 50404 29942 50428 29944
rect 50484 29942 50508 29944
rect 50564 29942 50588 29944
rect 50348 29922 50644 29942
rect 50348 28666 50644 28686
rect 50404 28664 50428 28666
rect 50484 28664 50508 28666
rect 50564 28664 50588 28666
rect 50426 28612 50428 28664
rect 50490 28612 50502 28664
rect 50564 28612 50566 28664
rect 50404 28610 50428 28612
rect 50484 28610 50508 28612
rect 50564 28610 50588 28612
rect 50348 28590 50644 28610
rect 50348 27334 50644 27354
rect 50404 27332 50428 27334
rect 50484 27332 50508 27334
rect 50564 27332 50588 27334
rect 50426 27280 50428 27332
rect 50490 27280 50502 27332
rect 50564 27280 50566 27332
rect 50404 27278 50428 27280
rect 50484 27278 50508 27280
rect 50564 27278 50588 27280
rect 50348 27258 50644 27278
rect 50348 26002 50644 26022
rect 50404 26000 50428 26002
rect 50484 26000 50508 26002
rect 50564 26000 50588 26002
rect 50426 25948 50428 26000
rect 50490 25948 50502 26000
rect 50564 25948 50566 26000
rect 50404 25946 50428 25948
rect 50484 25946 50508 25948
rect 50564 25946 50588 25948
rect 50348 25926 50644 25946
rect 50348 24670 50644 24690
rect 50404 24668 50428 24670
rect 50484 24668 50508 24670
rect 50564 24668 50588 24670
rect 50426 24616 50428 24668
rect 50490 24616 50502 24668
rect 50564 24616 50566 24668
rect 50404 24614 50428 24616
rect 50484 24614 50508 24616
rect 50564 24614 50588 24616
rect 50348 24594 50644 24614
rect 50348 23338 50644 23358
rect 50404 23336 50428 23338
rect 50484 23336 50508 23338
rect 50564 23336 50588 23338
rect 50426 23284 50428 23336
rect 50490 23284 50502 23336
rect 50564 23284 50566 23336
rect 50404 23282 50428 23284
rect 50484 23282 50508 23284
rect 50564 23282 50588 23284
rect 50348 23262 50644 23282
rect 50348 22006 50644 22026
rect 50404 22004 50428 22006
rect 50484 22004 50508 22006
rect 50564 22004 50588 22006
rect 50426 21952 50428 22004
rect 50490 21952 50502 22004
rect 50564 21952 50566 22004
rect 50404 21950 50428 21952
rect 50484 21950 50508 21952
rect 50564 21950 50588 21952
rect 50348 21930 50644 21950
rect 50818 20937 50846 56689
rect 51202 56161 51230 59200
rect 51670 56229 51722 56235
rect 51670 56171 51722 56177
rect 51190 56155 51242 56161
rect 51190 56097 51242 56103
rect 51574 55415 51626 55421
rect 51574 55357 51626 55363
rect 51286 49421 51338 49427
rect 51286 49363 51338 49369
rect 51190 24927 51242 24933
rect 51190 24869 51242 24875
rect 50806 20931 50858 20937
rect 50806 20873 50858 20879
rect 50348 20674 50644 20694
rect 50404 20672 50428 20674
rect 50484 20672 50508 20674
rect 50564 20672 50588 20674
rect 50426 20620 50428 20672
rect 50490 20620 50502 20672
rect 50564 20620 50566 20672
rect 50404 20618 50428 20620
rect 50484 20618 50508 20620
rect 50564 20618 50588 20620
rect 50348 20598 50644 20618
rect 50348 19342 50644 19362
rect 50404 19340 50428 19342
rect 50484 19340 50508 19342
rect 50564 19340 50588 19342
rect 50426 19288 50428 19340
rect 50490 19288 50502 19340
rect 50564 19288 50566 19340
rect 50404 19286 50428 19288
rect 50484 19286 50508 19288
rect 50564 19286 50588 19288
rect 50348 19266 50644 19286
rect 50998 18119 51050 18125
rect 50998 18061 51050 18067
rect 50348 18010 50644 18030
rect 50404 18008 50428 18010
rect 50484 18008 50508 18010
rect 50564 18008 50588 18010
rect 50426 17956 50428 18008
rect 50490 17956 50502 18008
rect 50564 17956 50566 18008
rect 50404 17954 50428 17956
rect 50484 17954 50508 17956
rect 50564 17954 50588 17956
rect 50348 17934 50644 17954
rect 51010 17829 51038 18061
rect 50998 17823 51050 17829
rect 50998 17765 51050 17771
rect 50348 16678 50644 16698
rect 50404 16676 50428 16678
rect 50484 16676 50508 16678
rect 50564 16676 50588 16678
rect 50426 16624 50428 16676
rect 50490 16624 50502 16676
rect 50564 16624 50566 16676
rect 50404 16622 50428 16624
rect 50484 16622 50508 16624
rect 50564 16622 50588 16624
rect 50348 16602 50644 16622
rect 50348 15346 50644 15366
rect 50404 15344 50428 15346
rect 50484 15344 50508 15346
rect 50564 15344 50588 15346
rect 50426 15292 50428 15344
rect 50490 15292 50502 15344
rect 50564 15292 50566 15344
rect 50404 15290 50428 15292
rect 50484 15290 50508 15292
rect 50564 15290 50588 15292
rect 50348 15270 50644 15290
rect 50348 14014 50644 14034
rect 50404 14012 50428 14014
rect 50484 14012 50508 14014
rect 50564 14012 50588 14014
rect 50426 13960 50428 14012
rect 50490 13960 50502 14012
rect 50564 13960 50566 14012
rect 50404 13958 50428 13960
rect 50484 13958 50508 13960
rect 50564 13958 50588 13960
rect 50348 13938 50644 13958
rect 50348 12682 50644 12702
rect 50404 12680 50428 12682
rect 50484 12680 50508 12682
rect 50564 12680 50588 12682
rect 50426 12628 50428 12680
rect 50490 12628 50502 12680
rect 50564 12628 50566 12680
rect 50404 12626 50428 12628
rect 50484 12626 50508 12628
rect 50564 12626 50588 12628
rect 50348 12606 50644 12626
rect 50348 11350 50644 11370
rect 50404 11348 50428 11350
rect 50484 11348 50508 11350
rect 50564 11348 50588 11350
rect 50426 11296 50428 11348
rect 50490 11296 50502 11348
rect 50564 11296 50566 11348
rect 50404 11294 50428 11296
rect 50484 11294 50508 11296
rect 50564 11294 50588 11296
rect 50348 11274 50644 11294
rect 50902 10793 50954 10799
rect 50902 10735 50954 10741
rect 50348 10018 50644 10038
rect 50404 10016 50428 10018
rect 50484 10016 50508 10018
rect 50564 10016 50588 10018
rect 50426 9964 50428 10016
rect 50490 9964 50502 10016
rect 50564 9964 50566 10016
rect 50404 9962 50428 9964
rect 50484 9962 50508 9964
rect 50564 9962 50588 9964
rect 50348 9942 50644 9962
rect 50348 8686 50644 8706
rect 50404 8684 50428 8686
rect 50484 8684 50508 8686
rect 50564 8684 50588 8686
rect 50426 8632 50428 8684
rect 50490 8632 50502 8684
rect 50564 8632 50566 8684
rect 50404 8630 50428 8632
rect 50484 8630 50508 8632
rect 50564 8630 50588 8632
rect 50348 8610 50644 8630
rect 50348 7354 50644 7374
rect 50404 7352 50428 7354
rect 50484 7352 50508 7354
rect 50564 7352 50588 7354
rect 50426 7300 50428 7352
rect 50490 7300 50502 7352
rect 50564 7300 50566 7352
rect 50404 7298 50428 7300
rect 50484 7298 50508 7300
rect 50564 7298 50588 7300
rect 50348 7278 50644 7298
rect 50230 7093 50282 7099
rect 50230 7035 50282 7041
rect 50134 6945 50186 6951
rect 50134 6887 50186 6893
rect 49750 6131 49802 6137
rect 49750 6073 49802 6079
rect 49654 5909 49706 5915
rect 49654 5851 49706 5857
rect 49654 5687 49706 5693
rect 49654 5629 49706 5635
rect 49666 3251 49694 5629
rect 49654 3245 49706 3251
rect 49654 3187 49706 3193
rect 49654 3023 49706 3029
rect 49654 2965 49706 2971
rect 49666 800 49694 2965
rect 49762 2012 49790 6073
rect 49846 4355 49898 4361
rect 49846 4297 49898 4303
rect 49858 2955 49886 4297
rect 49942 4281 49994 4287
rect 49942 4223 49994 4229
rect 49846 2949 49898 2955
rect 49846 2891 49898 2897
rect 49762 1984 49886 2012
rect 49858 800 49886 1984
rect 49954 800 49982 4223
rect 50038 2875 50090 2881
rect 50038 2817 50090 2823
rect 50050 800 50078 2817
rect 50146 800 50174 6887
rect 50914 6433 50942 10735
rect 51202 8357 51230 24869
rect 51190 8351 51242 8357
rect 51190 8293 51242 8299
rect 51298 6581 51326 49363
rect 51586 13759 51614 55357
rect 51682 18347 51710 56171
rect 51778 55717 51806 59200
rect 52258 56901 52286 59200
rect 52246 56895 52298 56901
rect 52834 56883 52862 59200
rect 52834 56855 52958 56883
rect 52246 56837 52298 56843
rect 52822 56747 52874 56753
rect 52822 56689 52874 56695
rect 51766 55711 51818 55717
rect 51766 55653 51818 55659
rect 52630 55637 52682 55643
rect 52630 55579 52682 55585
rect 52054 49421 52106 49427
rect 52054 49363 52106 49369
rect 52066 49131 52094 49363
rect 52054 49125 52106 49131
rect 52054 49067 52106 49073
rect 52342 38765 52394 38771
rect 52342 38707 52394 38713
rect 52354 38475 52382 38707
rect 52342 38469 52394 38475
rect 52342 38411 52394 38417
rect 51766 36915 51818 36921
rect 51766 36857 51818 36863
rect 51670 18341 51722 18347
rect 51670 18283 51722 18289
rect 51574 13753 51626 13759
rect 51574 13695 51626 13701
rect 51574 10275 51626 10281
rect 51574 10217 51626 10223
rect 51586 8431 51614 10217
rect 51670 9831 51722 9837
rect 51670 9773 51722 9779
rect 51682 9245 51710 9773
rect 51670 9239 51722 9245
rect 51670 9181 51722 9187
rect 51574 8425 51626 8431
rect 51574 8367 51626 8373
rect 51778 7765 51806 36857
rect 52054 31883 52106 31889
rect 52054 31825 52106 31831
rect 51766 7759 51818 7765
rect 51766 7701 51818 7707
rect 51670 7463 51722 7469
rect 51670 7405 51722 7411
rect 51382 6945 51434 6951
rect 51382 6887 51434 6893
rect 51286 6575 51338 6581
rect 51286 6517 51338 6523
rect 50902 6427 50954 6433
rect 50902 6369 50954 6375
rect 51094 6131 51146 6137
rect 51094 6073 51146 6079
rect 50348 6022 50644 6042
rect 50404 6020 50428 6022
rect 50484 6020 50508 6022
rect 50564 6020 50588 6022
rect 50426 5968 50428 6020
rect 50490 5968 50502 6020
rect 50564 5968 50566 6020
rect 50404 5966 50428 5968
rect 50484 5966 50508 5968
rect 50564 5966 50588 5968
rect 50348 5946 50644 5966
rect 50710 5687 50762 5693
rect 50710 5629 50762 5635
rect 50422 5021 50474 5027
rect 50422 4963 50474 4969
rect 50434 4824 50462 4963
rect 50242 4796 50462 4824
rect 50242 2604 50270 4796
rect 50348 4690 50644 4710
rect 50404 4688 50428 4690
rect 50484 4688 50508 4690
rect 50564 4688 50588 4690
rect 50426 4636 50428 4688
rect 50490 4636 50502 4688
rect 50564 4636 50566 4688
rect 50404 4634 50428 4636
rect 50484 4634 50508 4636
rect 50564 4634 50588 4636
rect 50348 4614 50644 4634
rect 50722 3843 50750 5629
rect 50902 5021 50954 5027
rect 50902 4963 50954 4969
rect 50710 3837 50762 3843
rect 50710 3779 50762 3785
rect 50710 3689 50762 3695
rect 50710 3631 50762 3637
rect 50806 3689 50858 3695
rect 50806 3631 50858 3637
rect 50348 3358 50644 3378
rect 50404 3356 50428 3358
rect 50484 3356 50508 3358
rect 50564 3356 50588 3358
rect 50426 3304 50428 3356
rect 50490 3304 50502 3356
rect 50564 3304 50566 3356
rect 50404 3302 50428 3304
rect 50484 3302 50508 3304
rect 50564 3302 50588 3304
rect 50348 3282 50644 3302
rect 50242 2576 50366 2604
rect 50338 800 50366 2576
rect 50722 1864 50750 3631
rect 50434 1836 50750 1864
rect 50434 800 50462 1836
rect 50518 1765 50570 1771
rect 50518 1707 50570 1713
rect 50530 800 50558 1707
rect 50710 1617 50762 1623
rect 50710 1559 50762 1565
rect 50722 800 50750 1559
rect 50818 800 50846 3631
rect 50914 1623 50942 4963
rect 50998 4281 51050 4287
rect 50998 4223 51050 4229
rect 50902 1617 50954 1623
rect 50902 1559 50954 1565
rect 50902 1469 50954 1475
rect 50902 1411 50954 1417
rect 50914 800 50942 1411
rect 51010 800 51038 4223
rect 51106 1771 51134 6073
rect 51286 3689 51338 3695
rect 51202 3649 51286 3677
rect 51094 1765 51146 1771
rect 51094 1707 51146 1713
rect 51202 800 51230 3649
rect 51286 3631 51338 3637
rect 51394 3492 51422 6887
rect 51574 6205 51626 6211
rect 51574 6147 51626 6153
rect 51298 3464 51422 3492
rect 51298 800 51326 3464
rect 51478 3023 51530 3029
rect 51478 2965 51530 2971
rect 51382 2949 51434 2955
rect 51382 2891 51434 2897
rect 51394 800 51422 2891
rect 51490 800 51518 2965
rect 51586 1475 51614 6147
rect 51574 1469 51626 1475
rect 51574 1411 51626 1417
rect 51682 800 51710 7405
rect 52066 7099 52094 31825
rect 52438 16121 52490 16127
rect 52438 16063 52490 16069
rect 52342 7463 52394 7469
rect 52342 7405 52394 7411
rect 52054 7093 52106 7099
rect 52054 7035 52106 7041
rect 52150 5687 52202 5693
rect 52150 5629 52202 5635
rect 51862 5021 51914 5027
rect 51862 4963 51914 4969
rect 51766 3097 51818 3103
rect 51766 3039 51818 3045
rect 51778 800 51806 3039
rect 51874 2955 51902 4963
rect 52054 3689 52106 3695
rect 51970 3649 52054 3677
rect 51862 2949 51914 2955
rect 51862 2891 51914 2897
rect 51970 1864 51998 3649
rect 52054 3631 52106 3637
rect 52054 3541 52106 3547
rect 52054 3483 52106 3489
rect 51874 1836 51998 1864
rect 51874 800 51902 1836
rect 52066 800 52094 3483
rect 52162 800 52190 5629
rect 52246 5021 52298 5027
rect 52246 4963 52298 4969
rect 52258 3103 52286 4963
rect 52246 3097 52298 3103
rect 52246 3039 52298 3045
rect 52246 2949 52298 2955
rect 52246 2891 52298 2897
rect 52258 800 52286 2891
rect 52354 800 52382 7405
rect 52450 6433 52478 16063
rect 52534 11607 52586 11613
rect 52534 11549 52586 11555
rect 52438 6427 52490 6433
rect 52438 6369 52490 6375
rect 52546 5860 52574 11549
rect 52642 7765 52670 55579
rect 52834 21529 52862 56689
rect 52930 56531 52958 56855
rect 53314 56531 53342 59200
rect 53890 56975 53918 59200
rect 53878 56969 53930 56975
rect 53878 56911 53930 56917
rect 54370 56531 54398 59200
rect 54946 56531 54974 59200
rect 55426 56901 55454 59200
rect 55414 56895 55466 56901
rect 55414 56837 55466 56843
rect 55414 56747 55466 56753
rect 55414 56689 55466 56695
rect 52918 56525 52970 56531
rect 52918 56467 52970 56473
rect 53302 56525 53354 56531
rect 53302 56467 53354 56473
rect 54358 56525 54410 56531
rect 54358 56467 54410 56473
rect 54934 56525 54986 56531
rect 54934 56467 54986 56473
rect 53686 56229 53738 56235
rect 53686 56171 53738 56177
rect 54550 56229 54602 56235
rect 54550 56171 54602 56177
rect 53014 54231 53066 54237
rect 53014 54173 53066 54179
rect 52918 51567 52970 51573
rect 52918 51509 52970 51515
rect 52822 21523 52874 21529
rect 52822 21465 52874 21471
rect 52930 7913 52958 51509
rect 53026 9245 53054 54173
rect 53206 45203 53258 45209
rect 53206 45145 53258 45151
rect 53014 9239 53066 9245
rect 53014 9181 53066 9187
rect 53218 8431 53246 45145
rect 53698 32185 53726 56171
rect 54262 47571 54314 47577
rect 54262 47513 54314 47519
rect 53686 32179 53738 32185
rect 53686 32121 53738 32127
rect 54274 17294 54302 47513
rect 54562 31075 54590 56171
rect 54550 31069 54602 31075
rect 54550 31011 54602 31017
rect 55426 22935 55454 56689
rect 56002 56531 56030 59200
rect 55990 56525 56042 56531
rect 55990 56467 56042 56473
rect 55510 56229 55562 56235
rect 55510 56171 55562 56177
rect 55414 22929 55466 22935
rect 55414 22871 55466 22877
rect 55522 20789 55550 56171
rect 56482 55717 56510 59200
rect 57058 56901 57086 59200
rect 57046 56895 57098 56901
rect 57046 56837 57098 56843
rect 56758 56747 56810 56753
rect 56758 56689 56810 56695
rect 56770 56457 56798 56689
rect 56758 56451 56810 56457
rect 56758 56393 56810 56399
rect 57538 55717 57566 59200
rect 56470 55711 56522 55717
rect 56470 55653 56522 55659
rect 57526 55711 57578 55717
rect 57526 55653 57578 55659
rect 55606 55415 55658 55421
rect 55606 55357 55658 55363
rect 56278 55415 56330 55421
rect 56278 55357 56330 55363
rect 57334 55415 57386 55421
rect 57334 55357 57386 55363
rect 55618 55199 55646 55357
rect 55606 55193 55658 55199
rect 55606 55135 55658 55141
rect 55798 54749 55850 54755
rect 55798 54691 55850 54697
rect 55810 54163 55838 54691
rect 55798 54157 55850 54163
rect 55798 54099 55850 54105
rect 55606 48977 55658 48983
rect 55606 48919 55658 48925
rect 55510 20783 55562 20789
rect 55510 20725 55562 20731
rect 54178 17266 54302 17294
rect 54070 16491 54122 16497
rect 54070 16433 54122 16439
rect 53878 8795 53930 8801
rect 53878 8737 53930 8743
rect 53206 8425 53258 8431
rect 53206 8367 53258 8373
rect 53494 8277 53546 8283
rect 53494 8219 53546 8225
rect 53110 8203 53162 8209
rect 53110 8145 53162 8151
rect 52918 7907 52970 7913
rect 52918 7849 52970 7855
rect 52630 7759 52682 7765
rect 52630 7701 52682 7707
rect 52726 7759 52778 7765
rect 52726 7701 52778 7707
rect 52450 5832 52574 5860
rect 52450 2807 52478 5832
rect 52534 5687 52586 5693
rect 52534 5629 52586 5635
rect 52438 2801 52490 2807
rect 52438 2743 52490 2749
rect 52546 800 52574 5629
rect 52630 4355 52682 4361
rect 52630 4297 52682 4303
rect 52642 800 52670 4297
rect 52738 800 52766 7701
rect 52930 7691 52958 7849
rect 52918 7685 52970 7691
rect 52918 7627 52970 7633
rect 52822 6945 52874 6951
rect 52822 6887 52874 6893
rect 52834 3547 52862 6887
rect 53014 4281 53066 4287
rect 53014 4223 53066 4229
rect 52822 3541 52874 3547
rect 52822 3483 52874 3489
rect 52918 2949 52970 2955
rect 52918 2891 52970 2897
rect 52930 800 52958 2891
rect 53026 800 53054 4223
rect 53122 800 53150 8145
rect 53302 5021 53354 5027
rect 53302 4963 53354 4969
rect 53314 2900 53342 4963
rect 53398 3689 53450 3695
rect 53398 3631 53450 3637
rect 53218 2872 53342 2900
rect 53218 800 53246 2872
rect 53410 800 53438 3631
rect 53506 800 53534 8219
rect 53686 5687 53738 5693
rect 53686 5629 53738 5635
rect 53590 5613 53642 5619
rect 53590 5555 53642 5561
rect 53602 800 53630 5555
rect 53698 2955 53726 5629
rect 53782 3023 53834 3029
rect 53782 2965 53834 2971
rect 53686 2949 53738 2955
rect 53686 2891 53738 2897
rect 53794 1568 53822 2965
rect 53698 1540 53822 1568
rect 53698 800 53726 1540
rect 53890 800 53918 8737
rect 54082 8431 54110 16433
rect 54070 8425 54122 8431
rect 54070 8367 54122 8373
rect 54178 7839 54206 17266
rect 54646 11607 54698 11613
rect 54646 11549 54698 11555
rect 54658 9763 54686 11549
rect 55126 9905 55178 9911
rect 55126 9847 55178 9853
rect 54646 9757 54698 9763
rect 54646 9699 54698 9705
rect 54262 9609 54314 9615
rect 54262 9551 54314 9557
rect 54934 9609 54986 9615
rect 54934 9551 54986 9557
rect 54166 7833 54218 7839
rect 54166 7775 54218 7781
rect 53974 6353 54026 6359
rect 53974 6295 54026 6301
rect 53986 800 54014 6295
rect 54070 4355 54122 4361
rect 54070 4297 54122 4303
rect 54082 800 54110 4297
rect 54274 800 54302 9551
rect 54550 9091 54602 9097
rect 54550 9033 54602 9039
rect 54358 6279 54410 6285
rect 54358 6221 54410 6227
rect 54370 800 54398 6221
rect 54454 3541 54506 3547
rect 54454 3483 54506 3489
rect 54466 800 54494 3483
rect 54562 800 54590 9033
rect 54742 7019 54794 7025
rect 54742 6961 54794 6967
rect 54754 800 54782 6961
rect 54838 2949 54890 2955
rect 54838 2891 54890 2897
rect 54850 800 54878 2891
rect 54946 800 54974 9551
rect 55030 6205 55082 6211
rect 55030 6147 55082 6153
rect 55042 800 55070 6147
rect 55138 3640 55166 9847
rect 55618 9245 55646 48919
rect 55990 38543 56042 38549
rect 55990 38485 56042 38491
rect 56002 17294 56030 38485
rect 56290 36107 56318 55357
rect 56854 50309 56906 50315
rect 56854 50251 56906 50257
rect 56278 36101 56330 36107
rect 56278 36043 56330 36049
rect 56002 17266 56126 17294
rect 55990 16935 56042 16941
rect 55990 16877 56042 16883
rect 56002 10429 56030 16877
rect 56098 11095 56126 17266
rect 56086 11089 56138 11095
rect 56086 11031 56138 11037
rect 56758 10941 56810 10947
rect 56758 10883 56810 10889
rect 55990 10423 56042 10429
rect 55990 10365 56042 10371
rect 56086 10423 56138 10429
rect 56086 10365 56138 10371
rect 55702 10127 55754 10133
rect 55702 10069 55754 10075
rect 55606 9239 55658 9245
rect 55606 9181 55658 9187
rect 55222 9017 55274 9023
rect 55222 8959 55274 8965
rect 55234 4213 55262 8959
rect 55414 7019 55466 7025
rect 55414 6961 55466 6967
rect 55222 4207 55274 4213
rect 55222 4149 55274 4155
rect 55138 3612 55358 3640
rect 55222 3467 55274 3473
rect 55222 3409 55274 3415
rect 55234 800 55262 3409
rect 55330 800 55358 3612
rect 55426 800 55454 6961
rect 55606 4355 55658 4361
rect 55606 4297 55658 4303
rect 55618 800 55646 4297
rect 55714 800 55742 10069
rect 55798 7685 55850 7691
rect 55798 7627 55850 7633
rect 55810 800 55838 7627
rect 55894 3763 55946 3769
rect 55894 3705 55946 3711
rect 55906 800 55934 3705
rect 56098 800 56126 10365
rect 56470 10127 56522 10133
rect 56470 10069 56522 10075
rect 56182 7685 56234 7691
rect 56182 7627 56234 7633
rect 56194 800 56222 7627
rect 56374 6945 56426 6951
rect 56374 6887 56426 6893
rect 56278 3615 56330 3621
rect 56278 3557 56330 3563
rect 56290 800 56318 3557
rect 56386 3473 56414 6887
rect 56374 3467 56426 3473
rect 56374 3409 56426 3415
rect 56482 800 56510 10069
rect 56662 7685 56714 7691
rect 56662 7627 56714 7633
rect 56674 7214 56702 7627
rect 56578 7186 56702 7214
rect 56578 800 56606 7186
rect 56662 4355 56714 4361
rect 56662 4297 56714 4303
rect 56674 800 56702 4297
rect 56770 800 56798 10883
rect 56866 10577 56894 50251
rect 57346 40399 57374 55357
rect 58006 54897 58058 54903
rect 58006 54839 58058 54845
rect 57622 54231 57674 54237
rect 57622 54173 57674 54179
rect 57634 53867 57662 54173
rect 57622 53861 57674 53867
rect 57622 53803 57674 53809
rect 57622 53417 57674 53423
rect 57622 53359 57674 53365
rect 57334 40393 57386 40399
rect 57334 40335 57386 40341
rect 56950 34251 57002 34257
rect 56950 34193 57002 34199
rect 56962 12427 56990 34193
rect 57634 22491 57662 53359
rect 57622 22485 57674 22491
rect 57622 22427 57674 22433
rect 58018 15091 58046 54839
rect 58114 54385 58142 59200
rect 58594 56309 58622 59200
rect 58582 56303 58634 56309
rect 58582 56245 58634 56251
rect 59170 55199 59198 59200
rect 59158 55193 59210 55199
rect 59158 55135 59210 55141
rect 58102 54379 58154 54385
rect 58102 54321 58154 54327
rect 59650 53867 59678 59200
rect 59638 53861 59690 53867
rect 59638 53803 59690 53809
rect 58006 15085 58058 15091
rect 58006 15027 58058 15033
rect 56950 12421 57002 12427
rect 56950 12363 57002 12369
rect 57526 12273 57578 12279
rect 57526 12215 57578 12221
rect 57142 11459 57194 11465
rect 57142 11401 57194 11407
rect 56854 10571 56906 10577
rect 56854 10513 56906 10519
rect 56866 10281 56894 10513
rect 56854 10275 56906 10281
rect 56854 10217 56906 10223
rect 56950 8351 57002 8357
rect 56950 8293 57002 8299
rect 56854 6427 56906 6433
rect 56854 6369 56906 6375
rect 56866 3251 56894 6369
rect 56854 3245 56906 3251
rect 56854 3187 56906 3193
rect 56962 800 56990 8293
rect 57046 5021 57098 5027
rect 57046 4963 57098 4969
rect 57058 800 57086 4963
rect 57154 800 57182 11401
rect 57238 9017 57290 9023
rect 57238 8959 57290 8965
rect 57250 800 57278 8959
rect 57334 8943 57386 8949
rect 57334 8885 57386 8891
rect 57346 4287 57374 8885
rect 57430 5687 57482 5693
rect 57430 5629 57482 5635
rect 57334 4281 57386 4287
rect 57334 4223 57386 4229
rect 57442 800 57470 5629
rect 57538 800 57566 12215
rect 58198 11607 58250 11613
rect 58198 11549 58250 11555
rect 57622 9683 57674 9689
rect 57622 9625 57674 9631
rect 57634 800 57662 9625
rect 58102 6353 58154 6359
rect 58102 6295 58154 6301
rect 57814 4947 57866 4953
rect 57814 4889 57866 4895
rect 57826 800 57854 4889
rect 57910 4207 57962 4213
rect 57910 4149 57962 4155
rect 57922 800 57950 4149
rect 58006 3245 58058 3251
rect 58006 3187 58058 3193
rect 58018 800 58046 3187
rect 58114 800 58142 6295
rect 58210 3695 58238 11549
rect 58294 10867 58346 10873
rect 58294 10809 58346 10815
rect 58198 3689 58250 3695
rect 58198 3631 58250 3637
rect 58306 800 58334 10809
rect 58582 10127 58634 10133
rect 58582 10069 58634 10075
rect 58390 8277 58442 8283
rect 58390 8219 58442 8225
rect 58402 800 58430 8219
rect 58486 7019 58538 7025
rect 58486 6961 58538 6967
rect 58498 800 58526 6961
rect 58594 800 58622 10069
rect 58966 8573 59018 8579
rect 58966 8515 59018 8521
rect 58774 7759 58826 7765
rect 58774 7701 58826 7707
rect 58786 800 58814 7701
rect 58870 6279 58922 6285
rect 58870 6221 58922 6227
rect 58882 800 58910 6221
rect 58978 800 59006 8515
rect 59830 8203 59882 8209
rect 59830 8145 59882 8151
rect 59350 7463 59402 7469
rect 59350 7405 59402 7411
rect 59254 4873 59306 4879
rect 59254 4815 59306 4821
rect 59158 4281 59210 4287
rect 59158 4223 59210 4229
rect 59170 800 59198 4223
rect 59266 800 59294 4815
rect 59362 800 59390 7405
rect 59638 5613 59690 5619
rect 59638 5555 59690 5561
rect 59446 3467 59498 3473
rect 59446 3409 59498 3415
rect 59458 800 59486 3409
rect 59650 800 59678 5555
rect 59734 3689 59786 3695
rect 59734 3631 59786 3637
rect 59746 800 59774 3631
rect 59842 800 59870 8145
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< via2 >>
rect 4268 57302 4324 57304
rect 4348 57302 4404 57304
rect 4428 57302 4484 57304
rect 4508 57302 4564 57304
rect 4268 57250 4294 57302
rect 4294 57250 4324 57302
rect 4348 57250 4358 57302
rect 4358 57250 4404 57302
rect 4428 57250 4474 57302
rect 4474 57250 4484 57302
rect 4508 57250 4538 57302
rect 4538 57250 4564 57302
rect 4268 57248 4324 57250
rect 4348 57248 4404 57250
rect 4428 57248 4484 57250
rect 4508 57248 4564 57250
rect 4268 55970 4324 55972
rect 4348 55970 4404 55972
rect 4428 55970 4484 55972
rect 4508 55970 4564 55972
rect 4268 55918 4294 55970
rect 4294 55918 4324 55970
rect 4348 55918 4358 55970
rect 4358 55918 4404 55970
rect 4428 55918 4474 55970
rect 4474 55918 4484 55970
rect 4508 55918 4538 55970
rect 4538 55918 4564 55970
rect 4268 55916 4324 55918
rect 4348 55916 4404 55918
rect 4428 55916 4484 55918
rect 4508 55916 4564 55918
rect 4268 54638 4324 54640
rect 4348 54638 4404 54640
rect 4428 54638 4484 54640
rect 4508 54638 4564 54640
rect 4268 54586 4294 54638
rect 4294 54586 4324 54638
rect 4348 54586 4358 54638
rect 4358 54586 4404 54638
rect 4428 54586 4474 54638
rect 4474 54586 4484 54638
rect 4508 54586 4538 54638
rect 4538 54586 4564 54638
rect 4268 54584 4324 54586
rect 4348 54584 4404 54586
rect 4428 54584 4484 54586
rect 4508 54584 4564 54586
rect 4268 53306 4324 53308
rect 4348 53306 4404 53308
rect 4428 53306 4484 53308
rect 4508 53306 4564 53308
rect 4268 53254 4294 53306
rect 4294 53254 4324 53306
rect 4348 53254 4358 53306
rect 4358 53254 4404 53306
rect 4428 53254 4474 53306
rect 4474 53254 4484 53306
rect 4508 53254 4538 53306
rect 4538 53254 4564 53306
rect 4268 53252 4324 53254
rect 4348 53252 4404 53254
rect 4428 53252 4484 53254
rect 4508 53252 4564 53254
rect 4268 51974 4324 51976
rect 4348 51974 4404 51976
rect 4428 51974 4484 51976
rect 4508 51974 4564 51976
rect 4268 51922 4294 51974
rect 4294 51922 4324 51974
rect 4348 51922 4358 51974
rect 4358 51922 4404 51974
rect 4428 51922 4474 51974
rect 4474 51922 4484 51974
rect 4508 51922 4538 51974
rect 4538 51922 4564 51974
rect 4268 51920 4324 51922
rect 4348 51920 4404 51922
rect 4428 51920 4484 51922
rect 4508 51920 4564 51922
rect 4268 50642 4324 50644
rect 4348 50642 4404 50644
rect 4428 50642 4484 50644
rect 4508 50642 4564 50644
rect 4268 50590 4294 50642
rect 4294 50590 4324 50642
rect 4348 50590 4358 50642
rect 4358 50590 4404 50642
rect 4428 50590 4474 50642
rect 4474 50590 4484 50642
rect 4508 50590 4538 50642
rect 4538 50590 4564 50642
rect 4268 50588 4324 50590
rect 4348 50588 4404 50590
rect 4428 50588 4484 50590
rect 4508 50588 4564 50590
rect 4268 49310 4324 49312
rect 4348 49310 4404 49312
rect 4428 49310 4484 49312
rect 4508 49310 4564 49312
rect 4268 49258 4294 49310
rect 4294 49258 4324 49310
rect 4348 49258 4358 49310
rect 4358 49258 4404 49310
rect 4428 49258 4474 49310
rect 4474 49258 4484 49310
rect 4508 49258 4538 49310
rect 4538 49258 4564 49310
rect 4268 49256 4324 49258
rect 4348 49256 4404 49258
rect 4428 49256 4484 49258
rect 4508 49256 4564 49258
rect 4268 47978 4324 47980
rect 4348 47978 4404 47980
rect 4428 47978 4484 47980
rect 4508 47978 4564 47980
rect 4268 47926 4294 47978
rect 4294 47926 4324 47978
rect 4348 47926 4358 47978
rect 4358 47926 4404 47978
rect 4428 47926 4474 47978
rect 4474 47926 4484 47978
rect 4508 47926 4538 47978
rect 4538 47926 4564 47978
rect 4268 47924 4324 47926
rect 4348 47924 4404 47926
rect 4428 47924 4484 47926
rect 4508 47924 4564 47926
rect 4268 46646 4324 46648
rect 4348 46646 4404 46648
rect 4428 46646 4484 46648
rect 4508 46646 4564 46648
rect 4268 46594 4294 46646
rect 4294 46594 4324 46646
rect 4348 46594 4358 46646
rect 4358 46594 4404 46646
rect 4428 46594 4474 46646
rect 4474 46594 4484 46646
rect 4508 46594 4538 46646
rect 4538 46594 4564 46646
rect 4268 46592 4324 46594
rect 4348 46592 4404 46594
rect 4428 46592 4484 46594
rect 4508 46592 4564 46594
rect 4268 45314 4324 45316
rect 4348 45314 4404 45316
rect 4428 45314 4484 45316
rect 4508 45314 4564 45316
rect 4268 45262 4294 45314
rect 4294 45262 4324 45314
rect 4348 45262 4358 45314
rect 4358 45262 4404 45314
rect 4428 45262 4474 45314
rect 4474 45262 4484 45314
rect 4508 45262 4538 45314
rect 4538 45262 4564 45314
rect 4268 45260 4324 45262
rect 4348 45260 4404 45262
rect 4428 45260 4484 45262
rect 4508 45260 4564 45262
rect 4268 43982 4324 43984
rect 4348 43982 4404 43984
rect 4428 43982 4484 43984
rect 4508 43982 4564 43984
rect 4268 43930 4294 43982
rect 4294 43930 4324 43982
rect 4348 43930 4358 43982
rect 4358 43930 4404 43982
rect 4428 43930 4474 43982
rect 4474 43930 4484 43982
rect 4508 43930 4538 43982
rect 4538 43930 4564 43982
rect 4268 43928 4324 43930
rect 4348 43928 4404 43930
rect 4428 43928 4484 43930
rect 4508 43928 4564 43930
rect 4268 42650 4324 42652
rect 4348 42650 4404 42652
rect 4428 42650 4484 42652
rect 4508 42650 4564 42652
rect 4268 42598 4294 42650
rect 4294 42598 4324 42650
rect 4348 42598 4358 42650
rect 4358 42598 4404 42650
rect 4428 42598 4474 42650
rect 4474 42598 4484 42650
rect 4508 42598 4538 42650
rect 4538 42598 4564 42650
rect 4268 42596 4324 42598
rect 4348 42596 4404 42598
rect 4428 42596 4484 42598
rect 4508 42596 4564 42598
rect 4268 41318 4324 41320
rect 4348 41318 4404 41320
rect 4428 41318 4484 41320
rect 4508 41318 4564 41320
rect 4268 41266 4294 41318
rect 4294 41266 4324 41318
rect 4348 41266 4358 41318
rect 4358 41266 4404 41318
rect 4428 41266 4474 41318
rect 4474 41266 4484 41318
rect 4508 41266 4538 41318
rect 4538 41266 4564 41318
rect 4268 41264 4324 41266
rect 4348 41264 4404 41266
rect 4428 41264 4484 41266
rect 4508 41264 4564 41266
rect 4268 39986 4324 39988
rect 4348 39986 4404 39988
rect 4428 39986 4484 39988
rect 4508 39986 4564 39988
rect 4268 39934 4294 39986
rect 4294 39934 4324 39986
rect 4348 39934 4358 39986
rect 4358 39934 4404 39986
rect 4428 39934 4474 39986
rect 4474 39934 4484 39986
rect 4508 39934 4538 39986
rect 4538 39934 4564 39986
rect 4268 39932 4324 39934
rect 4348 39932 4404 39934
rect 4428 39932 4484 39934
rect 4508 39932 4564 39934
rect 4268 38654 4324 38656
rect 4348 38654 4404 38656
rect 4428 38654 4484 38656
rect 4508 38654 4564 38656
rect 4268 38602 4294 38654
rect 4294 38602 4324 38654
rect 4348 38602 4358 38654
rect 4358 38602 4404 38654
rect 4428 38602 4474 38654
rect 4474 38602 4484 38654
rect 4508 38602 4538 38654
rect 4538 38602 4564 38654
rect 4268 38600 4324 38602
rect 4348 38600 4404 38602
rect 4428 38600 4484 38602
rect 4508 38600 4564 38602
rect 4268 37322 4324 37324
rect 4348 37322 4404 37324
rect 4428 37322 4484 37324
rect 4508 37322 4564 37324
rect 4268 37270 4294 37322
rect 4294 37270 4324 37322
rect 4348 37270 4358 37322
rect 4358 37270 4404 37322
rect 4428 37270 4474 37322
rect 4474 37270 4484 37322
rect 4508 37270 4538 37322
rect 4538 37270 4564 37322
rect 4268 37268 4324 37270
rect 4348 37268 4404 37270
rect 4428 37268 4484 37270
rect 4508 37268 4564 37270
rect 4268 35990 4324 35992
rect 4348 35990 4404 35992
rect 4428 35990 4484 35992
rect 4508 35990 4564 35992
rect 4268 35938 4294 35990
rect 4294 35938 4324 35990
rect 4348 35938 4358 35990
rect 4358 35938 4404 35990
rect 4428 35938 4474 35990
rect 4474 35938 4484 35990
rect 4508 35938 4538 35990
rect 4538 35938 4564 35990
rect 4268 35936 4324 35938
rect 4348 35936 4404 35938
rect 4428 35936 4484 35938
rect 4508 35936 4564 35938
rect 4268 34658 4324 34660
rect 4348 34658 4404 34660
rect 4428 34658 4484 34660
rect 4508 34658 4564 34660
rect 4268 34606 4294 34658
rect 4294 34606 4324 34658
rect 4348 34606 4358 34658
rect 4358 34606 4404 34658
rect 4428 34606 4474 34658
rect 4474 34606 4484 34658
rect 4508 34606 4538 34658
rect 4538 34606 4564 34658
rect 4268 34604 4324 34606
rect 4348 34604 4404 34606
rect 4428 34604 4484 34606
rect 4508 34604 4564 34606
rect 4268 33326 4324 33328
rect 4348 33326 4404 33328
rect 4428 33326 4484 33328
rect 4508 33326 4564 33328
rect 4268 33274 4294 33326
rect 4294 33274 4324 33326
rect 4348 33274 4358 33326
rect 4358 33274 4404 33326
rect 4428 33274 4474 33326
rect 4474 33274 4484 33326
rect 4508 33274 4538 33326
rect 4538 33274 4564 33326
rect 4268 33272 4324 33274
rect 4348 33272 4404 33274
rect 4428 33272 4484 33274
rect 4508 33272 4564 33274
rect 4268 31994 4324 31996
rect 4348 31994 4404 31996
rect 4428 31994 4484 31996
rect 4508 31994 4564 31996
rect 4268 31942 4294 31994
rect 4294 31942 4324 31994
rect 4348 31942 4358 31994
rect 4358 31942 4404 31994
rect 4428 31942 4474 31994
rect 4474 31942 4484 31994
rect 4508 31942 4538 31994
rect 4538 31942 4564 31994
rect 4268 31940 4324 31942
rect 4348 31940 4404 31942
rect 4428 31940 4484 31942
rect 4508 31940 4564 31942
rect 4268 30662 4324 30664
rect 4348 30662 4404 30664
rect 4428 30662 4484 30664
rect 4508 30662 4564 30664
rect 4268 30610 4294 30662
rect 4294 30610 4324 30662
rect 4348 30610 4358 30662
rect 4358 30610 4404 30662
rect 4428 30610 4474 30662
rect 4474 30610 4484 30662
rect 4508 30610 4538 30662
rect 4538 30610 4564 30662
rect 4268 30608 4324 30610
rect 4348 30608 4404 30610
rect 4428 30608 4484 30610
rect 4508 30608 4564 30610
rect 4268 29330 4324 29332
rect 4348 29330 4404 29332
rect 4428 29330 4484 29332
rect 4508 29330 4564 29332
rect 4268 29278 4294 29330
rect 4294 29278 4324 29330
rect 4348 29278 4358 29330
rect 4358 29278 4404 29330
rect 4428 29278 4474 29330
rect 4474 29278 4484 29330
rect 4508 29278 4538 29330
rect 4538 29278 4564 29330
rect 4268 29276 4324 29278
rect 4348 29276 4404 29278
rect 4428 29276 4484 29278
rect 4508 29276 4564 29278
rect 4268 27998 4324 28000
rect 4348 27998 4404 28000
rect 4428 27998 4484 28000
rect 4508 27998 4564 28000
rect 4268 27946 4294 27998
rect 4294 27946 4324 27998
rect 4348 27946 4358 27998
rect 4358 27946 4404 27998
rect 4428 27946 4474 27998
rect 4474 27946 4484 27998
rect 4508 27946 4538 27998
rect 4538 27946 4564 27998
rect 4268 27944 4324 27946
rect 4348 27944 4404 27946
rect 4428 27944 4484 27946
rect 4508 27944 4564 27946
rect 4268 26666 4324 26668
rect 4348 26666 4404 26668
rect 4428 26666 4484 26668
rect 4508 26666 4564 26668
rect 4268 26614 4294 26666
rect 4294 26614 4324 26666
rect 4348 26614 4358 26666
rect 4358 26614 4404 26666
rect 4428 26614 4474 26666
rect 4474 26614 4484 26666
rect 4508 26614 4538 26666
rect 4538 26614 4564 26666
rect 4268 26612 4324 26614
rect 4348 26612 4404 26614
rect 4428 26612 4484 26614
rect 4508 26612 4564 26614
rect 4268 25334 4324 25336
rect 4348 25334 4404 25336
rect 4428 25334 4484 25336
rect 4508 25334 4564 25336
rect 4268 25282 4294 25334
rect 4294 25282 4324 25334
rect 4348 25282 4358 25334
rect 4358 25282 4404 25334
rect 4428 25282 4474 25334
rect 4474 25282 4484 25334
rect 4508 25282 4538 25334
rect 4538 25282 4564 25334
rect 4268 25280 4324 25282
rect 4348 25280 4404 25282
rect 4428 25280 4484 25282
rect 4508 25280 4564 25282
rect 4268 24002 4324 24004
rect 4348 24002 4404 24004
rect 4428 24002 4484 24004
rect 4508 24002 4564 24004
rect 4268 23950 4294 24002
rect 4294 23950 4324 24002
rect 4348 23950 4358 24002
rect 4358 23950 4404 24002
rect 4428 23950 4474 24002
rect 4474 23950 4484 24002
rect 4508 23950 4538 24002
rect 4538 23950 4564 24002
rect 4268 23948 4324 23950
rect 4348 23948 4404 23950
rect 4428 23948 4484 23950
rect 4508 23948 4564 23950
rect 4268 22670 4324 22672
rect 4348 22670 4404 22672
rect 4428 22670 4484 22672
rect 4508 22670 4564 22672
rect 4268 22618 4294 22670
rect 4294 22618 4324 22670
rect 4348 22618 4358 22670
rect 4358 22618 4404 22670
rect 4428 22618 4474 22670
rect 4474 22618 4484 22670
rect 4508 22618 4538 22670
rect 4538 22618 4564 22670
rect 4268 22616 4324 22618
rect 4348 22616 4404 22618
rect 4428 22616 4484 22618
rect 4508 22616 4564 22618
rect 4268 21338 4324 21340
rect 4348 21338 4404 21340
rect 4428 21338 4484 21340
rect 4508 21338 4564 21340
rect 4268 21286 4294 21338
rect 4294 21286 4324 21338
rect 4348 21286 4358 21338
rect 4358 21286 4404 21338
rect 4428 21286 4474 21338
rect 4474 21286 4484 21338
rect 4508 21286 4538 21338
rect 4538 21286 4564 21338
rect 4268 21284 4324 21286
rect 4348 21284 4404 21286
rect 4428 21284 4484 21286
rect 4508 21284 4564 21286
rect 4268 20006 4324 20008
rect 4348 20006 4404 20008
rect 4428 20006 4484 20008
rect 4508 20006 4564 20008
rect 4268 19954 4294 20006
rect 4294 19954 4324 20006
rect 4348 19954 4358 20006
rect 4358 19954 4404 20006
rect 4428 19954 4474 20006
rect 4474 19954 4484 20006
rect 4508 19954 4538 20006
rect 4538 19954 4564 20006
rect 4268 19952 4324 19954
rect 4348 19952 4404 19954
rect 4428 19952 4484 19954
rect 4508 19952 4564 19954
rect 4268 18674 4324 18676
rect 4348 18674 4404 18676
rect 4428 18674 4484 18676
rect 4508 18674 4564 18676
rect 4268 18622 4294 18674
rect 4294 18622 4324 18674
rect 4348 18622 4358 18674
rect 4358 18622 4404 18674
rect 4428 18622 4474 18674
rect 4474 18622 4484 18674
rect 4508 18622 4538 18674
rect 4538 18622 4564 18674
rect 4268 18620 4324 18622
rect 4348 18620 4404 18622
rect 4428 18620 4484 18622
rect 4508 18620 4564 18622
rect 4268 17342 4324 17344
rect 4348 17342 4404 17344
rect 4428 17342 4484 17344
rect 4508 17342 4564 17344
rect 4268 17290 4294 17342
rect 4294 17290 4324 17342
rect 4348 17290 4358 17342
rect 4358 17290 4404 17342
rect 4428 17290 4474 17342
rect 4474 17290 4484 17342
rect 4508 17290 4538 17342
rect 4538 17290 4564 17342
rect 4268 17288 4324 17290
rect 4348 17288 4404 17290
rect 4428 17288 4484 17290
rect 4508 17288 4564 17290
rect 4268 16010 4324 16012
rect 4348 16010 4404 16012
rect 4428 16010 4484 16012
rect 4508 16010 4564 16012
rect 4268 15958 4294 16010
rect 4294 15958 4324 16010
rect 4348 15958 4358 16010
rect 4358 15958 4404 16010
rect 4428 15958 4474 16010
rect 4474 15958 4484 16010
rect 4508 15958 4538 16010
rect 4538 15958 4564 16010
rect 4268 15956 4324 15958
rect 4348 15956 4404 15958
rect 4428 15956 4484 15958
rect 4508 15956 4564 15958
rect 4268 14678 4324 14680
rect 4348 14678 4404 14680
rect 4428 14678 4484 14680
rect 4508 14678 4564 14680
rect 4268 14626 4294 14678
rect 4294 14626 4324 14678
rect 4348 14626 4358 14678
rect 4358 14626 4404 14678
rect 4428 14626 4474 14678
rect 4474 14626 4484 14678
rect 4508 14626 4538 14678
rect 4538 14626 4564 14678
rect 4268 14624 4324 14626
rect 4348 14624 4404 14626
rect 4428 14624 4484 14626
rect 4508 14624 4564 14626
rect 4268 13346 4324 13348
rect 4348 13346 4404 13348
rect 4428 13346 4484 13348
rect 4508 13346 4564 13348
rect 4268 13294 4294 13346
rect 4294 13294 4324 13346
rect 4348 13294 4358 13346
rect 4358 13294 4404 13346
rect 4428 13294 4474 13346
rect 4474 13294 4484 13346
rect 4508 13294 4538 13346
rect 4538 13294 4564 13346
rect 4268 13292 4324 13294
rect 4348 13292 4404 13294
rect 4428 13292 4484 13294
rect 4508 13292 4564 13294
rect 4268 12014 4324 12016
rect 4348 12014 4404 12016
rect 4428 12014 4484 12016
rect 4508 12014 4564 12016
rect 4268 11962 4294 12014
rect 4294 11962 4324 12014
rect 4348 11962 4358 12014
rect 4358 11962 4404 12014
rect 4428 11962 4474 12014
rect 4474 11962 4484 12014
rect 4508 11962 4538 12014
rect 4538 11962 4564 12014
rect 4268 11960 4324 11962
rect 4348 11960 4404 11962
rect 4428 11960 4484 11962
rect 4508 11960 4564 11962
rect 4268 10682 4324 10684
rect 4348 10682 4404 10684
rect 4428 10682 4484 10684
rect 4508 10682 4564 10684
rect 4268 10630 4294 10682
rect 4294 10630 4324 10682
rect 4348 10630 4358 10682
rect 4358 10630 4404 10682
rect 4428 10630 4474 10682
rect 4474 10630 4484 10682
rect 4508 10630 4538 10682
rect 4538 10630 4564 10682
rect 4268 10628 4324 10630
rect 4348 10628 4404 10630
rect 4428 10628 4484 10630
rect 4508 10628 4564 10630
rect 4268 9350 4324 9352
rect 4348 9350 4404 9352
rect 4428 9350 4484 9352
rect 4508 9350 4564 9352
rect 4268 9298 4294 9350
rect 4294 9298 4324 9350
rect 4348 9298 4358 9350
rect 4358 9298 4404 9350
rect 4428 9298 4474 9350
rect 4474 9298 4484 9350
rect 4508 9298 4538 9350
rect 4538 9298 4564 9350
rect 4268 9296 4324 9298
rect 4348 9296 4404 9298
rect 4428 9296 4484 9298
rect 4508 9296 4564 9298
rect 4268 8018 4324 8020
rect 4348 8018 4404 8020
rect 4428 8018 4484 8020
rect 4508 8018 4564 8020
rect 4268 7966 4294 8018
rect 4294 7966 4324 8018
rect 4348 7966 4358 8018
rect 4358 7966 4404 8018
rect 4428 7966 4474 8018
rect 4474 7966 4484 8018
rect 4508 7966 4538 8018
rect 4538 7966 4564 8018
rect 4268 7964 4324 7966
rect 4348 7964 4404 7966
rect 4428 7964 4484 7966
rect 4508 7964 4564 7966
rect 4268 6686 4324 6688
rect 4348 6686 4404 6688
rect 4428 6686 4484 6688
rect 4508 6686 4564 6688
rect 4268 6634 4294 6686
rect 4294 6634 4324 6686
rect 4348 6634 4358 6686
rect 4358 6634 4404 6686
rect 4428 6634 4474 6686
rect 4474 6634 4484 6686
rect 4508 6634 4538 6686
rect 4538 6634 4564 6686
rect 4268 6632 4324 6634
rect 4348 6632 4404 6634
rect 4428 6632 4484 6634
rect 4508 6632 4564 6634
rect 4268 5354 4324 5356
rect 4348 5354 4404 5356
rect 4428 5354 4484 5356
rect 4508 5354 4564 5356
rect 4268 5302 4294 5354
rect 4294 5302 4324 5354
rect 4348 5302 4358 5354
rect 4358 5302 4404 5354
rect 4428 5302 4474 5354
rect 4474 5302 4484 5354
rect 4508 5302 4538 5354
rect 4538 5302 4564 5354
rect 4268 5300 4324 5302
rect 4348 5300 4404 5302
rect 4428 5300 4484 5302
rect 4508 5300 4564 5302
rect 4268 4022 4324 4024
rect 4348 4022 4404 4024
rect 4428 4022 4484 4024
rect 4508 4022 4564 4024
rect 4268 3970 4294 4022
rect 4294 3970 4324 4022
rect 4348 3970 4358 4022
rect 4358 3970 4404 4022
rect 4428 3970 4474 4022
rect 4474 3970 4484 4022
rect 4508 3970 4538 4022
rect 4538 3970 4564 4022
rect 4268 3968 4324 3970
rect 4348 3968 4404 3970
rect 4428 3968 4484 3970
rect 4508 3968 4564 3970
rect 4268 2690 4324 2692
rect 4348 2690 4404 2692
rect 4428 2690 4484 2692
rect 4508 2690 4564 2692
rect 4268 2638 4294 2690
rect 4294 2638 4324 2690
rect 4348 2638 4358 2690
rect 4358 2638 4404 2690
rect 4428 2638 4474 2690
rect 4474 2638 4484 2690
rect 4508 2638 4538 2690
rect 4538 2638 4564 2690
rect 4268 2636 4324 2638
rect 4348 2636 4404 2638
rect 4428 2636 4484 2638
rect 4508 2636 4564 2638
rect 8276 19473 8278 19490
rect 8278 19473 8330 19490
rect 8330 19473 8332 19490
rect 8276 19434 8332 19473
rect 9044 19473 9046 19490
rect 9046 19473 9098 19490
rect 9098 19473 9100 19490
rect 9044 19434 9100 19473
rect 7940 7759 7996 7798
rect 7940 7742 7942 7759
rect 7942 7742 7994 7759
rect 7994 7742 7996 7759
rect 12980 7742 13036 7798
rect 19628 56636 19684 56638
rect 19708 56636 19764 56638
rect 19788 56636 19844 56638
rect 19868 56636 19924 56638
rect 19628 56584 19654 56636
rect 19654 56584 19684 56636
rect 19708 56584 19718 56636
rect 19718 56584 19764 56636
rect 19788 56584 19834 56636
rect 19834 56584 19844 56636
rect 19868 56584 19898 56636
rect 19898 56584 19924 56636
rect 19628 56582 19684 56584
rect 19708 56582 19764 56584
rect 19788 56582 19844 56584
rect 19868 56582 19924 56584
rect 19628 55304 19684 55306
rect 19708 55304 19764 55306
rect 19788 55304 19844 55306
rect 19868 55304 19924 55306
rect 19628 55252 19654 55304
rect 19654 55252 19684 55304
rect 19708 55252 19718 55304
rect 19718 55252 19764 55304
rect 19788 55252 19834 55304
rect 19834 55252 19844 55304
rect 19868 55252 19898 55304
rect 19898 55252 19924 55304
rect 19628 55250 19684 55252
rect 19708 55250 19764 55252
rect 19788 55250 19844 55252
rect 19868 55250 19924 55252
rect 19628 53972 19684 53974
rect 19708 53972 19764 53974
rect 19788 53972 19844 53974
rect 19868 53972 19924 53974
rect 19628 53920 19654 53972
rect 19654 53920 19684 53972
rect 19708 53920 19718 53972
rect 19718 53920 19764 53972
rect 19788 53920 19834 53972
rect 19834 53920 19844 53972
rect 19868 53920 19898 53972
rect 19898 53920 19924 53972
rect 19628 53918 19684 53920
rect 19708 53918 19764 53920
rect 19788 53918 19844 53920
rect 19868 53918 19924 53920
rect 19628 52640 19684 52642
rect 19708 52640 19764 52642
rect 19788 52640 19844 52642
rect 19868 52640 19924 52642
rect 19628 52588 19654 52640
rect 19654 52588 19684 52640
rect 19708 52588 19718 52640
rect 19718 52588 19764 52640
rect 19788 52588 19834 52640
rect 19834 52588 19844 52640
rect 19868 52588 19898 52640
rect 19898 52588 19924 52640
rect 19628 52586 19684 52588
rect 19708 52586 19764 52588
rect 19788 52586 19844 52588
rect 19868 52586 19924 52588
rect 19628 51308 19684 51310
rect 19708 51308 19764 51310
rect 19788 51308 19844 51310
rect 19868 51308 19924 51310
rect 19628 51256 19654 51308
rect 19654 51256 19684 51308
rect 19708 51256 19718 51308
rect 19718 51256 19764 51308
rect 19788 51256 19834 51308
rect 19834 51256 19844 51308
rect 19868 51256 19898 51308
rect 19898 51256 19924 51308
rect 19628 51254 19684 51256
rect 19708 51254 19764 51256
rect 19788 51254 19844 51256
rect 19868 51254 19924 51256
rect 19628 49976 19684 49978
rect 19708 49976 19764 49978
rect 19788 49976 19844 49978
rect 19868 49976 19924 49978
rect 19628 49924 19654 49976
rect 19654 49924 19684 49976
rect 19708 49924 19718 49976
rect 19718 49924 19764 49976
rect 19788 49924 19834 49976
rect 19834 49924 19844 49976
rect 19868 49924 19898 49976
rect 19898 49924 19924 49976
rect 19628 49922 19684 49924
rect 19708 49922 19764 49924
rect 19788 49922 19844 49924
rect 19868 49922 19924 49924
rect 19628 48644 19684 48646
rect 19708 48644 19764 48646
rect 19788 48644 19844 48646
rect 19868 48644 19924 48646
rect 19628 48592 19654 48644
rect 19654 48592 19684 48644
rect 19708 48592 19718 48644
rect 19718 48592 19764 48644
rect 19788 48592 19834 48644
rect 19834 48592 19844 48644
rect 19868 48592 19898 48644
rect 19898 48592 19924 48644
rect 19628 48590 19684 48592
rect 19708 48590 19764 48592
rect 19788 48590 19844 48592
rect 19868 48590 19924 48592
rect 19628 47312 19684 47314
rect 19708 47312 19764 47314
rect 19788 47312 19844 47314
rect 19868 47312 19924 47314
rect 19628 47260 19654 47312
rect 19654 47260 19684 47312
rect 19708 47260 19718 47312
rect 19718 47260 19764 47312
rect 19788 47260 19834 47312
rect 19834 47260 19844 47312
rect 19868 47260 19898 47312
rect 19898 47260 19924 47312
rect 19628 47258 19684 47260
rect 19708 47258 19764 47260
rect 19788 47258 19844 47260
rect 19868 47258 19924 47260
rect 19628 45980 19684 45982
rect 19708 45980 19764 45982
rect 19788 45980 19844 45982
rect 19868 45980 19924 45982
rect 19628 45928 19654 45980
rect 19654 45928 19684 45980
rect 19708 45928 19718 45980
rect 19718 45928 19764 45980
rect 19788 45928 19834 45980
rect 19834 45928 19844 45980
rect 19868 45928 19898 45980
rect 19898 45928 19924 45980
rect 19628 45926 19684 45928
rect 19708 45926 19764 45928
rect 19788 45926 19844 45928
rect 19868 45926 19924 45928
rect 19628 44648 19684 44650
rect 19708 44648 19764 44650
rect 19788 44648 19844 44650
rect 19868 44648 19924 44650
rect 19628 44596 19654 44648
rect 19654 44596 19684 44648
rect 19708 44596 19718 44648
rect 19718 44596 19764 44648
rect 19788 44596 19834 44648
rect 19834 44596 19844 44648
rect 19868 44596 19898 44648
rect 19898 44596 19924 44648
rect 19628 44594 19684 44596
rect 19708 44594 19764 44596
rect 19788 44594 19844 44596
rect 19868 44594 19924 44596
rect 19628 43316 19684 43318
rect 19708 43316 19764 43318
rect 19788 43316 19844 43318
rect 19868 43316 19924 43318
rect 19628 43264 19654 43316
rect 19654 43264 19684 43316
rect 19708 43264 19718 43316
rect 19718 43264 19764 43316
rect 19788 43264 19834 43316
rect 19834 43264 19844 43316
rect 19868 43264 19898 43316
rect 19898 43264 19924 43316
rect 19628 43262 19684 43264
rect 19708 43262 19764 43264
rect 19788 43262 19844 43264
rect 19868 43262 19924 43264
rect 19628 41984 19684 41986
rect 19708 41984 19764 41986
rect 19788 41984 19844 41986
rect 19868 41984 19924 41986
rect 19628 41932 19654 41984
rect 19654 41932 19684 41984
rect 19708 41932 19718 41984
rect 19718 41932 19764 41984
rect 19788 41932 19834 41984
rect 19834 41932 19844 41984
rect 19868 41932 19898 41984
rect 19898 41932 19924 41984
rect 19628 41930 19684 41932
rect 19708 41930 19764 41932
rect 19788 41930 19844 41932
rect 19868 41930 19924 41932
rect 19628 40652 19684 40654
rect 19708 40652 19764 40654
rect 19788 40652 19844 40654
rect 19868 40652 19924 40654
rect 19628 40600 19654 40652
rect 19654 40600 19684 40652
rect 19708 40600 19718 40652
rect 19718 40600 19764 40652
rect 19788 40600 19834 40652
rect 19834 40600 19844 40652
rect 19868 40600 19898 40652
rect 19898 40600 19924 40652
rect 19628 40598 19684 40600
rect 19708 40598 19764 40600
rect 19788 40598 19844 40600
rect 19868 40598 19924 40600
rect 19628 39320 19684 39322
rect 19708 39320 19764 39322
rect 19788 39320 19844 39322
rect 19868 39320 19924 39322
rect 19628 39268 19654 39320
rect 19654 39268 19684 39320
rect 19708 39268 19718 39320
rect 19718 39268 19764 39320
rect 19788 39268 19834 39320
rect 19834 39268 19844 39320
rect 19868 39268 19898 39320
rect 19898 39268 19924 39320
rect 19628 39266 19684 39268
rect 19708 39266 19764 39268
rect 19788 39266 19844 39268
rect 19868 39266 19924 39268
rect 19628 37988 19684 37990
rect 19708 37988 19764 37990
rect 19788 37988 19844 37990
rect 19868 37988 19924 37990
rect 19628 37936 19654 37988
rect 19654 37936 19684 37988
rect 19708 37936 19718 37988
rect 19718 37936 19764 37988
rect 19788 37936 19834 37988
rect 19834 37936 19844 37988
rect 19868 37936 19898 37988
rect 19898 37936 19924 37988
rect 19628 37934 19684 37936
rect 19708 37934 19764 37936
rect 19788 37934 19844 37936
rect 19868 37934 19924 37936
rect 19628 36656 19684 36658
rect 19708 36656 19764 36658
rect 19788 36656 19844 36658
rect 19868 36656 19924 36658
rect 19628 36604 19654 36656
rect 19654 36604 19684 36656
rect 19708 36604 19718 36656
rect 19718 36604 19764 36656
rect 19788 36604 19834 36656
rect 19834 36604 19844 36656
rect 19868 36604 19898 36656
rect 19898 36604 19924 36656
rect 19628 36602 19684 36604
rect 19708 36602 19764 36604
rect 19788 36602 19844 36604
rect 19868 36602 19924 36604
rect 19628 35324 19684 35326
rect 19708 35324 19764 35326
rect 19788 35324 19844 35326
rect 19868 35324 19924 35326
rect 19628 35272 19654 35324
rect 19654 35272 19684 35324
rect 19708 35272 19718 35324
rect 19718 35272 19764 35324
rect 19788 35272 19834 35324
rect 19834 35272 19844 35324
rect 19868 35272 19898 35324
rect 19898 35272 19924 35324
rect 19628 35270 19684 35272
rect 19708 35270 19764 35272
rect 19788 35270 19844 35272
rect 19868 35270 19924 35272
rect 19628 33992 19684 33994
rect 19708 33992 19764 33994
rect 19788 33992 19844 33994
rect 19868 33992 19924 33994
rect 19628 33940 19654 33992
rect 19654 33940 19684 33992
rect 19708 33940 19718 33992
rect 19718 33940 19764 33992
rect 19788 33940 19834 33992
rect 19834 33940 19844 33992
rect 19868 33940 19898 33992
rect 19898 33940 19924 33992
rect 19628 33938 19684 33940
rect 19708 33938 19764 33940
rect 19788 33938 19844 33940
rect 19868 33938 19924 33940
rect 19628 32660 19684 32662
rect 19708 32660 19764 32662
rect 19788 32660 19844 32662
rect 19868 32660 19924 32662
rect 19628 32608 19654 32660
rect 19654 32608 19684 32660
rect 19708 32608 19718 32660
rect 19718 32608 19764 32660
rect 19788 32608 19834 32660
rect 19834 32608 19844 32660
rect 19868 32608 19898 32660
rect 19898 32608 19924 32660
rect 19628 32606 19684 32608
rect 19708 32606 19764 32608
rect 19788 32606 19844 32608
rect 19868 32606 19924 32608
rect 19628 31328 19684 31330
rect 19708 31328 19764 31330
rect 19788 31328 19844 31330
rect 19868 31328 19924 31330
rect 19628 31276 19654 31328
rect 19654 31276 19684 31328
rect 19708 31276 19718 31328
rect 19718 31276 19764 31328
rect 19788 31276 19834 31328
rect 19834 31276 19844 31328
rect 19868 31276 19898 31328
rect 19898 31276 19924 31328
rect 19628 31274 19684 31276
rect 19708 31274 19764 31276
rect 19788 31274 19844 31276
rect 19868 31274 19924 31276
rect 19628 29996 19684 29998
rect 19708 29996 19764 29998
rect 19788 29996 19844 29998
rect 19868 29996 19924 29998
rect 19628 29944 19654 29996
rect 19654 29944 19684 29996
rect 19708 29944 19718 29996
rect 19718 29944 19764 29996
rect 19788 29944 19834 29996
rect 19834 29944 19844 29996
rect 19868 29944 19898 29996
rect 19898 29944 19924 29996
rect 19628 29942 19684 29944
rect 19708 29942 19764 29944
rect 19788 29942 19844 29944
rect 19868 29942 19924 29944
rect 19628 28664 19684 28666
rect 19708 28664 19764 28666
rect 19788 28664 19844 28666
rect 19868 28664 19924 28666
rect 19628 28612 19654 28664
rect 19654 28612 19684 28664
rect 19708 28612 19718 28664
rect 19718 28612 19764 28664
rect 19788 28612 19834 28664
rect 19834 28612 19844 28664
rect 19868 28612 19898 28664
rect 19898 28612 19924 28664
rect 19628 28610 19684 28612
rect 19708 28610 19764 28612
rect 19788 28610 19844 28612
rect 19868 28610 19924 28612
rect 19628 27332 19684 27334
rect 19708 27332 19764 27334
rect 19788 27332 19844 27334
rect 19868 27332 19924 27334
rect 19628 27280 19654 27332
rect 19654 27280 19684 27332
rect 19708 27280 19718 27332
rect 19718 27280 19764 27332
rect 19788 27280 19834 27332
rect 19834 27280 19844 27332
rect 19868 27280 19898 27332
rect 19898 27280 19924 27332
rect 19628 27278 19684 27280
rect 19708 27278 19764 27280
rect 19788 27278 19844 27280
rect 19868 27278 19924 27280
rect 19628 26000 19684 26002
rect 19708 26000 19764 26002
rect 19788 26000 19844 26002
rect 19868 26000 19924 26002
rect 19628 25948 19654 26000
rect 19654 25948 19684 26000
rect 19708 25948 19718 26000
rect 19718 25948 19764 26000
rect 19788 25948 19834 26000
rect 19834 25948 19844 26000
rect 19868 25948 19898 26000
rect 19898 25948 19924 26000
rect 19628 25946 19684 25948
rect 19708 25946 19764 25948
rect 19788 25946 19844 25948
rect 19868 25946 19924 25948
rect 19628 24668 19684 24670
rect 19708 24668 19764 24670
rect 19788 24668 19844 24670
rect 19868 24668 19924 24670
rect 19628 24616 19654 24668
rect 19654 24616 19684 24668
rect 19708 24616 19718 24668
rect 19718 24616 19764 24668
rect 19788 24616 19834 24668
rect 19834 24616 19844 24668
rect 19868 24616 19898 24668
rect 19898 24616 19924 24668
rect 19628 24614 19684 24616
rect 19708 24614 19764 24616
rect 19788 24614 19844 24616
rect 19868 24614 19924 24616
rect 19628 23336 19684 23338
rect 19708 23336 19764 23338
rect 19788 23336 19844 23338
rect 19868 23336 19924 23338
rect 19628 23284 19654 23336
rect 19654 23284 19684 23336
rect 19708 23284 19718 23336
rect 19718 23284 19764 23336
rect 19788 23284 19834 23336
rect 19834 23284 19844 23336
rect 19868 23284 19898 23336
rect 19898 23284 19924 23336
rect 19628 23282 19684 23284
rect 19708 23282 19764 23284
rect 19788 23282 19844 23284
rect 19868 23282 19924 23284
rect 19628 22004 19684 22006
rect 19708 22004 19764 22006
rect 19788 22004 19844 22006
rect 19868 22004 19924 22006
rect 19628 21952 19654 22004
rect 19654 21952 19684 22004
rect 19708 21952 19718 22004
rect 19718 21952 19764 22004
rect 19788 21952 19834 22004
rect 19834 21952 19844 22004
rect 19868 21952 19898 22004
rect 19898 21952 19924 22004
rect 19628 21950 19684 21952
rect 19708 21950 19764 21952
rect 19788 21950 19844 21952
rect 19868 21950 19924 21952
rect 19628 20672 19684 20674
rect 19708 20672 19764 20674
rect 19788 20672 19844 20674
rect 19868 20672 19924 20674
rect 19628 20620 19654 20672
rect 19654 20620 19684 20672
rect 19708 20620 19718 20672
rect 19718 20620 19764 20672
rect 19788 20620 19834 20672
rect 19834 20620 19844 20672
rect 19868 20620 19898 20672
rect 19898 20620 19924 20672
rect 19628 20618 19684 20620
rect 19708 20618 19764 20620
rect 19788 20618 19844 20620
rect 19868 20618 19924 20620
rect 19628 19340 19684 19342
rect 19708 19340 19764 19342
rect 19788 19340 19844 19342
rect 19868 19340 19924 19342
rect 19628 19288 19654 19340
rect 19654 19288 19684 19340
rect 19708 19288 19718 19340
rect 19718 19288 19764 19340
rect 19788 19288 19834 19340
rect 19834 19288 19844 19340
rect 19868 19288 19898 19340
rect 19898 19288 19924 19340
rect 19628 19286 19684 19288
rect 19708 19286 19764 19288
rect 19788 19286 19844 19288
rect 19868 19286 19924 19288
rect 19628 18008 19684 18010
rect 19708 18008 19764 18010
rect 19788 18008 19844 18010
rect 19868 18008 19924 18010
rect 19628 17956 19654 18008
rect 19654 17956 19684 18008
rect 19708 17956 19718 18008
rect 19718 17956 19764 18008
rect 19788 17956 19834 18008
rect 19834 17956 19844 18008
rect 19868 17956 19898 18008
rect 19898 17956 19924 18008
rect 19628 17954 19684 17956
rect 19708 17954 19764 17956
rect 19788 17954 19844 17956
rect 19868 17954 19924 17956
rect 19628 16676 19684 16678
rect 19708 16676 19764 16678
rect 19788 16676 19844 16678
rect 19868 16676 19924 16678
rect 19628 16624 19654 16676
rect 19654 16624 19684 16676
rect 19708 16624 19718 16676
rect 19718 16624 19764 16676
rect 19788 16624 19834 16676
rect 19834 16624 19844 16676
rect 19868 16624 19898 16676
rect 19898 16624 19924 16676
rect 19628 16622 19684 16624
rect 19708 16622 19764 16624
rect 19788 16622 19844 16624
rect 19868 16622 19924 16624
rect 19628 15344 19684 15346
rect 19708 15344 19764 15346
rect 19788 15344 19844 15346
rect 19868 15344 19924 15346
rect 19628 15292 19654 15344
rect 19654 15292 19684 15344
rect 19708 15292 19718 15344
rect 19718 15292 19764 15344
rect 19788 15292 19834 15344
rect 19834 15292 19844 15344
rect 19868 15292 19898 15344
rect 19898 15292 19924 15344
rect 19628 15290 19684 15292
rect 19708 15290 19764 15292
rect 19788 15290 19844 15292
rect 19868 15290 19924 15292
rect 19628 14012 19684 14014
rect 19708 14012 19764 14014
rect 19788 14012 19844 14014
rect 19868 14012 19924 14014
rect 19628 13960 19654 14012
rect 19654 13960 19684 14012
rect 19708 13960 19718 14012
rect 19718 13960 19764 14012
rect 19788 13960 19834 14012
rect 19834 13960 19844 14012
rect 19868 13960 19898 14012
rect 19898 13960 19924 14012
rect 19628 13958 19684 13960
rect 19708 13958 19764 13960
rect 19788 13958 19844 13960
rect 19868 13958 19924 13960
rect 19628 12680 19684 12682
rect 19708 12680 19764 12682
rect 19788 12680 19844 12682
rect 19868 12680 19924 12682
rect 19628 12628 19654 12680
rect 19654 12628 19684 12680
rect 19708 12628 19718 12680
rect 19718 12628 19764 12680
rect 19788 12628 19834 12680
rect 19834 12628 19844 12680
rect 19868 12628 19898 12680
rect 19898 12628 19924 12680
rect 19628 12626 19684 12628
rect 19708 12626 19764 12628
rect 19788 12626 19844 12628
rect 19868 12626 19924 12628
rect 19628 11348 19684 11350
rect 19708 11348 19764 11350
rect 19788 11348 19844 11350
rect 19868 11348 19924 11350
rect 19628 11296 19654 11348
rect 19654 11296 19684 11348
rect 19708 11296 19718 11348
rect 19718 11296 19764 11348
rect 19788 11296 19834 11348
rect 19834 11296 19844 11348
rect 19868 11296 19898 11348
rect 19898 11296 19924 11348
rect 19628 11294 19684 11296
rect 19708 11294 19764 11296
rect 19788 11294 19844 11296
rect 19868 11294 19924 11296
rect 19628 10016 19684 10018
rect 19708 10016 19764 10018
rect 19788 10016 19844 10018
rect 19868 10016 19924 10018
rect 19628 9964 19654 10016
rect 19654 9964 19684 10016
rect 19708 9964 19718 10016
rect 19718 9964 19764 10016
rect 19788 9964 19834 10016
rect 19834 9964 19844 10016
rect 19868 9964 19898 10016
rect 19898 9964 19924 10016
rect 19628 9962 19684 9964
rect 19708 9962 19764 9964
rect 19788 9962 19844 9964
rect 19868 9962 19924 9964
rect 19628 8684 19684 8686
rect 19708 8684 19764 8686
rect 19788 8684 19844 8686
rect 19868 8684 19924 8686
rect 19628 8632 19654 8684
rect 19654 8632 19684 8684
rect 19708 8632 19718 8684
rect 19718 8632 19764 8684
rect 19788 8632 19834 8684
rect 19834 8632 19844 8684
rect 19868 8632 19898 8684
rect 19898 8632 19924 8684
rect 19628 8630 19684 8632
rect 19708 8630 19764 8632
rect 19788 8630 19844 8632
rect 19868 8630 19924 8632
rect 19628 7352 19684 7354
rect 19708 7352 19764 7354
rect 19788 7352 19844 7354
rect 19868 7352 19924 7354
rect 19628 7300 19654 7352
rect 19654 7300 19684 7352
rect 19708 7300 19718 7352
rect 19718 7300 19764 7352
rect 19788 7300 19834 7352
rect 19834 7300 19844 7352
rect 19868 7300 19898 7352
rect 19898 7300 19924 7352
rect 19628 7298 19684 7300
rect 19708 7298 19764 7300
rect 19788 7298 19844 7300
rect 19868 7298 19924 7300
rect 19628 6020 19684 6022
rect 19708 6020 19764 6022
rect 19788 6020 19844 6022
rect 19868 6020 19924 6022
rect 19628 5968 19654 6020
rect 19654 5968 19684 6020
rect 19708 5968 19718 6020
rect 19718 5968 19764 6020
rect 19788 5968 19834 6020
rect 19834 5968 19844 6020
rect 19868 5968 19898 6020
rect 19898 5968 19924 6020
rect 19628 5966 19684 5968
rect 19708 5966 19764 5968
rect 19788 5966 19844 5968
rect 19868 5966 19924 5968
rect 19628 4688 19684 4690
rect 19708 4688 19764 4690
rect 19788 4688 19844 4690
rect 19868 4688 19924 4690
rect 19628 4636 19654 4688
rect 19654 4636 19684 4688
rect 19708 4636 19718 4688
rect 19718 4636 19764 4688
rect 19788 4636 19834 4688
rect 19834 4636 19844 4688
rect 19868 4636 19898 4688
rect 19898 4636 19924 4688
rect 19628 4634 19684 4636
rect 19708 4634 19764 4636
rect 19788 4634 19844 4636
rect 19868 4634 19924 4636
rect 19628 3356 19684 3358
rect 19708 3356 19764 3358
rect 19788 3356 19844 3358
rect 19868 3356 19924 3358
rect 19628 3304 19654 3356
rect 19654 3304 19684 3356
rect 19708 3304 19718 3356
rect 19718 3304 19764 3356
rect 19788 3304 19834 3356
rect 19834 3304 19844 3356
rect 19868 3304 19898 3356
rect 19898 3304 19924 3356
rect 19628 3302 19684 3304
rect 19708 3302 19764 3304
rect 19788 3302 19844 3304
rect 19868 3302 19924 3304
rect 34988 57302 35044 57304
rect 35068 57302 35124 57304
rect 35148 57302 35204 57304
rect 35228 57302 35284 57304
rect 34988 57250 35014 57302
rect 35014 57250 35044 57302
rect 35068 57250 35078 57302
rect 35078 57250 35124 57302
rect 35148 57250 35194 57302
rect 35194 57250 35204 57302
rect 35228 57250 35258 57302
rect 35258 57250 35284 57302
rect 34988 57248 35044 57250
rect 35068 57248 35124 57250
rect 35148 57248 35204 57250
rect 35228 57248 35284 57250
rect 34988 55970 35044 55972
rect 35068 55970 35124 55972
rect 35148 55970 35204 55972
rect 35228 55970 35284 55972
rect 34988 55918 35014 55970
rect 35014 55918 35044 55970
rect 35068 55918 35078 55970
rect 35078 55918 35124 55970
rect 35148 55918 35194 55970
rect 35194 55918 35204 55970
rect 35228 55918 35258 55970
rect 35258 55918 35284 55970
rect 34988 55916 35044 55918
rect 35068 55916 35124 55918
rect 35148 55916 35204 55918
rect 35228 55916 35284 55918
rect 34988 54638 35044 54640
rect 35068 54638 35124 54640
rect 35148 54638 35204 54640
rect 35228 54638 35284 54640
rect 34988 54586 35014 54638
rect 35014 54586 35044 54638
rect 35068 54586 35078 54638
rect 35078 54586 35124 54638
rect 35148 54586 35194 54638
rect 35194 54586 35204 54638
rect 35228 54586 35258 54638
rect 35258 54586 35284 54638
rect 34988 54584 35044 54586
rect 35068 54584 35124 54586
rect 35148 54584 35204 54586
rect 35228 54584 35284 54586
rect 34988 53306 35044 53308
rect 35068 53306 35124 53308
rect 35148 53306 35204 53308
rect 35228 53306 35284 53308
rect 34988 53254 35014 53306
rect 35014 53254 35044 53306
rect 35068 53254 35078 53306
rect 35078 53254 35124 53306
rect 35148 53254 35194 53306
rect 35194 53254 35204 53306
rect 35228 53254 35258 53306
rect 35258 53254 35284 53306
rect 34988 53252 35044 53254
rect 35068 53252 35124 53254
rect 35148 53252 35204 53254
rect 35228 53252 35284 53254
rect 34988 51974 35044 51976
rect 35068 51974 35124 51976
rect 35148 51974 35204 51976
rect 35228 51974 35284 51976
rect 34988 51922 35014 51974
rect 35014 51922 35044 51974
rect 35068 51922 35078 51974
rect 35078 51922 35124 51974
rect 35148 51922 35194 51974
rect 35194 51922 35204 51974
rect 35228 51922 35258 51974
rect 35258 51922 35284 51974
rect 34988 51920 35044 51922
rect 35068 51920 35124 51922
rect 35148 51920 35204 51922
rect 35228 51920 35284 51922
rect 34988 50642 35044 50644
rect 35068 50642 35124 50644
rect 35148 50642 35204 50644
rect 35228 50642 35284 50644
rect 34988 50590 35014 50642
rect 35014 50590 35044 50642
rect 35068 50590 35078 50642
rect 35078 50590 35124 50642
rect 35148 50590 35194 50642
rect 35194 50590 35204 50642
rect 35228 50590 35258 50642
rect 35258 50590 35284 50642
rect 34988 50588 35044 50590
rect 35068 50588 35124 50590
rect 35148 50588 35204 50590
rect 35228 50588 35284 50590
rect 34988 49310 35044 49312
rect 35068 49310 35124 49312
rect 35148 49310 35204 49312
rect 35228 49310 35284 49312
rect 34988 49258 35014 49310
rect 35014 49258 35044 49310
rect 35068 49258 35078 49310
rect 35078 49258 35124 49310
rect 35148 49258 35194 49310
rect 35194 49258 35204 49310
rect 35228 49258 35258 49310
rect 35258 49258 35284 49310
rect 34988 49256 35044 49258
rect 35068 49256 35124 49258
rect 35148 49256 35204 49258
rect 35228 49256 35284 49258
rect 34988 47978 35044 47980
rect 35068 47978 35124 47980
rect 35148 47978 35204 47980
rect 35228 47978 35284 47980
rect 34988 47926 35014 47978
rect 35014 47926 35044 47978
rect 35068 47926 35078 47978
rect 35078 47926 35124 47978
rect 35148 47926 35194 47978
rect 35194 47926 35204 47978
rect 35228 47926 35258 47978
rect 35258 47926 35284 47978
rect 34988 47924 35044 47926
rect 35068 47924 35124 47926
rect 35148 47924 35204 47926
rect 35228 47924 35284 47926
rect 34988 46646 35044 46648
rect 35068 46646 35124 46648
rect 35148 46646 35204 46648
rect 35228 46646 35284 46648
rect 34988 46594 35014 46646
rect 35014 46594 35044 46646
rect 35068 46594 35078 46646
rect 35078 46594 35124 46646
rect 35148 46594 35194 46646
rect 35194 46594 35204 46646
rect 35228 46594 35258 46646
rect 35258 46594 35284 46646
rect 34988 46592 35044 46594
rect 35068 46592 35124 46594
rect 35148 46592 35204 46594
rect 35228 46592 35284 46594
rect 34988 45314 35044 45316
rect 35068 45314 35124 45316
rect 35148 45314 35204 45316
rect 35228 45314 35284 45316
rect 34988 45262 35014 45314
rect 35014 45262 35044 45314
rect 35068 45262 35078 45314
rect 35078 45262 35124 45314
rect 35148 45262 35194 45314
rect 35194 45262 35204 45314
rect 35228 45262 35258 45314
rect 35258 45262 35284 45314
rect 34988 45260 35044 45262
rect 35068 45260 35124 45262
rect 35148 45260 35204 45262
rect 35228 45260 35284 45262
rect 34988 43982 35044 43984
rect 35068 43982 35124 43984
rect 35148 43982 35204 43984
rect 35228 43982 35284 43984
rect 34988 43930 35014 43982
rect 35014 43930 35044 43982
rect 35068 43930 35078 43982
rect 35078 43930 35124 43982
rect 35148 43930 35194 43982
rect 35194 43930 35204 43982
rect 35228 43930 35258 43982
rect 35258 43930 35284 43982
rect 34988 43928 35044 43930
rect 35068 43928 35124 43930
rect 35148 43928 35204 43930
rect 35228 43928 35284 43930
rect 34988 42650 35044 42652
rect 35068 42650 35124 42652
rect 35148 42650 35204 42652
rect 35228 42650 35284 42652
rect 34988 42598 35014 42650
rect 35014 42598 35044 42650
rect 35068 42598 35078 42650
rect 35078 42598 35124 42650
rect 35148 42598 35194 42650
rect 35194 42598 35204 42650
rect 35228 42598 35258 42650
rect 35258 42598 35284 42650
rect 34988 42596 35044 42598
rect 35068 42596 35124 42598
rect 35148 42596 35204 42598
rect 35228 42596 35284 42598
rect 34988 41318 35044 41320
rect 35068 41318 35124 41320
rect 35148 41318 35204 41320
rect 35228 41318 35284 41320
rect 34988 41266 35014 41318
rect 35014 41266 35044 41318
rect 35068 41266 35078 41318
rect 35078 41266 35124 41318
rect 35148 41266 35194 41318
rect 35194 41266 35204 41318
rect 35228 41266 35258 41318
rect 35258 41266 35284 41318
rect 34988 41264 35044 41266
rect 35068 41264 35124 41266
rect 35148 41264 35204 41266
rect 35228 41264 35284 41266
rect 34988 39986 35044 39988
rect 35068 39986 35124 39988
rect 35148 39986 35204 39988
rect 35228 39986 35284 39988
rect 34988 39934 35014 39986
rect 35014 39934 35044 39986
rect 35068 39934 35078 39986
rect 35078 39934 35124 39986
rect 35148 39934 35194 39986
rect 35194 39934 35204 39986
rect 35228 39934 35258 39986
rect 35258 39934 35284 39986
rect 34988 39932 35044 39934
rect 35068 39932 35124 39934
rect 35148 39932 35204 39934
rect 35228 39932 35284 39934
rect 34988 38654 35044 38656
rect 35068 38654 35124 38656
rect 35148 38654 35204 38656
rect 35228 38654 35284 38656
rect 34988 38602 35014 38654
rect 35014 38602 35044 38654
rect 35068 38602 35078 38654
rect 35078 38602 35124 38654
rect 35148 38602 35194 38654
rect 35194 38602 35204 38654
rect 35228 38602 35258 38654
rect 35258 38602 35284 38654
rect 34988 38600 35044 38602
rect 35068 38600 35124 38602
rect 35148 38600 35204 38602
rect 35228 38600 35284 38602
rect 34988 37322 35044 37324
rect 35068 37322 35124 37324
rect 35148 37322 35204 37324
rect 35228 37322 35284 37324
rect 34988 37270 35014 37322
rect 35014 37270 35044 37322
rect 35068 37270 35078 37322
rect 35078 37270 35124 37322
rect 35148 37270 35194 37322
rect 35194 37270 35204 37322
rect 35228 37270 35258 37322
rect 35258 37270 35284 37322
rect 34988 37268 35044 37270
rect 35068 37268 35124 37270
rect 35148 37268 35204 37270
rect 35228 37268 35284 37270
rect 34988 35990 35044 35992
rect 35068 35990 35124 35992
rect 35148 35990 35204 35992
rect 35228 35990 35284 35992
rect 34988 35938 35014 35990
rect 35014 35938 35044 35990
rect 35068 35938 35078 35990
rect 35078 35938 35124 35990
rect 35148 35938 35194 35990
rect 35194 35938 35204 35990
rect 35228 35938 35258 35990
rect 35258 35938 35284 35990
rect 34988 35936 35044 35938
rect 35068 35936 35124 35938
rect 35148 35936 35204 35938
rect 35228 35936 35284 35938
rect 34988 34658 35044 34660
rect 35068 34658 35124 34660
rect 35148 34658 35204 34660
rect 35228 34658 35284 34660
rect 34988 34606 35014 34658
rect 35014 34606 35044 34658
rect 35068 34606 35078 34658
rect 35078 34606 35124 34658
rect 35148 34606 35194 34658
rect 35194 34606 35204 34658
rect 35228 34606 35258 34658
rect 35258 34606 35284 34658
rect 34988 34604 35044 34606
rect 35068 34604 35124 34606
rect 35148 34604 35204 34606
rect 35228 34604 35284 34606
rect 34988 33326 35044 33328
rect 35068 33326 35124 33328
rect 35148 33326 35204 33328
rect 35228 33326 35284 33328
rect 34988 33274 35014 33326
rect 35014 33274 35044 33326
rect 35068 33274 35078 33326
rect 35078 33274 35124 33326
rect 35148 33274 35194 33326
rect 35194 33274 35204 33326
rect 35228 33274 35258 33326
rect 35258 33274 35284 33326
rect 34988 33272 35044 33274
rect 35068 33272 35124 33274
rect 35148 33272 35204 33274
rect 35228 33272 35284 33274
rect 34988 31994 35044 31996
rect 35068 31994 35124 31996
rect 35148 31994 35204 31996
rect 35228 31994 35284 31996
rect 34988 31942 35014 31994
rect 35014 31942 35044 31994
rect 35068 31942 35078 31994
rect 35078 31942 35124 31994
rect 35148 31942 35194 31994
rect 35194 31942 35204 31994
rect 35228 31942 35258 31994
rect 35258 31942 35284 31994
rect 34988 31940 35044 31942
rect 35068 31940 35124 31942
rect 35148 31940 35204 31942
rect 35228 31940 35284 31942
rect 34988 30662 35044 30664
rect 35068 30662 35124 30664
rect 35148 30662 35204 30664
rect 35228 30662 35284 30664
rect 34988 30610 35014 30662
rect 35014 30610 35044 30662
rect 35068 30610 35078 30662
rect 35078 30610 35124 30662
rect 35148 30610 35194 30662
rect 35194 30610 35204 30662
rect 35228 30610 35258 30662
rect 35258 30610 35284 30662
rect 34988 30608 35044 30610
rect 35068 30608 35124 30610
rect 35148 30608 35204 30610
rect 35228 30608 35284 30610
rect 34988 29330 35044 29332
rect 35068 29330 35124 29332
rect 35148 29330 35204 29332
rect 35228 29330 35284 29332
rect 34988 29278 35014 29330
rect 35014 29278 35044 29330
rect 35068 29278 35078 29330
rect 35078 29278 35124 29330
rect 35148 29278 35194 29330
rect 35194 29278 35204 29330
rect 35228 29278 35258 29330
rect 35258 29278 35284 29330
rect 34988 29276 35044 29278
rect 35068 29276 35124 29278
rect 35148 29276 35204 29278
rect 35228 29276 35284 29278
rect 34988 27998 35044 28000
rect 35068 27998 35124 28000
rect 35148 27998 35204 28000
rect 35228 27998 35284 28000
rect 34988 27946 35014 27998
rect 35014 27946 35044 27998
rect 35068 27946 35078 27998
rect 35078 27946 35124 27998
rect 35148 27946 35194 27998
rect 35194 27946 35204 27998
rect 35228 27946 35258 27998
rect 35258 27946 35284 27998
rect 34988 27944 35044 27946
rect 35068 27944 35124 27946
rect 35148 27944 35204 27946
rect 35228 27944 35284 27946
rect 34988 26666 35044 26668
rect 35068 26666 35124 26668
rect 35148 26666 35204 26668
rect 35228 26666 35284 26668
rect 34988 26614 35014 26666
rect 35014 26614 35044 26666
rect 35068 26614 35078 26666
rect 35078 26614 35124 26666
rect 35148 26614 35194 26666
rect 35194 26614 35204 26666
rect 35228 26614 35258 26666
rect 35258 26614 35284 26666
rect 34988 26612 35044 26614
rect 35068 26612 35124 26614
rect 35148 26612 35204 26614
rect 35228 26612 35284 26614
rect 34988 25334 35044 25336
rect 35068 25334 35124 25336
rect 35148 25334 35204 25336
rect 35228 25334 35284 25336
rect 34988 25282 35014 25334
rect 35014 25282 35044 25334
rect 35068 25282 35078 25334
rect 35078 25282 35124 25334
rect 35148 25282 35194 25334
rect 35194 25282 35204 25334
rect 35228 25282 35258 25334
rect 35258 25282 35284 25334
rect 34988 25280 35044 25282
rect 35068 25280 35124 25282
rect 35148 25280 35204 25282
rect 35228 25280 35284 25282
rect 34988 24002 35044 24004
rect 35068 24002 35124 24004
rect 35148 24002 35204 24004
rect 35228 24002 35284 24004
rect 34988 23950 35014 24002
rect 35014 23950 35044 24002
rect 35068 23950 35078 24002
rect 35078 23950 35124 24002
rect 35148 23950 35194 24002
rect 35194 23950 35204 24002
rect 35228 23950 35258 24002
rect 35258 23950 35284 24002
rect 34988 23948 35044 23950
rect 35068 23948 35124 23950
rect 35148 23948 35204 23950
rect 35228 23948 35284 23950
rect 34988 22670 35044 22672
rect 35068 22670 35124 22672
rect 35148 22670 35204 22672
rect 35228 22670 35284 22672
rect 34988 22618 35014 22670
rect 35014 22618 35044 22670
rect 35068 22618 35078 22670
rect 35078 22618 35124 22670
rect 35148 22618 35194 22670
rect 35194 22618 35204 22670
rect 35228 22618 35258 22670
rect 35258 22618 35284 22670
rect 34988 22616 35044 22618
rect 35068 22616 35124 22618
rect 35148 22616 35204 22618
rect 35228 22616 35284 22618
rect 34988 21338 35044 21340
rect 35068 21338 35124 21340
rect 35148 21338 35204 21340
rect 35228 21338 35284 21340
rect 34988 21286 35014 21338
rect 35014 21286 35044 21338
rect 35068 21286 35078 21338
rect 35078 21286 35124 21338
rect 35148 21286 35194 21338
rect 35194 21286 35204 21338
rect 35228 21286 35258 21338
rect 35258 21286 35284 21338
rect 34988 21284 35044 21286
rect 35068 21284 35124 21286
rect 35148 21284 35204 21286
rect 35228 21284 35284 21286
rect 34988 20006 35044 20008
rect 35068 20006 35124 20008
rect 35148 20006 35204 20008
rect 35228 20006 35284 20008
rect 34988 19954 35014 20006
rect 35014 19954 35044 20006
rect 35068 19954 35078 20006
rect 35078 19954 35124 20006
rect 35148 19954 35194 20006
rect 35194 19954 35204 20006
rect 35228 19954 35258 20006
rect 35258 19954 35284 20006
rect 34988 19952 35044 19954
rect 35068 19952 35124 19954
rect 35148 19952 35204 19954
rect 35228 19952 35284 19954
rect 34988 18674 35044 18676
rect 35068 18674 35124 18676
rect 35148 18674 35204 18676
rect 35228 18674 35284 18676
rect 34988 18622 35014 18674
rect 35014 18622 35044 18674
rect 35068 18622 35078 18674
rect 35078 18622 35124 18674
rect 35148 18622 35194 18674
rect 35194 18622 35204 18674
rect 35228 18622 35258 18674
rect 35258 18622 35284 18674
rect 34988 18620 35044 18622
rect 35068 18620 35124 18622
rect 35148 18620 35204 18622
rect 35228 18620 35284 18622
rect 34988 17342 35044 17344
rect 35068 17342 35124 17344
rect 35148 17342 35204 17344
rect 35228 17342 35284 17344
rect 34988 17290 35014 17342
rect 35014 17290 35044 17342
rect 35068 17290 35078 17342
rect 35078 17290 35124 17342
rect 35148 17290 35194 17342
rect 35194 17290 35204 17342
rect 35228 17290 35258 17342
rect 35258 17290 35284 17342
rect 34988 17288 35044 17290
rect 35068 17288 35124 17290
rect 35148 17288 35204 17290
rect 35228 17288 35284 17290
rect 34988 16010 35044 16012
rect 35068 16010 35124 16012
rect 35148 16010 35204 16012
rect 35228 16010 35284 16012
rect 34988 15958 35014 16010
rect 35014 15958 35044 16010
rect 35068 15958 35078 16010
rect 35078 15958 35124 16010
rect 35148 15958 35194 16010
rect 35194 15958 35204 16010
rect 35228 15958 35258 16010
rect 35258 15958 35284 16010
rect 34988 15956 35044 15958
rect 35068 15956 35124 15958
rect 35148 15956 35204 15958
rect 35228 15956 35284 15958
rect 34988 14678 35044 14680
rect 35068 14678 35124 14680
rect 35148 14678 35204 14680
rect 35228 14678 35284 14680
rect 34988 14626 35014 14678
rect 35014 14626 35044 14678
rect 35068 14626 35078 14678
rect 35078 14626 35124 14678
rect 35148 14626 35194 14678
rect 35194 14626 35204 14678
rect 35228 14626 35258 14678
rect 35258 14626 35284 14678
rect 34988 14624 35044 14626
rect 35068 14624 35124 14626
rect 35148 14624 35204 14626
rect 35228 14624 35284 14626
rect 34988 13346 35044 13348
rect 35068 13346 35124 13348
rect 35148 13346 35204 13348
rect 35228 13346 35284 13348
rect 34988 13294 35014 13346
rect 35014 13294 35044 13346
rect 35068 13294 35078 13346
rect 35078 13294 35124 13346
rect 35148 13294 35194 13346
rect 35194 13294 35204 13346
rect 35228 13294 35258 13346
rect 35258 13294 35284 13346
rect 34988 13292 35044 13294
rect 35068 13292 35124 13294
rect 35148 13292 35204 13294
rect 35228 13292 35284 13294
rect 34988 12014 35044 12016
rect 35068 12014 35124 12016
rect 35148 12014 35204 12016
rect 35228 12014 35284 12016
rect 34988 11962 35014 12014
rect 35014 11962 35044 12014
rect 35068 11962 35078 12014
rect 35078 11962 35124 12014
rect 35148 11962 35194 12014
rect 35194 11962 35204 12014
rect 35228 11962 35258 12014
rect 35258 11962 35284 12014
rect 34988 11960 35044 11962
rect 35068 11960 35124 11962
rect 35148 11960 35204 11962
rect 35228 11960 35284 11962
rect 34988 10682 35044 10684
rect 35068 10682 35124 10684
rect 35148 10682 35204 10684
rect 35228 10682 35284 10684
rect 34988 10630 35014 10682
rect 35014 10630 35044 10682
rect 35068 10630 35078 10682
rect 35078 10630 35124 10682
rect 35148 10630 35194 10682
rect 35194 10630 35204 10682
rect 35228 10630 35258 10682
rect 35258 10630 35284 10682
rect 34988 10628 35044 10630
rect 35068 10628 35124 10630
rect 35148 10628 35204 10630
rect 35228 10628 35284 10630
rect 34988 9350 35044 9352
rect 35068 9350 35124 9352
rect 35148 9350 35204 9352
rect 35228 9350 35284 9352
rect 34988 9298 35014 9350
rect 35014 9298 35044 9350
rect 35068 9298 35078 9350
rect 35078 9298 35124 9350
rect 35148 9298 35194 9350
rect 35194 9298 35204 9350
rect 35228 9298 35258 9350
rect 35258 9298 35284 9350
rect 34988 9296 35044 9298
rect 35068 9296 35124 9298
rect 35148 9296 35204 9298
rect 35228 9296 35284 9298
rect 34988 8018 35044 8020
rect 35068 8018 35124 8020
rect 35148 8018 35204 8020
rect 35228 8018 35284 8020
rect 34988 7966 35014 8018
rect 35014 7966 35044 8018
rect 35068 7966 35078 8018
rect 35078 7966 35124 8018
rect 35148 7966 35194 8018
rect 35194 7966 35204 8018
rect 35228 7966 35258 8018
rect 35258 7966 35284 8018
rect 34988 7964 35044 7966
rect 35068 7964 35124 7966
rect 35148 7964 35204 7966
rect 35228 7964 35284 7966
rect 34988 6686 35044 6688
rect 35068 6686 35124 6688
rect 35148 6686 35204 6688
rect 35228 6686 35284 6688
rect 34988 6634 35014 6686
rect 35014 6634 35044 6686
rect 35068 6634 35078 6686
rect 35078 6634 35124 6686
rect 35148 6634 35194 6686
rect 35194 6634 35204 6686
rect 35228 6634 35258 6686
rect 35258 6634 35284 6686
rect 34988 6632 35044 6634
rect 35068 6632 35124 6634
rect 35148 6632 35204 6634
rect 35228 6632 35284 6634
rect 34988 5354 35044 5356
rect 35068 5354 35124 5356
rect 35148 5354 35204 5356
rect 35228 5354 35284 5356
rect 34988 5302 35014 5354
rect 35014 5302 35044 5354
rect 35068 5302 35078 5354
rect 35078 5302 35124 5354
rect 35148 5302 35194 5354
rect 35194 5302 35204 5354
rect 35228 5302 35258 5354
rect 35258 5302 35284 5354
rect 34988 5300 35044 5302
rect 35068 5300 35124 5302
rect 35148 5300 35204 5302
rect 35228 5300 35284 5302
rect 34988 4022 35044 4024
rect 35068 4022 35124 4024
rect 35148 4022 35204 4024
rect 35228 4022 35284 4024
rect 34988 3970 35014 4022
rect 35014 3970 35044 4022
rect 35068 3970 35078 4022
rect 35078 3970 35124 4022
rect 35148 3970 35194 4022
rect 35194 3970 35204 4022
rect 35228 3970 35258 4022
rect 35258 3970 35284 4022
rect 34988 3968 35044 3970
rect 35068 3968 35124 3970
rect 35148 3968 35204 3970
rect 35228 3968 35284 3970
rect 34988 2690 35044 2692
rect 35068 2690 35124 2692
rect 35148 2690 35204 2692
rect 35228 2690 35284 2692
rect 34988 2638 35014 2690
rect 35014 2638 35044 2690
rect 35068 2638 35078 2690
rect 35078 2638 35124 2690
rect 35148 2638 35194 2690
rect 35194 2638 35204 2690
rect 35228 2638 35258 2690
rect 35258 2638 35284 2690
rect 34988 2636 35044 2638
rect 35068 2636 35124 2638
rect 35148 2636 35204 2638
rect 35228 2636 35284 2638
rect 50348 56636 50404 56638
rect 50428 56636 50484 56638
rect 50508 56636 50564 56638
rect 50588 56636 50644 56638
rect 50348 56584 50374 56636
rect 50374 56584 50404 56636
rect 50428 56584 50438 56636
rect 50438 56584 50484 56636
rect 50508 56584 50554 56636
rect 50554 56584 50564 56636
rect 50588 56584 50618 56636
rect 50618 56584 50644 56636
rect 50348 56582 50404 56584
rect 50428 56582 50484 56584
rect 50508 56582 50564 56584
rect 50588 56582 50644 56584
rect 50348 55304 50404 55306
rect 50428 55304 50484 55306
rect 50508 55304 50564 55306
rect 50588 55304 50644 55306
rect 50348 55252 50374 55304
rect 50374 55252 50404 55304
rect 50428 55252 50438 55304
rect 50438 55252 50484 55304
rect 50508 55252 50554 55304
rect 50554 55252 50564 55304
rect 50588 55252 50618 55304
rect 50618 55252 50644 55304
rect 50348 55250 50404 55252
rect 50428 55250 50484 55252
rect 50508 55250 50564 55252
rect 50588 55250 50644 55252
rect 50348 53972 50404 53974
rect 50428 53972 50484 53974
rect 50508 53972 50564 53974
rect 50588 53972 50644 53974
rect 50348 53920 50374 53972
rect 50374 53920 50404 53972
rect 50428 53920 50438 53972
rect 50438 53920 50484 53972
rect 50508 53920 50554 53972
rect 50554 53920 50564 53972
rect 50588 53920 50618 53972
rect 50618 53920 50644 53972
rect 50348 53918 50404 53920
rect 50428 53918 50484 53920
rect 50508 53918 50564 53920
rect 50588 53918 50644 53920
rect 50348 52640 50404 52642
rect 50428 52640 50484 52642
rect 50508 52640 50564 52642
rect 50588 52640 50644 52642
rect 50348 52588 50374 52640
rect 50374 52588 50404 52640
rect 50428 52588 50438 52640
rect 50438 52588 50484 52640
rect 50508 52588 50554 52640
rect 50554 52588 50564 52640
rect 50588 52588 50618 52640
rect 50618 52588 50644 52640
rect 50348 52586 50404 52588
rect 50428 52586 50484 52588
rect 50508 52586 50564 52588
rect 50588 52586 50644 52588
rect 50348 51308 50404 51310
rect 50428 51308 50484 51310
rect 50508 51308 50564 51310
rect 50588 51308 50644 51310
rect 50348 51256 50374 51308
rect 50374 51256 50404 51308
rect 50428 51256 50438 51308
rect 50438 51256 50484 51308
rect 50508 51256 50554 51308
rect 50554 51256 50564 51308
rect 50588 51256 50618 51308
rect 50618 51256 50644 51308
rect 50348 51254 50404 51256
rect 50428 51254 50484 51256
rect 50508 51254 50564 51256
rect 50588 51254 50644 51256
rect 50348 49976 50404 49978
rect 50428 49976 50484 49978
rect 50508 49976 50564 49978
rect 50588 49976 50644 49978
rect 50348 49924 50374 49976
rect 50374 49924 50404 49976
rect 50428 49924 50438 49976
rect 50438 49924 50484 49976
rect 50508 49924 50554 49976
rect 50554 49924 50564 49976
rect 50588 49924 50618 49976
rect 50618 49924 50644 49976
rect 50348 49922 50404 49924
rect 50428 49922 50484 49924
rect 50508 49922 50564 49924
rect 50588 49922 50644 49924
rect 50348 48644 50404 48646
rect 50428 48644 50484 48646
rect 50508 48644 50564 48646
rect 50588 48644 50644 48646
rect 50348 48592 50374 48644
rect 50374 48592 50404 48644
rect 50428 48592 50438 48644
rect 50438 48592 50484 48644
rect 50508 48592 50554 48644
rect 50554 48592 50564 48644
rect 50588 48592 50618 48644
rect 50618 48592 50644 48644
rect 50348 48590 50404 48592
rect 50428 48590 50484 48592
rect 50508 48590 50564 48592
rect 50588 48590 50644 48592
rect 50348 47312 50404 47314
rect 50428 47312 50484 47314
rect 50508 47312 50564 47314
rect 50588 47312 50644 47314
rect 50348 47260 50374 47312
rect 50374 47260 50404 47312
rect 50428 47260 50438 47312
rect 50438 47260 50484 47312
rect 50508 47260 50554 47312
rect 50554 47260 50564 47312
rect 50588 47260 50618 47312
rect 50618 47260 50644 47312
rect 50348 47258 50404 47260
rect 50428 47258 50484 47260
rect 50508 47258 50564 47260
rect 50588 47258 50644 47260
rect 50348 45980 50404 45982
rect 50428 45980 50484 45982
rect 50508 45980 50564 45982
rect 50588 45980 50644 45982
rect 50348 45928 50374 45980
rect 50374 45928 50404 45980
rect 50428 45928 50438 45980
rect 50438 45928 50484 45980
rect 50508 45928 50554 45980
rect 50554 45928 50564 45980
rect 50588 45928 50618 45980
rect 50618 45928 50644 45980
rect 50348 45926 50404 45928
rect 50428 45926 50484 45928
rect 50508 45926 50564 45928
rect 50588 45926 50644 45928
rect 50348 44648 50404 44650
rect 50428 44648 50484 44650
rect 50508 44648 50564 44650
rect 50588 44648 50644 44650
rect 50348 44596 50374 44648
rect 50374 44596 50404 44648
rect 50428 44596 50438 44648
rect 50438 44596 50484 44648
rect 50508 44596 50554 44648
rect 50554 44596 50564 44648
rect 50588 44596 50618 44648
rect 50618 44596 50644 44648
rect 50348 44594 50404 44596
rect 50428 44594 50484 44596
rect 50508 44594 50564 44596
rect 50588 44594 50644 44596
rect 50348 43316 50404 43318
rect 50428 43316 50484 43318
rect 50508 43316 50564 43318
rect 50588 43316 50644 43318
rect 50348 43264 50374 43316
rect 50374 43264 50404 43316
rect 50428 43264 50438 43316
rect 50438 43264 50484 43316
rect 50508 43264 50554 43316
rect 50554 43264 50564 43316
rect 50588 43264 50618 43316
rect 50618 43264 50644 43316
rect 50348 43262 50404 43264
rect 50428 43262 50484 43264
rect 50508 43262 50564 43264
rect 50588 43262 50644 43264
rect 50348 41984 50404 41986
rect 50428 41984 50484 41986
rect 50508 41984 50564 41986
rect 50588 41984 50644 41986
rect 50348 41932 50374 41984
rect 50374 41932 50404 41984
rect 50428 41932 50438 41984
rect 50438 41932 50484 41984
rect 50508 41932 50554 41984
rect 50554 41932 50564 41984
rect 50588 41932 50618 41984
rect 50618 41932 50644 41984
rect 50348 41930 50404 41932
rect 50428 41930 50484 41932
rect 50508 41930 50564 41932
rect 50588 41930 50644 41932
rect 50348 40652 50404 40654
rect 50428 40652 50484 40654
rect 50508 40652 50564 40654
rect 50588 40652 50644 40654
rect 50348 40600 50374 40652
rect 50374 40600 50404 40652
rect 50428 40600 50438 40652
rect 50438 40600 50484 40652
rect 50508 40600 50554 40652
rect 50554 40600 50564 40652
rect 50588 40600 50618 40652
rect 50618 40600 50644 40652
rect 50348 40598 50404 40600
rect 50428 40598 50484 40600
rect 50508 40598 50564 40600
rect 50588 40598 50644 40600
rect 50348 39320 50404 39322
rect 50428 39320 50484 39322
rect 50508 39320 50564 39322
rect 50588 39320 50644 39322
rect 50348 39268 50374 39320
rect 50374 39268 50404 39320
rect 50428 39268 50438 39320
rect 50438 39268 50484 39320
rect 50508 39268 50554 39320
rect 50554 39268 50564 39320
rect 50588 39268 50618 39320
rect 50618 39268 50644 39320
rect 50348 39266 50404 39268
rect 50428 39266 50484 39268
rect 50508 39266 50564 39268
rect 50588 39266 50644 39268
rect 50348 37988 50404 37990
rect 50428 37988 50484 37990
rect 50508 37988 50564 37990
rect 50588 37988 50644 37990
rect 50348 37936 50374 37988
rect 50374 37936 50404 37988
rect 50428 37936 50438 37988
rect 50438 37936 50484 37988
rect 50508 37936 50554 37988
rect 50554 37936 50564 37988
rect 50588 37936 50618 37988
rect 50618 37936 50644 37988
rect 50348 37934 50404 37936
rect 50428 37934 50484 37936
rect 50508 37934 50564 37936
rect 50588 37934 50644 37936
rect 50348 36656 50404 36658
rect 50428 36656 50484 36658
rect 50508 36656 50564 36658
rect 50588 36656 50644 36658
rect 50348 36604 50374 36656
rect 50374 36604 50404 36656
rect 50428 36604 50438 36656
rect 50438 36604 50484 36656
rect 50508 36604 50554 36656
rect 50554 36604 50564 36656
rect 50588 36604 50618 36656
rect 50618 36604 50644 36656
rect 50348 36602 50404 36604
rect 50428 36602 50484 36604
rect 50508 36602 50564 36604
rect 50588 36602 50644 36604
rect 50348 35324 50404 35326
rect 50428 35324 50484 35326
rect 50508 35324 50564 35326
rect 50588 35324 50644 35326
rect 50348 35272 50374 35324
rect 50374 35272 50404 35324
rect 50428 35272 50438 35324
rect 50438 35272 50484 35324
rect 50508 35272 50554 35324
rect 50554 35272 50564 35324
rect 50588 35272 50618 35324
rect 50618 35272 50644 35324
rect 50348 35270 50404 35272
rect 50428 35270 50484 35272
rect 50508 35270 50564 35272
rect 50588 35270 50644 35272
rect 50348 33992 50404 33994
rect 50428 33992 50484 33994
rect 50508 33992 50564 33994
rect 50588 33992 50644 33994
rect 50348 33940 50374 33992
rect 50374 33940 50404 33992
rect 50428 33940 50438 33992
rect 50438 33940 50484 33992
rect 50508 33940 50554 33992
rect 50554 33940 50564 33992
rect 50588 33940 50618 33992
rect 50618 33940 50644 33992
rect 50348 33938 50404 33940
rect 50428 33938 50484 33940
rect 50508 33938 50564 33940
rect 50588 33938 50644 33940
rect 50348 32660 50404 32662
rect 50428 32660 50484 32662
rect 50508 32660 50564 32662
rect 50588 32660 50644 32662
rect 50348 32608 50374 32660
rect 50374 32608 50404 32660
rect 50428 32608 50438 32660
rect 50438 32608 50484 32660
rect 50508 32608 50554 32660
rect 50554 32608 50564 32660
rect 50588 32608 50618 32660
rect 50618 32608 50644 32660
rect 50348 32606 50404 32608
rect 50428 32606 50484 32608
rect 50508 32606 50564 32608
rect 50588 32606 50644 32608
rect 50348 31328 50404 31330
rect 50428 31328 50484 31330
rect 50508 31328 50564 31330
rect 50588 31328 50644 31330
rect 50348 31276 50374 31328
rect 50374 31276 50404 31328
rect 50428 31276 50438 31328
rect 50438 31276 50484 31328
rect 50508 31276 50554 31328
rect 50554 31276 50564 31328
rect 50588 31276 50618 31328
rect 50618 31276 50644 31328
rect 50348 31274 50404 31276
rect 50428 31274 50484 31276
rect 50508 31274 50564 31276
rect 50588 31274 50644 31276
rect 50348 29996 50404 29998
rect 50428 29996 50484 29998
rect 50508 29996 50564 29998
rect 50588 29996 50644 29998
rect 50348 29944 50374 29996
rect 50374 29944 50404 29996
rect 50428 29944 50438 29996
rect 50438 29944 50484 29996
rect 50508 29944 50554 29996
rect 50554 29944 50564 29996
rect 50588 29944 50618 29996
rect 50618 29944 50644 29996
rect 50348 29942 50404 29944
rect 50428 29942 50484 29944
rect 50508 29942 50564 29944
rect 50588 29942 50644 29944
rect 50348 28664 50404 28666
rect 50428 28664 50484 28666
rect 50508 28664 50564 28666
rect 50588 28664 50644 28666
rect 50348 28612 50374 28664
rect 50374 28612 50404 28664
rect 50428 28612 50438 28664
rect 50438 28612 50484 28664
rect 50508 28612 50554 28664
rect 50554 28612 50564 28664
rect 50588 28612 50618 28664
rect 50618 28612 50644 28664
rect 50348 28610 50404 28612
rect 50428 28610 50484 28612
rect 50508 28610 50564 28612
rect 50588 28610 50644 28612
rect 50348 27332 50404 27334
rect 50428 27332 50484 27334
rect 50508 27332 50564 27334
rect 50588 27332 50644 27334
rect 50348 27280 50374 27332
rect 50374 27280 50404 27332
rect 50428 27280 50438 27332
rect 50438 27280 50484 27332
rect 50508 27280 50554 27332
rect 50554 27280 50564 27332
rect 50588 27280 50618 27332
rect 50618 27280 50644 27332
rect 50348 27278 50404 27280
rect 50428 27278 50484 27280
rect 50508 27278 50564 27280
rect 50588 27278 50644 27280
rect 50348 26000 50404 26002
rect 50428 26000 50484 26002
rect 50508 26000 50564 26002
rect 50588 26000 50644 26002
rect 50348 25948 50374 26000
rect 50374 25948 50404 26000
rect 50428 25948 50438 26000
rect 50438 25948 50484 26000
rect 50508 25948 50554 26000
rect 50554 25948 50564 26000
rect 50588 25948 50618 26000
rect 50618 25948 50644 26000
rect 50348 25946 50404 25948
rect 50428 25946 50484 25948
rect 50508 25946 50564 25948
rect 50588 25946 50644 25948
rect 50348 24668 50404 24670
rect 50428 24668 50484 24670
rect 50508 24668 50564 24670
rect 50588 24668 50644 24670
rect 50348 24616 50374 24668
rect 50374 24616 50404 24668
rect 50428 24616 50438 24668
rect 50438 24616 50484 24668
rect 50508 24616 50554 24668
rect 50554 24616 50564 24668
rect 50588 24616 50618 24668
rect 50618 24616 50644 24668
rect 50348 24614 50404 24616
rect 50428 24614 50484 24616
rect 50508 24614 50564 24616
rect 50588 24614 50644 24616
rect 50348 23336 50404 23338
rect 50428 23336 50484 23338
rect 50508 23336 50564 23338
rect 50588 23336 50644 23338
rect 50348 23284 50374 23336
rect 50374 23284 50404 23336
rect 50428 23284 50438 23336
rect 50438 23284 50484 23336
rect 50508 23284 50554 23336
rect 50554 23284 50564 23336
rect 50588 23284 50618 23336
rect 50618 23284 50644 23336
rect 50348 23282 50404 23284
rect 50428 23282 50484 23284
rect 50508 23282 50564 23284
rect 50588 23282 50644 23284
rect 50348 22004 50404 22006
rect 50428 22004 50484 22006
rect 50508 22004 50564 22006
rect 50588 22004 50644 22006
rect 50348 21952 50374 22004
rect 50374 21952 50404 22004
rect 50428 21952 50438 22004
rect 50438 21952 50484 22004
rect 50508 21952 50554 22004
rect 50554 21952 50564 22004
rect 50588 21952 50618 22004
rect 50618 21952 50644 22004
rect 50348 21950 50404 21952
rect 50428 21950 50484 21952
rect 50508 21950 50564 21952
rect 50588 21950 50644 21952
rect 50348 20672 50404 20674
rect 50428 20672 50484 20674
rect 50508 20672 50564 20674
rect 50588 20672 50644 20674
rect 50348 20620 50374 20672
rect 50374 20620 50404 20672
rect 50428 20620 50438 20672
rect 50438 20620 50484 20672
rect 50508 20620 50554 20672
rect 50554 20620 50564 20672
rect 50588 20620 50618 20672
rect 50618 20620 50644 20672
rect 50348 20618 50404 20620
rect 50428 20618 50484 20620
rect 50508 20618 50564 20620
rect 50588 20618 50644 20620
rect 50348 19340 50404 19342
rect 50428 19340 50484 19342
rect 50508 19340 50564 19342
rect 50588 19340 50644 19342
rect 50348 19288 50374 19340
rect 50374 19288 50404 19340
rect 50428 19288 50438 19340
rect 50438 19288 50484 19340
rect 50508 19288 50554 19340
rect 50554 19288 50564 19340
rect 50588 19288 50618 19340
rect 50618 19288 50644 19340
rect 50348 19286 50404 19288
rect 50428 19286 50484 19288
rect 50508 19286 50564 19288
rect 50588 19286 50644 19288
rect 50348 18008 50404 18010
rect 50428 18008 50484 18010
rect 50508 18008 50564 18010
rect 50588 18008 50644 18010
rect 50348 17956 50374 18008
rect 50374 17956 50404 18008
rect 50428 17956 50438 18008
rect 50438 17956 50484 18008
rect 50508 17956 50554 18008
rect 50554 17956 50564 18008
rect 50588 17956 50618 18008
rect 50618 17956 50644 18008
rect 50348 17954 50404 17956
rect 50428 17954 50484 17956
rect 50508 17954 50564 17956
rect 50588 17954 50644 17956
rect 50348 16676 50404 16678
rect 50428 16676 50484 16678
rect 50508 16676 50564 16678
rect 50588 16676 50644 16678
rect 50348 16624 50374 16676
rect 50374 16624 50404 16676
rect 50428 16624 50438 16676
rect 50438 16624 50484 16676
rect 50508 16624 50554 16676
rect 50554 16624 50564 16676
rect 50588 16624 50618 16676
rect 50618 16624 50644 16676
rect 50348 16622 50404 16624
rect 50428 16622 50484 16624
rect 50508 16622 50564 16624
rect 50588 16622 50644 16624
rect 50348 15344 50404 15346
rect 50428 15344 50484 15346
rect 50508 15344 50564 15346
rect 50588 15344 50644 15346
rect 50348 15292 50374 15344
rect 50374 15292 50404 15344
rect 50428 15292 50438 15344
rect 50438 15292 50484 15344
rect 50508 15292 50554 15344
rect 50554 15292 50564 15344
rect 50588 15292 50618 15344
rect 50618 15292 50644 15344
rect 50348 15290 50404 15292
rect 50428 15290 50484 15292
rect 50508 15290 50564 15292
rect 50588 15290 50644 15292
rect 50348 14012 50404 14014
rect 50428 14012 50484 14014
rect 50508 14012 50564 14014
rect 50588 14012 50644 14014
rect 50348 13960 50374 14012
rect 50374 13960 50404 14012
rect 50428 13960 50438 14012
rect 50438 13960 50484 14012
rect 50508 13960 50554 14012
rect 50554 13960 50564 14012
rect 50588 13960 50618 14012
rect 50618 13960 50644 14012
rect 50348 13958 50404 13960
rect 50428 13958 50484 13960
rect 50508 13958 50564 13960
rect 50588 13958 50644 13960
rect 50348 12680 50404 12682
rect 50428 12680 50484 12682
rect 50508 12680 50564 12682
rect 50588 12680 50644 12682
rect 50348 12628 50374 12680
rect 50374 12628 50404 12680
rect 50428 12628 50438 12680
rect 50438 12628 50484 12680
rect 50508 12628 50554 12680
rect 50554 12628 50564 12680
rect 50588 12628 50618 12680
rect 50618 12628 50644 12680
rect 50348 12626 50404 12628
rect 50428 12626 50484 12628
rect 50508 12626 50564 12628
rect 50588 12626 50644 12628
rect 50348 11348 50404 11350
rect 50428 11348 50484 11350
rect 50508 11348 50564 11350
rect 50588 11348 50644 11350
rect 50348 11296 50374 11348
rect 50374 11296 50404 11348
rect 50428 11296 50438 11348
rect 50438 11296 50484 11348
rect 50508 11296 50554 11348
rect 50554 11296 50564 11348
rect 50588 11296 50618 11348
rect 50618 11296 50644 11348
rect 50348 11294 50404 11296
rect 50428 11294 50484 11296
rect 50508 11294 50564 11296
rect 50588 11294 50644 11296
rect 50348 10016 50404 10018
rect 50428 10016 50484 10018
rect 50508 10016 50564 10018
rect 50588 10016 50644 10018
rect 50348 9964 50374 10016
rect 50374 9964 50404 10016
rect 50428 9964 50438 10016
rect 50438 9964 50484 10016
rect 50508 9964 50554 10016
rect 50554 9964 50564 10016
rect 50588 9964 50618 10016
rect 50618 9964 50644 10016
rect 50348 9962 50404 9964
rect 50428 9962 50484 9964
rect 50508 9962 50564 9964
rect 50588 9962 50644 9964
rect 50348 8684 50404 8686
rect 50428 8684 50484 8686
rect 50508 8684 50564 8686
rect 50588 8684 50644 8686
rect 50348 8632 50374 8684
rect 50374 8632 50404 8684
rect 50428 8632 50438 8684
rect 50438 8632 50484 8684
rect 50508 8632 50554 8684
rect 50554 8632 50564 8684
rect 50588 8632 50618 8684
rect 50618 8632 50644 8684
rect 50348 8630 50404 8632
rect 50428 8630 50484 8632
rect 50508 8630 50564 8632
rect 50588 8630 50644 8632
rect 50348 7352 50404 7354
rect 50428 7352 50484 7354
rect 50508 7352 50564 7354
rect 50588 7352 50644 7354
rect 50348 7300 50374 7352
rect 50374 7300 50404 7352
rect 50428 7300 50438 7352
rect 50438 7300 50484 7352
rect 50508 7300 50554 7352
rect 50554 7300 50564 7352
rect 50588 7300 50618 7352
rect 50618 7300 50644 7352
rect 50348 7298 50404 7300
rect 50428 7298 50484 7300
rect 50508 7298 50564 7300
rect 50588 7298 50644 7300
rect 50348 6020 50404 6022
rect 50428 6020 50484 6022
rect 50508 6020 50564 6022
rect 50588 6020 50644 6022
rect 50348 5968 50374 6020
rect 50374 5968 50404 6020
rect 50428 5968 50438 6020
rect 50438 5968 50484 6020
rect 50508 5968 50554 6020
rect 50554 5968 50564 6020
rect 50588 5968 50618 6020
rect 50618 5968 50644 6020
rect 50348 5966 50404 5968
rect 50428 5966 50484 5968
rect 50508 5966 50564 5968
rect 50588 5966 50644 5968
rect 50348 4688 50404 4690
rect 50428 4688 50484 4690
rect 50508 4688 50564 4690
rect 50588 4688 50644 4690
rect 50348 4636 50374 4688
rect 50374 4636 50404 4688
rect 50428 4636 50438 4688
rect 50438 4636 50484 4688
rect 50508 4636 50554 4688
rect 50554 4636 50564 4688
rect 50588 4636 50618 4688
rect 50618 4636 50644 4688
rect 50348 4634 50404 4636
rect 50428 4634 50484 4636
rect 50508 4634 50564 4636
rect 50588 4634 50644 4636
rect 50348 3356 50404 3358
rect 50428 3356 50484 3358
rect 50508 3356 50564 3358
rect 50588 3356 50644 3358
rect 50348 3304 50374 3356
rect 50374 3304 50404 3356
rect 50428 3304 50438 3356
rect 50438 3304 50484 3356
rect 50508 3304 50554 3356
rect 50554 3304 50564 3356
rect 50588 3304 50618 3356
rect 50618 3304 50644 3356
rect 50348 3302 50404 3304
rect 50428 3302 50484 3304
rect 50508 3302 50564 3304
rect 50588 3302 50644 3304
<< metal3 >>
rect 4256 57308 4576 57309
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 57243 4576 57244
rect 34976 57308 35296 57309
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 57243 35296 57244
rect 19616 56642 19936 56643
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 56577 19936 56578
rect 50336 56642 50656 56643
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 56577 50656 56578
rect 4256 55976 4576 55977
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 55911 4576 55912
rect 34976 55976 35296 55977
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 55911 35296 55912
rect 19616 55310 19936 55311
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 55245 19936 55246
rect 50336 55310 50656 55311
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 55245 50656 55246
rect 4256 54644 4576 54645
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 54579 4576 54580
rect 34976 54644 35296 54645
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 54579 35296 54580
rect 19616 53978 19936 53979
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 53913 19936 53914
rect 50336 53978 50656 53979
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 53913 50656 53914
rect 4256 53312 4576 53313
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 53247 4576 53248
rect 34976 53312 35296 53313
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 53247 35296 53248
rect 19616 52646 19936 52647
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 52581 19936 52582
rect 50336 52646 50656 52647
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 52581 50656 52582
rect 4256 51980 4576 51981
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 51915 4576 51916
rect 34976 51980 35296 51981
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 51915 35296 51916
rect 19616 51314 19936 51315
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 51249 19936 51250
rect 50336 51314 50656 51315
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 51249 50656 51250
rect 4256 50648 4576 50649
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 50583 4576 50584
rect 34976 50648 35296 50649
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 50583 35296 50584
rect 19616 49982 19936 49983
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 49917 19936 49918
rect 50336 49982 50656 49983
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 49917 50656 49918
rect 4256 49316 4576 49317
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 49251 4576 49252
rect 34976 49316 35296 49317
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 49251 35296 49252
rect 19616 48650 19936 48651
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 48585 19936 48586
rect 50336 48650 50656 48651
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 48585 50656 48586
rect 4256 47984 4576 47985
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 47919 4576 47920
rect 34976 47984 35296 47985
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 47919 35296 47920
rect 19616 47318 19936 47319
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 47253 19936 47254
rect 50336 47318 50656 47319
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 47253 50656 47254
rect 4256 46652 4576 46653
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 46587 4576 46588
rect 34976 46652 35296 46653
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 46587 35296 46588
rect 19616 45986 19936 45987
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 45921 19936 45922
rect 50336 45986 50656 45987
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 45921 50656 45922
rect 4256 45320 4576 45321
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 45255 4576 45256
rect 34976 45320 35296 45321
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 45255 35296 45256
rect 19616 44654 19936 44655
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 44589 19936 44590
rect 50336 44654 50656 44655
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 44589 50656 44590
rect 4256 43988 4576 43989
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 43923 4576 43924
rect 34976 43988 35296 43989
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 43923 35296 43924
rect 19616 43322 19936 43323
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 43257 19936 43258
rect 50336 43322 50656 43323
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 43257 50656 43258
rect 4256 42656 4576 42657
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 42591 4576 42592
rect 34976 42656 35296 42657
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 42591 35296 42592
rect 19616 41990 19936 41991
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 41925 19936 41926
rect 50336 41990 50656 41991
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 41925 50656 41926
rect 4256 41324 4576 41325
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 41259 4576 41260
rect 34976 41324 35296 41325
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 41259 35296 41260
rect 19616 40658 19936 40659
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 40593 19936 40594
rect 50336 40658 50656 40659
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 40593 50656 40594
rect 4256 39992 4576 39993
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 39927 4576 39928
rect 34976 39992 35296 39993
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 39927 35296 39928
rect 19616 39326 19936 39327
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 39261 19936 39262
rect 50336 39326 50656 39327
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 39261 50656 39262
rect 4256 38660 4576 38661
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 38595 4576 38596
rect 34976 38660 35296 38661
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 38595 35296 38596
rect 19616 37994 19936 37995
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 37929 19936 37930
rect 50336 37994 50656 37995
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 37929 50656 37930
rect 4256 37328 4576 37329
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 37263 4576 37264
rect 34976 37328 35296 37329
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 37263 35296 37264
rect 19616 36662 19936 36663
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 36597 19936 36598
rect 50336 36662 50656 36663
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 36597 50656 36598
rect 4256 35996 4576 35997
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 35931 4576 35932
rect 34976 35996 35296 35997
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 35931 35296 35932
rect 19616 35330 19936 35331
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 35265 19936 35266
rect 50336 35330 50656 35331
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 35265 50656 35266
rect 4256 34664 4576 34665
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 34599 4576 34600
rect 34976 34664 35296 34665
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 34599 35296 34600
rect 19616 33998 19936 33999
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 33933 19936 33934
rect 50336 33998 50656 33999
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 33933 50656 33934
rect 4256 33332 4576 33333
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 33267 4576 33268
rect 34976 33332 35296 33333
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 33267 35296 33268
rect 19616 32666 19936 32667
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 32601 19936 32602
rect 50336 32666 50656 32667
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 32601 50656 32602
rect 4256 32000 4576 32001
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 31935 4576 31936
rect 34976 32000 35296 32001
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 31935 35296 31936
rect 19616 31334 19936 31335
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 31269 19936 31270
rect 50336 31334 50656 31335
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 31269 50656 31270
rect 4256 30668 4576 30669
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 30603 4576 30604
rect 34976 30668 35296 30669
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 30603 35296 30604
rect 19616 30002 19936 30003
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 29937 19936 29938
rect 50336 30002 50656 30003
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 29937 50656 29938
rect 4256 29336 4576 29337
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 29271 4576 29272
rect 34976 29336 35296 29337
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 29271 35296 29272
rect 19616 28670 19936 28671
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 28605 19936 28606
rect 50336 28670 50656 28671
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 28605 50656 28606
rect 4256 28004 4576 28005
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 27939 4576 27940
rect 34976 28004 35296 28005
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 27939 35296 27940
rect 19616 27338 19936 27339
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 27273 19936 27274
rect 50336 27338 50656 27339
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 27273 50656 27274
rect 4256 26672 4576 26673
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 26607 4576 26608
rect 34976 26672 35296 26673
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 26607 35296 26608
rect 19616 26006 19936 26007
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 25941 19936 25942
rect 50336 26006 50656 26007
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 25941 50656 25942
rect 4256 25340 4576 25341
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 25275 4576 25276
rect 34976 25340 35296 25341
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 25275 35296 25276
rect 19616 24674 19936 24675
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 24609 19936 24610
rect 50336 24674 50656 24675
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 24609 50656 24610
rect 4256 24008 4576 24009
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 23943 4576 23944
rect 34976 24008 35296 24009
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 23943 35296 23944
rect 19616 23342 19936 23343
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 23277 19936 23278
rect 50336 23342 50656 23343
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 23277 50656 23278
rect 4256 22676 4576 22677
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 22611 4576 22612
rect 34976 22676 35296 22677
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 22611 35296 22612
rect 19616 22010 19936 22011
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 21945 19936 21946
rect 50336 22010 50656 22011
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 21945 50656 21946
rect 4256 21344 4576 21345
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 21279 4576 21280
rect 34976 21344 35296 21345
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 21279 35296 21280
rect 19616 20678 19936 20679
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 20613 19936 20614
rect 50336 20678 50656 20679
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 20613 50656 20614
rect 4256 20012 4576 20013
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 19947 4576 19948
rect 34976 20012 35296 20013
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 19947 35296 19948
rect 8271 19492 8337 19495
rect 9039 19492 9105 19495
rect 8271 19490 9105 19492
rect 8271 19434 8276 19490
rect 8332 19434 9044 19490
rect 9100 19434 9105 19490
rect 8271 19432 9105 19434
rect 8271 19429 8337 19432
rect 9039 19429 9105 19432
rect 19616 19346 19936 19347
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 19281 19936 19282
rect 50336 19346 50656 19347
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 19281 50656 19282
rect 4256 18680 4576 18681
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 18615 4576 18616
rect 34976 18680 35296 18681
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 18615 35296 18616
rect 19616 18014 19936 18015
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 17949 19936 17950
rect 50336 18014 50656 18015
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 17949 50656 17950
rect 4256 17348 4576 17349
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 17283 4576 17284
rect 34976 17348 35296 17349
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 17283 35296 17284
rect 19616 16682 19936 16683
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 16617 19936 16618
rect 50336 16682 50656 16683
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 16617 50656 16618
rect 4256 16016 4576 16017
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 15951 4576 15952
rect 34976 16016 35296 16017
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 15951 35296 15952
rect 19616 15350 19936 15351
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 15285 19936 15286
rect 50336 15350 50656 15351
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 15285 50656 15286
rect 4256 14684 4576 14685
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 14619 4576 14620
rect 34976 14684 35296 14685
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 14619 35296 14620
rect 19616 14018 19936 14019
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 13953 19936 13954
rect 50336 14018 50656 14019
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 13953 50656 13954
rect 4256 13352 4576 13353
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 13287 4576 13288
rect 34976 13352 35296 13353
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 13287 35296 13288
rect 19616 12686 19936 12687
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 12621 19936 12622
rect 50336 12686 50656 12687
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 12621 50656 12622
rect 4256 12020 4576 12021
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 11955 4576 11956
rect 34976 12020 35296 12021
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 11955 35296 11956
rect 19616 11354 19936 11355
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 11289 19936 11290
rect 50336 11354 50656 11355
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 11289 50656 11290
rect 4256 10688 4576 10689
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 10623 4576 10624
rect 34976 10688 35296 10689
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 10623 35296 10624
rect 19616 10022 19936 10023
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 9957 19936 9958
rect 50336 10022 50656 10023
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 9957 50656 9958
rect 4256 9356 4576 9357
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 9291 4576 9292
rect 34976 9356 35296 9357
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 9291 35296 9292
rect 19616 8690 19936 8691
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 8625 19936 8626
rect 50336 8690 50656 8691
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 8625 50656 8626
rect 4256 8024 4576 8025
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 7959 4576 7960
rect 34976 8024 35296 8025
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 7959 35296 7960
rect 7935 7800 8001 7803
rect 12975 7800 13041 7803
rect 7935 7798 13041 7800
rect 7935 7742 7940 7798
rect 7996 7742 12980 7798
rect 13036 7742 13041 7798
rect 7935 7740 13041 7742
rect 7935 7737 8001 7740
rect 12975 7737 13041 7740
rect 19616 7358 19936 7359
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 7293 19936 7294
rect 50336 7358 50656 7359
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 7293 50656 7294
rect 4256 6692 4576 6693
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 6627 4576 6628
rect 34976 6692 35296 6693
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 6627 35296 6628
rect 19616 6026 19936 6027
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 5961 19936 5962
rect 50336 6026 50656 6027
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 5961 50656 5962
rect 4256 5360 4576 5361
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 5295 4576 5296
rect 34976 5360 35296 5361
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 5295 35296 5296
rect 19616 4694 19936 4695
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 4629 19936 4630
rect 50336 4694 50656 4695
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 4629 50656 4630
rect 4256 4028 4576 4029
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 3963 4576 3964
rect 34976 4028 35296 4029
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 3963 35296 3964
rect 19616 3362 19936 3363
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 19616 3297 19936 3298
rect 50336 3362 50656 3363
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 50336 3297 50656 3298
rect 4256 2696 4576 2697
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4256 2631 4576 2632
rect 34976 2696 35296 2697
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 34976 2631 35296 2632
<< via3 >>
rect 4264 57304 4328 57308
rect 4264 57248 4268 57304
rect 4268 57248 4324 57304
rect 4324 57248 4328 57304
rect 4264 57244 4328 57248
rect 4344 57304 4408 57308
rect 4344 57248 4348 57304
rect 4348 57248 4404 57304
rect 4404 57248 4408 57304
rect 4344 57244 4408 57248
rect 4424 57304 4488 57308
rect 4424 57248 4428 57304
rect 4428 57248 4484 57304
rect 4484 57248 4488 57304
rect 4424 57244 4488 57248
rect 4504 57304 4568 57308
rect 4504 57248 4508 57304
rect 4508 57248 4564 57304
rect 4564 57248 4568 57304
rect 4504 57244 4568 57248
rect 34984 57304 35048 57308
rect 34984 57248 34988 57304
rect 34988 57248 35044 57304
rect 35044 57248 35048 57304
rect 34984 57244 35048 57248
rect 35064 57304 35128 57308
rect 35064 57248 35068 57304
rect 35068 57248 35124 57304
rect 35124 57248 35128 57304
rect 35064 57244 35128 57248
rect 35144 57304 35208 57308
rect 35144 57248 35148 57304
rect 35148 57248 35204 57304
rect 35204 57248 35208 57304
rect 35144 57244 35208 57248
rect 35224 57304 35288 57308
rect 35224 57248 35228 57304
rect 35228 57248 35284 57304
rect 35284 57248 35288 57304
rect 35224 57244 35288 57248
rect 19624 56638 19688 56642
rect 19624 56582 19628 56638
rect 19628 56582 19684 56638
rect 19684 56582 19688 56638
rect 19624 56578 19688 56582
rect 19704 56638 19768 56642
rect 19704 56582 19708 56638
rect 19708 56582 19764 56638
rect 19764 56582 19768 56638
rect 19704 56578 19768 56582
rect 19784 56638 19848 56642
rect 19784 56582 19788 56638
rect 19788 56582 19844 56638
rect 19844 56582 19848 56638
rect 19784 56578 19848 56582
rect 19864 56638 19928 56642
rect 19864 56582 19868 56638
rect 19868 56582 19924 56638
rect 19924 56582 19928 56638
rect 19864 56578 19928 56582
rect 50344 56638 50408 56642
rect 50344 56582 50348 56638
rect 50348 56582 50404 56638
rect 50404 56582 50408 56638
rect 50344 56578 50408 56582
rect 50424 56638 50488 56642
rect 50424 56582 50428 56638
rect 50428 56582 50484 56638
rect 50484 56582 50488 56638
rect 50424 56578 50488 56582
rect 50504 56638 50568 56642
rect 50504 56582 50508 56638
rect 50508 56582 50564 56638
rect 50564 56582 50568 56638
rect 50504 56578 50568 56582
rect 50584 56638 50648 56642
rect 50584 56582 50588 56638
rect 50588 56582 50644 56638
rect 50644 56582 50648 56638
rect 50584 56578 50648 56582
rect 4264 55972 4328 55976
rect 4264 55916 4268 55972
rect 4268 55916 4324 55972
rect 4324 55916 4328 55972
rect 4264 55912 4328 55916
rect 4344 55972 4408 55976
rect 4344 55916 4348 55972
rect 4348 55916 4404 55972
rect 4404 55916 4408 55972
rect 4344 55912 4408 55916
rect 4424 55972 4488 55976
rect 4424 55916 4428 55972
rect 4428 55916 4484 55972
rect 4484 55916 4488 55972
rect 4424 55912 4488 55916
rect 4504 55972 4568 55976
rect 4504 55916 4508 55972
rect 4508 55916 4564 55972
rect 4564 55916 4568 55972
rect 4504 55912 4568 55916
rect 34984 55972 35048 55976
rect 34984 55916 34988 55972
rect 34988 55916 35044 55972
rect 35044 55916 35048 55972
rect 34984 55912 35048 55916
rect 35064 55972 35128 55976
rect 35064 55916 35068 55972
rect 35068 55916 35124 55972
rect 35124 55916 35128 55972
rect 35064 55912 35128 55916
rect 35144 55972 35208 55976
rect 35144 55916 35148 55972
rect 35148 55916 35204 55972
rect 35204 55916 35208 55972
rect 35144 55912 35208 55916
rect 35224 55972 35288 55976
rect 35224 55916 35228 55972
rect 35228 55916 35284 55972
rect 35284 55916 35288 55972
rect 35224 55912 35288 55916
rect 19624 55306 19688 55310
rect 19624 55250 19628 55306
rect 19628 55250 19684 55306
rect 19684 55250 19688 55306
rect 19624 55246 19688 55250
rect 19704 55306 19768 55310
rect 19704 55250 19708 55306
rect 19708 55250 19764 55306
rect 19764 55250 19768 55306
rect 19704 55246 19768 55250
rect 19784 55306 19848 55310
rect 19784 55250 19788 55306
rect 19788 55250 19844 55306
rect 19844 55250 19848 55306
rect 19784 55246 19848 55250
rect 19864 55306 19928 55310
rect 19864 55250 19868 55306
rect 19868 55250 19924 55306
rect 19924 55250 19928 55306
rect 19864 55246 19928 55250
rect 50344 55306 50408 55310
rect 50344 55250 50348 55306
rect 50348 55250 50404 55306
rect 50404 55250 50408 55306
rect 50344 55246 50408 55250
rect 50424 55306 50488 55310
rect 50424 55250 50428 55306
rect 50428 55250 50484 55306
rect 50484 55250 50488 55306
rect 50424 55246 50488 55250
rect 50504 55306 50568 55310
rect 50504 55250 50508 55306
rect 50508 55250 50564 55306
rect 50564 55250 50568 55306
rect 50504 55246 50568 55250
rect 50584 55306 50648 55310
rect 50584 55250 50588 55306
rect 50588 55250 50644 55306
rect 50644 55250 50648 55306
rect 50584 55246 50648 55250
rect 4264 54640 4328 54644
rect 4264 54584 4268 54640
rect 4268 54584 4324 54640
rect 4324 54584 4328 54640
rect 4264 54580 4328 54584
rect 4344 54640 4408 54644
rect 4344 54584 4348 54640
rect 4348 54584 4404 54640
rect 4404 54584 4408 54640
rect 4344 54580 4408 54584
rect 4424 54640 4488 54644
rect 4424 54584 4428 54640
rect 4428 54584 4484 54640
rect 4484 54584 4488 54640
rect 4424 54580 4488 54584
rect 4504 54640 4568 54644
rect 4504 54584 4508 54640
rect 4508 54584 4564 54640
rect 4564 54584 4568 54640
rect 4504 54580 4568 54584
rect 34984 54640 35048 54644
rect 34984 54584 34988 54640
rect 34988 54584 35044 54640
rect 35044 54584 35048 54640
rect 34984 54580 35048 54584
rect 35064 54640 35128 54644
rect 35064 54584 35068 54640
rect 35068 54584 35124 54640
rect 35124 54584 35128 54640
rect 35064 54580 35128 54584
rect 35144 54640 35208 54644
rect 35144 54584 35148 54640
rect 35148 54584 35204 54640
rect 35204 54584 35208 54640
rect 35144 54580 35208 54584
rect 35224 54640 35288 54644
rect 35224 54584 35228 54640
rect 35228 54584 35284 54640
rect 35284 54584 35288 54640
rect 35224 54580 35288 54584
rect 19624 53974 19688 53978
rect 19624 53918 19628 53974
rect 19628 53918 19684 53974
rect 19684 53918 19688 53974
rect 19624 53914 19688 53918
rect 19704 53974 19768 53978
rect 19704 53918 19708 53974
rect 19708 53918 19764 53974
rect 19764 53918 19768 53974
rect 19704 53914 19768 53918
rect 19784 53974 19848 53978
rect 19784 53918 19788 53974
rect 19788 53918 19844 53974
rect 19844 53918 19848 53974
rect 19784 53914 19848 53918
rect 19864 53974 19928 53978
rect 19864 53918 19868 53974
rect 19868 53918 19924 53974
rect 19924 53918 19928 53974
rect 19864 53914 19928 53918
rect 50344 53974 50408 53978
rect 50344 53918 50348 53974
rect 50348 53918 50404 53974
rect 50404 53918 50408 53974
rect 50344 53914 50408 53918
rect 50424 53974 50488 53978
rect 50424 53918 50428 53974
rect 50428 53918 50484 53974
rect 50484 53918 50488 53974
rect 50424 53914 50488 53918
rect 50504 53974 50568 53978
rect 50504 53918 50508 53974
rect 50508 53918 50564 53974
rect 50564 53918 50568 53974
rect 50504 53914 50568 53918
rect 50584 53974 50648 53978
rect 50584 53918 50588 53974
rect 50588 53918 50644 53974
rect 50644 53918 50648 53974
rect 50584 53914 50648 53918
rect 4264 53308 4328 53312
rect 4264 53252 4268 53308
rect 4268 53252 4324 53308
rect 4324 53252 4328 53308
rect 4264 53248 4328 53252
rect 4344 53308 4408 53312
rect 4344 53252 4348 53308
rect 4348 53252 4404 53308
rect 4404 53252 4408 53308
rect 4344 53248 4408 53252
rect 4424 53308 4488 53312
rect 4424 53252 4428 53308
rect 4428 53252 4484 53308
rect 4484 53252 4488 53308
rect 4424 53248 4488 53252
rect 4504 53308 4568 53312
rect 4504 53252 4508 53308
rect 4508 53252 4564 53308
rect 4564 53252 4568 53308
rect 4504 53248 4568 53252
rect 34984 53308 35048 53312
rect 34984 53252 34988 53308
rect 34988 53252 35044 53308
rect 35044 53252 35048 53308
rect 34984 53248 35048 53252
rect 35064 53308 35128 53312
rect 35064 53252 35068 53308
rect 35068 53252 35124 53308
rect 35124 53252 35128 53308
rect 35064 53248 35128 53252
rect 35144 53308 35208 53312
rect 35144 53252 35148 53308
rect 35148 53252 35204 53308
rect 35204 53252 35208 53308
rect 35144 53248 35208 53252
rect 35224 53308 35288 53312
rect 35224 53252 35228 53308
rect 35228 53252 35284 53308
rect 35284 53252 35288 53308
rect 35224 53248 35288 53252
rect 19624 52642 19688 52646
rect 19624 52586 19628 52642
rect 19628 52586 19684 52642
rect 19684 52586 19688 52642
rect 19624 52582 19688 52586
rect 19704 52642 19768 52646
rect 19704 52586 19708 52642
rect 19708 52586 19764 52642
rect 19764 52586 19768 52642
rect 19704 52582 19768 52586
rect 19784 52642 19848 52646
rect 19784 52586 19788 52642
rect 19788 52586 19844 52642
rect 19844 52586 19848 52642
rect 19784 52582 19848 52586
rect 19864 52642 19928 52646
rect 19864 52586 19868 52642
rect 19868 52586 19924 52642
rect 19924 52586 19928 52642
rect 19864 52582 19928 52586
rect 50344 52642 50408 52646
rect 50344 52586 50348 52642
rect 50348 52586 50404 52642
rect 50404 52586 50408 52642
rect 50344 52582 50408 52586
rect 50424 52642 50488 52646
rect 50424 52586 50428 52642
rect 50428 52586 50484 52642
rect 50484 52586 50488 52642
rect 50424 52582 50488 52586
rect 50504 52642 50568 52646
rect 50504 52586 50508 52642
rect 50508 52586 50564 52642
rect 50564 52586 50568 52642
rect 50504 52582 50568 52586
rect 50584 52642 50648 52646
rect 50584 52586 50588 52642
rect 50588 52586 50644 52642
rect 50644 52586 50648 52642
rect 50584 52582 50648 52586
rect 4264 51976 4328 51980
rect 4264 51920 4268 51976
rect 4268 51920 4324 51976
rect 4324 51920 4328 51976
rect 4264 51916 4328 51920
rect 4344 51976 4408 51980
rect 4344 51920 4348 51976
rect 4348 51920 4404 51976
rect 4404 51920 4408 51976
rect 4344 51916 4408 51920
rect 4424 51976 4488 51980
rect 4424 51920 4428 51976
rect 4428 51920 4484 51976
rect 4484 51920 4488 51976
rect 4424 51916 4488 51920
rect 4504 51976 4568 51980
rect 4504 51920 4508 51976
rect 4508 51920 4564 51976
rect 4564 51920 4568 51976
rect 4504 51916 4568 51920
rect 34984 51976 35048 51980
rect 34984 51920 34988 51976
rect 34988 51920 35044 51976
rect 35044 51920 35048 51976
rect 34984 51916 35048 51920
rect 35064 51976 35128 51980
rect 35064 51920 35068 51976
rect 35068 51920 35124 51976
rect 35124 51920 35128 51976
rect 35064 51916 35128 51920
rect 35144 51976 35208 51980
rect 35144 51920 35148 51976
rect 35148 51920 35204 51976
rect 35204 51920 35208 51976
rect 35144 51916 35208 51920
rect 35224 51976 35288 51980
rect 35224 51920 35228 51976
rect 35228 51920 35284 51976
rect 35284 51920 35288 51976
rect 35224 51916 35288 51920
rect 19624 51310 19688 51314
rect 19624 51254 19628 51310
rect 19628 51254 19684 51310
rect 19684 51254 19688 51310
rect 19624 51250 19688 51254
rect 19704 51310 19768 51314
rect 19704 51254 19708 51310
rect 19708 51254 19764 51310
rect 19764 51254 19768 51310
rect 19704 51250 19768 51254
rect 19784 51310 19848 51314
rect 19784 51254 19788 51310
rect 19788 51254 19844 51310
rect 19844 51254 19848 51310
rect 19784 51250 19848 51254
rect 19864 51310 19928 51314
rect 19864 51254 19868 51310
rect 19868 51254 19924 51310
rect 19924 51254 19928 51310
rect 19864 51250 19928 51254
rect 50344 51310 50408 51314
rect 50344 51254 50348 51310
rect 50348 51254 50404 51310
rect 50404 51254 50408 51310
rect 50344 51250 50408 51254
rect 50424 51310 50488 51314
rect 50424 51254 50428 51310
rect 50428 51254 50484 51310
rect 50484 51254 50488 51310
rect 50424 51250 50488 51254
rect 50504 51310 50568 51314
rect 50504 51254 50508 51310
rect 50508 51254 50564 51310
rect 50564 51254 50568 51310
rect 50504 51250 50568 51254
rect 50584 51310 50648 51314
rect 50584 51254 50588 51310
rect 50588 51254 50644 51310
rect 50644 51254 50648 51310
rect 50584 51250 50648 51254
rect 4264 50644 4328 50648
rect 4264 50588 4268 50644
rect 4268 50588 4324 50644
rect 4324 50588 4328 50644
rect 4264 50584 4328 50588
rect 4344 50644 4408 50648
rect 4344 50588 4348 50644
rect 4348 50588 4404 50644
rect 4404 50588 4408 50644
rect 4344 50584 4408 50588
rect 4424 50644 4488 50648
rect 4424 50588 4428 50644
rect 4428 50588 4484 50644
rect 4484 50588 4488 50644
rect 4424 50584 4488 50588
rect 4504 50644 4568 50648
rect 4504 50588 4508 50644
rect 4508 50588 4564 50644
rect 4564 50588 4568 50644
rect 4504 50584 4568 50588
rect 34984 50644 35048 50648
rect 34984 50588 34988 50644
rect 34988 50588 35044 50644
rect 35044 50588 35048 50644
rect 34984 50584 35048 50588
rect 35064 50644 35128 50648
rect 35064 50588 35068 50644
rect 35068 50588 35124 50644
rect 35124 50588 35128 50644
rect 35064 50584 35128 50588
rect 35144 50644 35208 50648
rect 35144 50588 35148 50644
rect 35148 50588 35204 50644
rect 35204 50588 35208 50644
rect 35144 50584 35208 50588
rect 35224 50644 35288 50648
rect 35224 50588 35228 50644
rect 35228 50588 35284 50644
rect 35284 50588 35288 50644
rect 35224 50584 35288 50588
rect 19624 49978 19688 49982
rect 19624 49922 19628 49978
rect 19628 49922 19684 49978
rect 19684 49922 19688 49978
rect 19624 49918 19688 49922
rect 19704 49978 19768 49982
rect 19704 49922 19708 49978
rect 19708 49922 19764 49978
rect 19764 49922 19768 49978
rect 19704 49918 19768 49922
rect 19784 49978 19848 49982
rect 19784 49922 19788 49978
rect 19788 49922 19844 49978
rect 19844 49922 19848 49978
rect 19784 49918 19848 49922
rect 19864 49978 19928 49982
rect 19864 49922 19868 49978
rect 19868 49922 19924 49978
rect 19924 49922 19928 49978
rect 19864 49918 19928 49922
rect 50344 49978 50408 49982
rect 50344 49922 50348 49978
rect 50348 49922 50404 49978
rect 50404 49922 50408 49978
rect 50344 49918 50408 49922
rect 50424 49978 50488 49982
rect 50424 49922 50428 49978
rect 50428 49922 50484 49978
rect 50484 49922 50488 49978
rect 50424 49918 50488 49922
rect 50504 49978 50568 49982
rect 50504 49922 50508 49978
rect 50508 49922 50564 49978
rect 50564 49922 50568 49978
rect 50504 49918 50568 49922
rect 50584 49978 50648 49982
rect 50584 49922 50588 49978
rect 50588 49922 50644 49978
rect 50644 49922 50648 49978
rect 50584 49918 50648 49922
rect 4264 49312 4328 49316
rect 4264 49256 4268 49312
rect 4268 49256 4324 49312
rect 4324 49256 4328 49312
rect 4264 49252 4328 49256
rect 4344 49312 4408 49316
rect 4344 49256 4348 49312
rect 4348 49256 4404 49312
rect 4404 49256 4408 49312
rect 4344 49252 4408 49256
rect 4424 49312 4488 49316
rect 4424 49256 4428 49312
rect 4428 49256 4484 49312
rect 4484 49256 4488 49312
rect 4424 49252 4488 49256
rect 4504 49312 4568 49316
rect 4504 49256 4508 49312
rect 4508 49256 4564 49312
rect 4564 49256 4568 49312
rect 4504 49252 4568 49256
rect 34984 49312 35048 49316
rect 34984 49256 34988 49312
rect 34988 49256 35044 49312
rect 35044 49256 35048 49312
rect 34984 49252 35048 49256
rect 35064 49312 35128 49316
rect 35064 49256 35068 49312
rect 35068 49256 35124 49312
rect 35124 49256 35128 49312
rect 35064 49252 35128 49256
rect 35144 49312 35208 49316
rect 35144 49256 35148 49312
rect 35148 49256 35204 49312
rect 35204 49256 35208 49312
rect 35144 49252 35208 49256
rect 35224 49312 35288 49316
rect 35224 49256 35228 49312
rect 35228 49256 35284 49312
rect 35284 49256 35288 49312
rect 35224 49252 35288 49256
rect 19624 48646 19688 48650
rect 19624 48590 19628 48646
rect 19628 48590 19684 48646
rect 19684 48590 19688 48646
rect 19624 48586 19688 48590
rect 19704 48646 19768 48650
rect 19704 48590 19708 48646
rect 19708 48590 19764 48646
rect 19764 48590 19768 48646
rect 19704 48586 19768 48590
rect 19784 48646 19848 48650
rect 19784 48590 19788 48646
rect 19788 48590 19844 48646
rect 19844 48590 19848 48646
rect 19784 48586 19848 48590
rect 19864 48646 19928 48650
rect 19864 48590 19868 48646
rect 19868 48590 19924 48646
rect 19924 48590 19928 48646
rect 19864 48586 19928 48590
rect 50344 48646 50408 48650
rect 50344 48590 50348 48646
rect 50348 48590 50404 48646
rect 50404 48590 50408 48646
rect 50344 48586 50408 48590
rect 50424 48646 50488 48650
rect 50424 48590 50428 48646
rect 50428 48590 50484 48646
rect 50484 48590 50488 48646
rect 50424 48586 50488 48590
rect 50504 48646 50568 48650
rect 50504 48590 50508 48646
rect 50508 48590 50564 48646
rect 50564 48590 50568 48646
rect 50504 48586 50568 48590
rect 50584 48646 50648 48650
rect 50584 48590 50588 48646
rect 50588 48590 50644 48646
rect 50644 48590 50648 48646
rect 50584 48586 50648 48590
rect 4264 47980 4328 47984
rect 4264 47924 4268 47980
rect 4268 47924 4324 47980
rect 4324 47924 4328 47980
rect 4264 47920 4328 47924
rect 4344 47980 4408 47984
rect 4344 47924 4348 47980
rect 4348 47924 4404 47980
rect 4404 47924 4408 47980
rect 4344 47920 4408 47924
rect 4424 47980 4488 47984
rect 4424 47924 4428 47980
rect 4428 47924 4484 47980
rect 4484 47924 4488 47980
rect 4424 47920 4488 47924
rect 4504 47980 4568 47984
rect 4504 47924 4508 47980
rect 4508 47924 4564 47980
rect 4564 47924 4568 47980
rect 4504 47920 4568 47924
rect 34984 47980 35048 47984
rect 34984 47924 34988 47980
rect 34988 47924 35044 47980
rect 35044 47924 35048 47980
rect 34984 47920 35048 47924
rect 35064 47980 35128 47984
rect 35064 47924 35068 47980
rect 35068 47924 35124 47980
rect 35124 47924 35128 47980
rect 35064 47920 35128 47924
rect 35144 47980 35208 47984
rect 35144 47924 35148 47980
rect 35148 47924 35204 47980
rect 35204 47924 35208 47980
rect 35144 47920 35208 47924
rect 35224 47980 35288 47984
rect 35224 47924 35228 47980
rect 35228 47924 35284 47980
rect 35284 47924 35288 47980
rect 35224 47920 35288 47924
rect 19624 47314 19688 47318
rect 19624 47258 19628 47314
rect 19628 47258 19684 47314
rect 19684 47258 19688 47314
rect 19624 47254 19688 47258
rect 19704 47314 19768 47318
rect 19704 47258 19708 47314
rect 19708 47258 19764 47314
rect 19764 47258 19768 47314
rect 19704 47254 19768 47258
rect 19784 47314 19848 47318
rect 19784 47258 19788 47314
rect 19788 47258 19844 47314
rect 19844 47258 19848 47314
rect 19784 47254 19848 47258
rect 19864 47314 19928 47318
rect 19864 47258 19868 47314
rect 19868 47258 19924 47314
rect 19924 47258 19928 47314
rect 19864 47254 19928 47258
rect 50344 47314 50408 47318
rect 50344 47258 50348 47314
rect 50348 47258 50404 47314
rect 50404 47258 50408 47314
rect 50344 47254 50408 47258
rect 50424 47314 50488 47318
rect 50424 47258 50428 47314
rect 50428 47258 50484 47314
rect 50484 47258 50488 47314
rect 50424 47254 50488 47258
rect 50504 47314 50568 47318
rect 50504 47258 50508 47314
rect 50508 47258 50564 47314
rect 50564 47258 50568 47314
rect 50504 47254 50568 47258
rect 50584 47314 50648 47318
rect 50584 47258 50588 47314
rect 50588 47258 50644 47314
rect 50644 47258 50648 47314
rect 50584 47254 50648 47258
rect 4264 46648 4328 46652
rect 4264 46592 4268 46648
rect 4268 46592 4324 46648
rect 4324 46592 4328 46648
rect 4264 46588 4328 46592
rect 4344 46648 4408 46652
rect 4344 46592 4348 46648
rect 4348 46592 4404 46648
rect 4404 46592 4408 46648
rect 4344 46588 4408 46592
rect 4424 46648 4488 46652
rect 4424 46592 4428 46648
rect 4428 46592 4484 46648
rect 4484 46592 4488 46648
rect 4424 46588 4488 46592
rect 4504 46648 4568 46652
rect 4504 46592 4508 46648
rect 4508 46592 4564 46648
rect 4564 46592 4568 46648
rect 4504 46588 4568 46592
rect 34984 46648 35048 46652
rect 34984 46592 34988 46648
rect 34988 46592 35044 46648
rect 35044 46592 35048 46648
rect 34984 46588 35048 46592
rect 35064 46648 35128 46652
rect 35064 46592 35068 46648
rect 35068 46592 35124 46648
rect 35124 46592 35128 46648
rect 35064 46588 35128 46592
rect 35144 46648 35208 46652
rect 35144 46592 35148 46648
rect 35148 46592 35204 46648
rect 35204 46592 35208 46648
rect 35144 46588 35208 46592
rect 35224 46648 35288 46652
rect 35224 46592 35228 46648
rect 35228 46592 35284 46648
rect 35284 46592 35288 46648
rect 35224 46588 35288 46592
rect 19624 45982 19688 45986
rect 19624 45926 19628 45982
rect 19628 45926 19684 45982
rect 19684 45926 19688 45982
rect 19624 45922 19688 45926
rect 19704 45982 19768 45986
rect 19704 45926 19708 45982
rect 19708 45926 19764 45982
rect 19764 45926 19768 45982
rect 19704 45922 19768 45926
rect 19784 45982 19848 45986
rect 19784 45926 19788 45982
rect 19788 45926 19844 45982
rect 19844 45926 19848 45982
rect 19784 45922 19848 45926
rect 19864 45982 19928 45986
rect 19864 45926 19868 45982
rect 19868 45926 19924 45982
rect 19924 45926 19928 45982
rect 19864 45922 19928 45926
rect 50344 45982 50408 45986
rect 50344 45926 50348 45982
rect 50348 45926 50404 45982
rect 50404 45926 50408 45982
rect 50344 45922 50408 45926
rect 50424 45982 50488 45986
rect 50424 45926 50428 45982
rect 50428 45926 50484 45982
rect 50484 45926 50488 45982
rect 50424 45922 50488 45926
rect 50504 45982 50568 45986
rect 50504 45926 50508 45982
rect 50508 45926 50564 45982
rect 50564 45926 50568 45982
rect 50504 45922 50568 45926
rect 50584 45982 50648 45986
rect 50584 45926 50588 45982
rect 50588 45926 50644 45982
rect 50644 45926 50648 45982
rect 50584 45922 50648 45926
rect 4264 45316 4328 45320
rect 4264 45260 4268 45316
rect 4268 45260 4324 45316
rect 4324 45260 4328 45316
rect 4264 45256 4328 45260
rect 4344 45316 4408 45320
rect 4344 45260 4348 45316
rect 4348 45260 4404 45316
rect 4404 45260 4408 45316
rect 4344 45256 4408 45260
rect 4424 45316 4488 45320
rect 4424 45260 4428 45316
rect 4428 45260 4484 45316
rect 4484 45260 4488 45316
rect 4424 45256 4488 45260
rect 4504 45316 4568 45320
rect 4504 45260 4508 45316
rect 4508 45260 4564 45316
rect 4564 45260 4568 45316
rect 4504 45256 4568 45260
rect 34984 45316 35048 45320
rect 34984 45260 34988 45316
rect 34988 45260 35044 45316
rect 35044 45260 35048 45316
rect 34984 45256 35048 45260
rect 35064 45316 35128 45320
rect 35064 45260 35068 45316
rect 35068 45260 35124 45316
rect 35124 45260 35128 45316
rect 35064 45256 35128 45260
rect 35144 45316 35208 45320
rect 35144 45260 35148 45316
rect 35148 45260 35204 45316
rect 35204 45260 35208 45316
rect 35144 45256 35208 45260
rect 35224 45316 35288 45320
rect 35224 45260 35228 45316
rect 35228 45260 35284 45316
rect 35284 45260 35288 45316
rect 35224 45256 35288 45260
rect 19624 44650 19688 44654
rect 19624 44594 19628 44650
rect 19628 44594 19684 44650
rect 19684 44594 19688 44650
rect 19624 44590 19688 44594
rect 19704 44650 19768 44654
rect 19704 44594 19708 44650
rect 19708 44594 19764 44650
rect 19764 44594 19768 44650
rect 19704 44590 19768 44594
rect 19784 44650 19848 44654
rect 19784 44594 19788 44650
rect 19788 44594 19844 44650
rect 19844 44594 19848 44650
rect 19784 44590 19848 44594
rect 19864 44650 19928 44654
rect 19864 44594 19868 44650
rect 19868 44594 19924 44650
rect 19924 44594 19928 44650
rect 19864 44590 19928 44594
rect 50344 44650 50408 44654
rect 50344 44594 50348 44650
rect 50348 44594 50404 44650
rect 50404 44594 50408 44650
rect 50344 44590 50408 44594
rect 50424 44650 50488 44654
rect 50424 44594 50428 44650
rect 50428 44594 50484 44650
rect 50484 44594 50488 44650
rect 50424 44590 50488 44594
rect 50504 44650 50568 44654
rect 50504 44594 50508 44650
rect 50508 44594 50564 44650
rect 50564 44594 50568 44650
rect 50504 44590 50568 44594
rect 50584 44650 50648 44654
rect 50584 44594 50588 44650
rect 50588 44594 50644 44650
rect 50644 44594 50648 44650
rect 50584 44590 50648 44594
rect 4264 43984 4328 43988
rect 4264 43928 4268 43984
rect 4268 43928 4324 43984
rect 4324 43928 4328 43984
rect 4264 43924 4328 43928
rect 4344 43984 4408 43988
rect 4344 43928 4348 43984
rect 4348 43928 4404 43984
rect 4404 43928 4408 43984
rect 4344 43924 4408 43928
rect 4424 43984 4488 43988
rect 4424 43928 4428 43984
rect 4428 43928 4484 43984
rect 4484 43928 4488 43984
rect 4424 43924 4488 43928
rect 4504 43984 4568 43988
rect 4504 43928 4508 43984
rect 4508 43928 4564 43984
rect 4564 43928 4568 43984
rect 4504 43924 4568 43928
rect 34984 43984 35048 43988
rect 34984 43928 34988 43984
rect 34988 43928 35044 43984
rect 35044 43928 35048 43984
rect 34984 43924 35048 43928
rect 35064 43984 35128 43988
rect 35064 43928 35068 43984
rect 35068 43928 35124 43984
rect 35124 43928 35128 43984
rect 35064 43924 35128 43928
rect 35144 43984 35208 43988
rect 35144 43928 35148 43984
rect 35148 43928 35204 43984
rect 35204 43928 35208 43984
rect 35144 43924 35208 43928
rect 35224 43984 35288 43988
rect 35224 43928 35228 43984
rect 35228 43928 35284 43984
rect 35284 43928 35288 43984
rect 35224 43924 35288 43928
rect 19624 43318 19688 43322
rect 19624 43262 19628 43318
rect 19628 43262 19684 43318
rect 19684 43262 19688 43318
rect 19624 43258 19688 43262
rect 19704 43318 19768 43322
rect 19704 43262 19708 43318
rect 19708 43262 19764 43318
rect 19764 43262 19768 43318
rect 19704 43258 19768 43262
rect 19784 43318 19848 43322
rect 19784 43262 19788 43318
rect 19788 43262 19844 43318
rect 19844 43262 19848 43318
rect 19784 43258 19848 43262
rect 19864 43318 19928 43322
rect 19864 43262 19868 43318
rect 19868 43262 19924 43318
rect 19924 43262 19928 43318
rect 19864 43258 19928 43262
rect 50344 43318 50408 43322
rect 50344 43262 50348 43318
rect 50348 43262 50404 43318
rect 50404 43262 50408 43318
rect 50344 43258 50408 43262
rect 50424 43318 50488 43322
rect 50424 43262 50428 43318
rect 50428 43262 50484 43318
rect 50484 43262 50488 43318
rect 50424 43258 50488 43262
rect 50504 43318 50568 43322
rect 50504 43262 50508 43318
rect 50508 43262 50564 43318
rect 50564 43262 50568 43318
rect 50504 43258 50568 43262
rect 50584 43318 50648 43322
rect 50584 43262 50588 43318
rect 50588 43262 50644 43318
rect 50644 43262 50648 43318
rect 50584 43258 50648 43262
rect 4264 42652 4328 42656
rect 4264 42596 4268 42652
rect 4268 42596 4324 42652
rect 4324 42596 4328 42652
rect 4264 42592 4328 42596
rect 4344 42652 4408 42656
rect 4344 42596 4348 42652
rect 4348 42596 4404 42652
rect 4404 42596 4408 42652
rect 4344 42592 4408 42596
rect 4424 42652 4488 42656
rect 4424 42596 4428 42652
rect 4428 42596 4484 42652
rect 4484 42596 4488 42652
rect 4424 42592 4488 42596
rect 4504 42652 4568 42656
rect 4504 42596 4508 42652
rect 4508 42596 4564 42652
rect 4564 42596 4568 42652
rect 4504 42592 4568 42596
rect 34984 42652 35048 42656
rect 34984 42596 34988 42652
rect 34988 42596 35044 42652
rect 35044 42596 35048 42652
rect 34984 42592 35048 42596
rect 35064 42652 35128 42656
rect 35064 42596 35068 42652
rect 35068 42596 35124 42652
rect 35124 42596 35128 42652
rect 35064 42592 35128 42596
rect 35144 42652 35208 42656
rect 35144 42596 35148 42652
rect 35148 42596 35204 42652
rect 35204 42596 35208 42652
rect 35144 42592 35208 42596
rect 35224 42652 35288 42656
rect 35224 42596 35228 42652
rect 35228 42596 35284 42652
rect 35284 42596 35288 42652
rect 35224 42592 35288 42596
rect 19624 41986 19688 41990
rect 19624 41930 19628 41986
rect 19628 41930 19684 41986
rect 19684 41930 19688 41986
rect 19624 41926 19688 41930
rect 19704 41986 19768 41990
rect 19704 41930 19708 41986
rect 19708 41930 19764 41986
rect 19764 41930 19768 41986
rect 19704 41926 19768 41930
rect 19784 41986 19848 41990
rect 19784 41930 19788 41986
rect 19788 41930 19844 41986
rect 19844 41930 19848 41986
rect 19784 41926 19848 41930
rect 19864 41986 19928 41990
rect 19864 41930 19868 41986
rect 19868 41930 19924 41986
rect 19924 41930 19928 41986
rect 19864 41926 19928 41930
rect 50344 41986 50408 41990
rect 50344 41930 50348 41986
rect 50348 41930 50404 41986
rect 50404 41930 50408 41986
rect 50344 41926 50408 41930
rect 50424 41986 50488 41990
rect 50424 41930 50428 41986
rect 50428 41930 50484 41986
rect 50484 41930 50488 41986
rect 50424 41926 50488 41930
rect 50504 41986 50568 41990
rect 50504 41930 50508 41986
rect 50508 41930 50564 41986
rect 50564 41930 50568 41986
rect 50504 41926 50568 41930
rect 50584 41986 50648 41990
rect 50584 41930 50588 41986
rect 50588 41930 50644 41986
rect 50644 41930 50648 41986
rect 50584 41926 50648 41930
rect 4264 41320 4328 41324
rect 4264 41264 4268 41320
rect 4268 41264 4324 41320
rect 4324 41264 4328 41320
rect 4264 41260 4328 41264
rect 4344 41320 4408 41324
rect 4344 41264 4348 41320
rect 4348 41264 4404 41320
rect 4404 41264 4408 41320
rect 4344 41260 4408 41264
rect 4424 41320 4488 41324
rect 4424 41264 4428 41320
rect 4428 41264 4484 41320
rect 4484 41264 4488 41320
rect 4424 41260 4488 41264
rect 4504 41320 4568 41324
rect 4504 41264 4508 41320
rect 4508 41264 4564 41320
rect 4564 41264 4568 41320
rect 4504 41260 4568 41264
rect 34984 41320 35048 41324
rect 34984 41264 34988 41320
rect 34988 41264 35044 41320
rect 35044 41264 35048 41320
rect 34984 41260 35048 41264
rect 35064 41320 35128 41324
rect 35064 41264 35068 41320
rect 35068 41264 35124 41320
rect 35124 41264 35128 41320
rect 35064 41260 35128 41264
rect 35144 41320 35208 41324
rect 35144 41264 35148 41320
rect 35148 41264 35204 41320
rect 35204 41264 35208 41320
rect 35144 41260 35208 41264
rect 35224 41320 35288 41324
rect 35224 41264 35228 41320
rect 35228 41264 35284 41320
rect 35284 41264 35288 41320
rect 35224 41260 35288 41264
rect 19624 40654 19688 40658
rect 19624 40598 19628 40654
rect 19628 40598 19684 40654
rect 19684 40598 19688 40654
rect 19624 40594 19688 40598
rect 19704 40654 19768 40658
rect 19704 40598 19708 40654
rect 19708 40598 19764 40654
rect 19764 40598 19768 40654
rect 19704 40594 19768 40598
rect 19784 40654 19848 40658
rect 19784 40598 19788 40654
rect 19788 40598 19844 40654
rect 19844 40598 19848 40654
rect 19784 40594 19848 40598
rect 19864 40654 19928 40658
rect 19864 40598 19868 40654
rect 19868 40598 19924 40654
rect 19924 40598 19928 40654
rect 19864 40594 19928 40598
rect 50344 40654 50408 40658
rect 50344 40598 50348 40654
rect 50348 40598 50404 40654
rect 50404 40598 50408 40654
rect 50344 40594 50408 40598
rect 50424 40654 50488 40658
rect 50424 40598 50428 40654
rect 50428 40598 50484 40654
rect 50484 40598 50488 40654
rect 50424 40594 50488 40598
rect 50504 40654 50568 40658
rect 50504 40598 50508 40654
rect 50508 40598 50564 40654
rect 50564 40598 50568 40654
rect 50504 40594 50568 40598
rect 50584 40654 50648 40658
rect 50584 40598 50588 40654
rect 50588 40598 50644 40654
rect 50644 40598 50648 40654
rect 50584 40594 50648 40598
rect 4264 39988 4328 39992
rect 4264 39932 4268 39988
rect 4268 39932 4324 39988
rect 4324 39932 4328 39988
rect 4264 39928 4328 39932
rect 4344 39988 4408 39992
rect 4344 39932 4348 39988
rect 4348 39932 4404 39988
rect 4404 39932 4408 39988
rect 4344 39928 4408 39932
rect 4424 39988 4488 39992
rect 4424 39932 4428 39988
rect 4428 39932 4484 39988
rect 4484 39932 4488 39988
rect 4424 39928 4488 39932
rect 4504 39988 4568 39992
rect 4504 39932 4508 39988
rect 4508 39932 4564 39988
rect 4564 39932 4568 39988
rect 4504 39928 4568 39932
rect 34984 39988 35048 39992
rect 34984 39932 34988 39988
rect 34988 39932 35044 39988
rect 35044 39932 35048 39988
rect 34984 39928 35048 39932
rect 35064 39988 35128 39992
rect 35064 39932 35068 39988
rect 35068 39932 35124 39988
rect 35124 39932 35128 39988
rect 35064 39928 35128 39932
rect 35144 39988 35208 39992
rect 35144 39932 35148 39988
rect 35148 39932 35204 39988
rect 35204 39932 35208 39988
rect 35144 39928 35208 39932
rect 35224 39988 35288 39992
rect 35224 39932 35228 39988
rect 35228 39932 35284 39988
rect 35284 39932 35288 39988
rect 35224 39928 35288 39932
rect 19624 39322 19688 39326
rect 19624 39266 19628 39322
rect 19628 39266 19684 39322
rect 19684 39266 19688 39322
rect 19624 39262 19688 39266
rect 19704 39322 19768 39326
rect 19704 39266 19708 39322
rect 19708 39266 19764 39322
rect 19764 39266 19768 39322
rect 19704 39262 19768 39266
rect 19784 39322 19848 39326
rect 19784 39266 19788 39322
rect 19788 39266 19844 39322
rect 19844 39266 19848 39322
rect 19784 39262 19848 39266
rect 19864 39322 19928 39326
rect 19864 39266 19868 39322
rect 19868 39266 19924 39322
rect 19924 39266 19928 39322
rect 19864 39262 19928 39266
rect 50344 39322 50408 39326
rect 50344 39266 50348 39322
rect 50348 39266 50404 39322
rect 50404 39266 50408 39322
rect 50344 39262 50408 39266
rect 50424 39322 50488 39326
rect 50424 39266 50428 39322
rect 50428 39266 50484 39322
rect 50484 39266 50488 39322
rect 50424 39262 50488 39266
rect 50504 39322 50568 39326
rect 50504 39266 50508 39322
rect 50508 39266 50564 39322
rect 50564 39266 50568 39322
rect 50504 39262 50568 39266
rect 50584 39322 50648 39326
rect 50584 39266 50588 39322
rect 50588 39266 50644 39322
rect 50644 39266 50648 39322
rect 50584 39262 50648 39266
rect 4264 38656 4328 38660
rect 4264 38600 4268 38656
rect 4268 38600 4324 38656
rect 4324 38600 4328 38656
rect 4264 38596 4328 38600
rect 4344 38656 4408 38660
rect 4344 38600 4348 38656
rect 4348 38600 4404 38656
rect 4404 38600 4408 38656
rect 4344 38596 4408 38600
rect 4424 38656 4488 38660
rect 4424 38600 4428 38656
rect 4428 38600 4484 38656
rect 4484 38600 4488 38656
rect 4424 38596 4488 38600
rect 4504 38656 4568 38660
rect 4504 38600 4508 38656
rect 4508 38600 4564 38656
rect 4564 38600 4568 38656
rect 4504 38596 4568 38600
rect 34984 38656 35048 38660
rect 34984 38600 34988 38656
rect 34988 38600 35044 38656
rect 35044 38600 35048 38656
rect 34984 38596 35048 38600
rect 35064 38656 35128 38660
rect 35064 38600 35068 38656
rect 35068 38600 35124 38656
rect 35124 38600 35128 38656
rect 35064 38596 35128 38600
rect 35144 38656 35208 38660
rect 35144 38600 35148 38656
rect 35148 38600 35204 38656
rect 35204 38600 35208 38656
rect 35144 38596 35208 38600
rect 35224 38656 35288 38660
rect 35224 38600 35228 38656
rect 35228 38600 35284 38656
rect 35284 38600 35288 38656
rect 35224 38596 35288 38600
rect 19624 37990 19688 37994
rect 19624 37934 19628 37990
rect 19628 37934 19684 37990
rect 19684 37934 19688 37990
rect 19624 37930 19688 37934
rect 19704 37990 19768 37994
rect 19704 37934 19708 37990
rect 19708 37934 19764 37990
rect 19764 37934 19768 37990
rect 19704 37930 19768 37934
rect 19784 37990 19848 37994
rect 19784 37934 19788 37990
rect 19788 37934 19844 37990
rect 19844 37934 19848 37990
rect 19784 37930 19848 37934
rect 19864 37990 19928 37994
rect 19864 37934 19868 37990
rect 19868 37934 19924 37990
rect 19924 37934 19928 37990
rect 19864 37930 19928 37934
rect 50344 37990 50408 37994
rect 50344 37934 50348 37990
rect 50348 37934 50404 37990
rect 50404 37934 50408 37990
rect 50344 37930 50408 37934
rect 50424 37990 50488 37994
rect 50424 37934 50428 37990
rect 50428 37934 50484 37990
rect 50484 37934 50488 37990
rect 50424 37930 50488 37934
rect 50504 37990 50568 37994
rect 50504 37934 50508 37990
rect 50508 37934 50564 37990
rect 50564 37934 50568 37990
rect 50504 37930 50568 37934
rect 50584 37990 50648 37994
rect 50584 37934 50588 37990
rect 50588 37934 50644 37990
rect 50644 37934 50648 37990
rect 50584 37930 50648 37934
rect 4264 37324 4328 37328
rect 4264 37268 4268 37324
rect 4268 37268 4324 37324
rect 4324 37268 4328 37324
rect 4264 37264 4328 37268
rect 4344 37324 4408 37328
rect 4344 37268 4348 37324
rect 4348 37268 4404 37324
rect 4404 37268 4408 37324
rect 4344 37264 4408 37268
rect 4424 37324 4488 37328
rect 4424 37268 4428 37324
rect 4428 37268 4484 37324
rect 4484 37268 4488 37324
rect 4424 37264 4488 37268
rect 4504 37324 4568 37328
rect 4504 37268 4508 37324
rect 4508 37268 4564 37324
rect 4564 37268 4568 37324
rect 4504 37264 4568 37268
rect 34984 37324 35048 37328
rect 34984 37268 34988 37324
rect 34988 37268 35044 37324
rect 35044 37268 35048 37324
rect 34984 37264 35048 37268
rect 35064 37324 35128 37328
rect 35064 37268 35068 37324
rect 35068 37268 35124 37324
rect 35124 37268 35128 37324
rect 35064 37264 35128 37268
rect 35144 37324 35208 37328
rect 35144 37268 35148 37324
rect 35148 37268 35204 37324
rect 35204 37268 35208 37324
rect 35144 37264 35208 37268
rect 35224 37324 35288 37328
rect 35224 37268 35228 37324
rect 35228 37268 35284 37324
rect 35284 37268 35288 37324
rect 35224 37264 35288 37268
rect 19624 36658 19688 36662
rect 19624 36602 19628 36658
rect 19628 36602 19684 36658
rect 19684 36602 19688 36658
rect 19624 36598 19688 36602
rect 19704 36658 19768 36662
rect 19704 36602 19708 36658
rect 19708 36602 19764 36658
rect 19764 36602 19768 36658
rect 19704 36598 19768 36602
rect 19784 36658 19848 36662
rect 19784 36602 19788 36658
rect 19788 36602 19844 36658
rect 19844 36602 19848 36658
rect 19784 36598 19848 36602
rect 19864 36658 19928 36662
rect 19864 36602 19868 36658
rect 19868 36602 19924 36658
rect 19924 36602 19928 36658
rect 19864 36598 19928 36602
rect 50344 36658 50408 36662
rect 50344 36602 50348 36658
rect 50348 36602 50404 36658
rect 50404 36602 50408 36658
rect 50344 36598 50408 36602
rect 50424 36658 50488 36662
rect 50424 36602 50428 36658
rect 50428 36602 50484 36658
rect 50484 36602 50488 36658
rect 50424 36598 50488 36602
rect 50504 36658 50568 36662
rect 50504 36602 50508 36658
rect 50508 36602 50564 36658
rect 50564 36602 50568 36658
rect 50504 36598 50568 36602
rect 50584 36658 50648 36662
rect 50584 36602 50588 36658
rect 50588 36602 50644 36658
rect 50644 36602 50648 36658
rect 50584 36598 50648 36602
rect 4264 35992 4328 35996
rect 4264 35936 4268 35992
rect 4268 35936 4324 35992
rect 4324 35936 4328 35992
rect 4264 35932 4328 35936
rect 4344 35992 4408 35996
rect 4344 35936 4348 35992
rect 4348 35936 4404 35992
rect 4404 35936 4408 35992
rect 4344 35932 4408 35936
rect 4424 35992 4488 35996
rect 4424 35936 4428 35992
rect 4428 35936 4484 35992
rect 4484 35936 4488 35992
rect 4424 35932 4488 35936
rect 4504 35992 4568 35996
rect 4504 35936 4508 35992
rect 4508 35936 4564 35992
rect 4564 35936 4568 35992
rect 4504 35932 4568 35936
rect 34984 35992 35048 35996
rect 34984 35936 34988 35992
rect 34988 35936 35044 35992
rect 35044 35936 35048 35992
rect 34984 35932 35048 35936
rect 35064 35992 35128 35996
rect 35064 35936 35068 35992
rect 35068 35936 35124 35992
rect 35124 35936 35128 35992
rect 35064 35932 35128 35936
rect 35144 35992 35208 35996
rect 35144 35936 35148 35992
rect 35148 35936 35204 35992
rect 35204 35936 35208 35992
rect 35144 35932 35208 35936
rect 35224 35992 35288 35996
rect 35224 35936 35228 35992
rect 35228 35936 35284 35992
rect 35284 35936 35288 35992
rect 35224 35932 35288 35936
rect 19624 35326 19688 35330
rect 19624 35270 19628 35326
rect 19628 35270 19684 35326
rect 19684 35270 19688 35326
rect 19624 35266 19688 35270
rect 19704 35326 19768 35330
rect 19704 35270 19708 35326
rect 19708 35270 19764 35326
rect 19764 35270 19768 35326
rect 19704 35266 19768 35270
rect 19784 35326 19848 35330
rect 19784 35270 19788 35326
rect 19788 35270 19844 35326
rect 19844 35270 19848 35326
rect 19784 35266 19848 35270
rect 19864 35326 19928 35330
rect 19864 35270 19868 35326
rect 19868 35270 19924 35326
rect 19924 35270 19928 35326
rect 19864 35266 19928 35270
rect 50344 35326 50408 35330
rect 50344 35270 50348 35326
rect 50348 35270 50404 35326
rect 50404 35270 50408 35326
rect 50344 35266 50408 35270
rect 50424 35326 50488 35330
rect 50424 35270 50428 35326
rect 50428 35270 50484 35326
rect 50484 35270 50488 35326
rect 50424 35266 50488 35270
rect 50504 35326 50568 35330
rect 50504 35270 50508 35326
rect 50508 35270 50564 35326
rect 50564 35270 50568 35326
rect 50504 35266 50568 35270
rect 50584 35326 50648 35330
rect 50584 35270 50588 35326
rect 50588 35270 50644 35326
rect 50644 35270 50648 35326
rect 50584 35266 50648 35270
rect 4264 34660 4328 34664
rect 4264 34604 4268 34660
rect 4268 34604 4324 34660
rect 4324 34604 4328 34660
rect 4264 34600 4328 34604
rect 4344 34660 4408 34664
rect 4344 34604 4348 34660
rect 4348 34604 4404 34660
rect 4404 34604 4408 34660
rect 4344 34600 4408 34604
rect 4424 34660 4488 34664
rect 4424 34604 4428 34660
rect 4428 34604 4484 34660
rect 4484 34604 4488 34660
rect 4424 34600 4488 34604
rect 4504 34660 4568 34664
rect 4504 34604 4508 34660
rect 4508 34604 4564 34660
rect 4564 34604 4568 34660
rect 4504 34600 4568 34604
rect 34984 34660 35048 34664
rect 34984 34604 34988 34660
rect 34988 34604 35044 34660
rect 35044 34604 35048 34660
rect 34984 34600 35048 34604
rect 35064 34660 35128 34664
rect 35064 34604 35068 34660
rect 35068 34604 35124 34660
rect 35124 34604 35128 34660
rect 35064 34600 35128 34604
rect 35144 34660 35208 34664
rect 35144 34604 35148 34660
rect 35148 34604 35204 34660
rect 35204 34604 35208 34660
rect 35144 34600 35208 34604
rect 35224 34660 35288 34664
rect 35224 34604 35228 34660
rect 35228 34604 35284 34660
rect 35284 34604 35288 34660
rect 35224 34600 35288 34604
rect 19624 33994 19688 33998
rect 19624 33938 19628 33994
rect 19628 33938 19684 33994
rect 19684 33938 19688 33994
rect 19624 33934 19688 33938
rect 19704 33994 19768 33998
rect 19704 33938 19708 33994
rect 19708 33938 19764 33994
rect 19764 33938 19768 33994
rect 19704 33934 19768 33938
rect 19784 33994 19848 33998
rect 19784 33938 19788 33994
rect 19788 33938 19844 33994
rect 19844 33938 19848 33994
rect 19784 33934 19848 33938
rect 19864 33994 19928 33998
rect 19864 33938 19868 33994
rect 19868 33938 19924 33994
rect 19924 33938 19928 33994
rect 19864 33934 19928 33938
rect 50344 33994 50408 33998
rect 50344 33938 50348 33994
rect 50348 33938 50404 33994
rect 50404 33938 50408 33994
rect 50344 33934 50408 33938
rect 50424 33994 50488 33998
rect 50424 33938 50428 33994
rect 50428 33938 50484 33994
rect 50484 33938 50488 33994
rect 50424 33934 50488 33938
rect 50504 33994 50568 33998
rect 50504 33938 50508 33994
rect 50508 33938 50564 33994
rect 50564 33938 50568 33994
rect 50504 33934 50568 33938
rect 50584 33994 50648 33998
rect 50584 33938 50588 33994
rect 50588 33938 50644 33994
rect 50644 33938 50648 33994
rect 50584 33934 50648 33938
rect 4264 33328 4328 33332
rect 4264 33272 4268 33328
rect 4268 33272 4324 33328
rect 4324 33272 4328 33328
rect 4264 33268 4328 33272
rect 4344 33328 4408 33332
rect 4344 33272 4348 33328
rect 4348 33272 4404 33328
rect 4404 33272 4408 33328
rect 4344 33268 4408 33272
rect 4424 33328 4488 33332
rect 4424 33272 4428 33328
rect 4428 33272 4484 33328
rect 4484 33272 4488 33328
rect 4424 33268 4488 33272
rect 4504 33328 4568 33332
rect 4504 33272 4508 33328
rect 4508 33272 4564 33328
rect 4564 33272 4568 33328
rect 4504 33268 4568 33272
rect 34984 33328 35048 33332
rect 34984 33272 34988 33328
rect 34988 33272 35044 33328
rect 35044 33272 35048 33328
rect 34984 33268 35048 33272
rect 35064 33328 35128 33332
rect 35064 33272 35068 33328
rect 35068 33272 35124 33328
rect 35124 33272 35128 33328
rect 35064 33268 35128 33272
rect 35144 33328 35208 33332
rect 35144 33272 35148 33328
rect 35148 33272 35204 33328
rect 35204 33272 35208 33328
rect 35144 33268 35208 33272
rect 35224 33328 35288 33332
rect 35224 33272 35228 33328
rect 35228 33272 35284 33328
rect 35284 33272 35288 33328
rect 35224 33268 35288 33272
rect 19624 32662 19688 32666
rect 19624 32606 19628 32662
rect 19628 32606 19684 32662
rect 19684 32606 19688 32662
rect 19624 32602 19688 32606
rect 19704 32662 19768 32666
rect 19704 32606 19708 32662
rect 19708 32606 19764 32662
rect 19764 32606 19768 32662
rect 19704 32602 19768 32606
rect 19784 32662 19848 32666
rect 19784 32606 19788 32662
rect 19788 32606 19844 32662
rect 19844 32606 19848 32662
rect 19784 32602 19848 32606
rect 19864 32662 19928 32666
rect 19864 32606 19868 32662
rect 19868 32606 19924 32662
rect 19924 32606 19928 32662
rect 19864 32602 19928 32606
rect 50344 32662 50408 32666
rect 50344 32606 50348 32662
rect 50348 32606 50404 32662
rect 50404 32606 50408 32662
rect 50344 32602 50408 32606
rect 50424 32662 50488 32666
rect 50424 32606 50428 32662
rect 50428 32606 50484 32662
rect 50484 32606 50488 32662
rect 50424 32602 50488 32606
rect 50504 32662 50568 32666
rect 50504 32606 50508 32662
rect 50508 32606 50564 32662
rect 50564 32606 50568 32662
rect 50504 32602 50568 32606
rect 50584 32662 50648 32666
rect 50584 32606 50588 32662
rect 50588 32606 50644 32662
rect 50644 32606 50648 32662
rect 50584 32602 50648 32606
rect 4264 31996 4328 32000
rect 4264 31940 4268 31996
rect 4268 31940 4324 31996
rect 4324 31940 4328 31996
rect 4264 31936 4328 31940
rect 4344 31996 4408 32000
rect 4344 31940 4348 31996
rect 4348 31940 4404 31996
rect 4404 31940 4408 31996
rect 4344 31936 4408 31940
rect 4424 31996 4488 32000
rect 4424 31940 4428 31996
rect 4428 31940 4484 31996
rect 4484 31940 4488 31996
rect 4424 31936 4488 31940
rect 4504 31996 4568 32000
rect 4504 31940 4508 31996
rect 4508 31940 4564 31996
rect 4564 31940 4568 31996
rect 4504 31936 4568 31940
rect 34984 31996 35048 32000
rect 34984 31940 34988 31996
rect 34988 31940 35044 31996
rect 35044 31940 35048 31996
rect 34984 31936 35048 31940
rect 35064 31996 35128 32000
rect 35064 31940 35068 31996
rect 35068 31940 35124 31996
rect 35124 31940 35128 31996
rect 35064 31936 35128 31940
rect 35144 31996 35208 32000
rect 35144 31940 35148 31996
rect 35148 31940 35204 31996
rect 35204 31940 35208 31996
rect 35144 31936 35208 31940
rect 35224 31996 35288 32000
rect 35224 31940 35228 31996
rect 35228 31940 35284 31996
rect 35284 31940 35288 31996
rect 35224 31936 35288 31940
rect 19624 31330 19688 31334
rect 19624 31274 19628 31330
rect 19628 31274 19684 31330
rect 19684 31274 19688 31330
rect 19624 31270 19688 31274
rect 19704 31330 19768 31334
rect 19704 31274 19708 31330
rect 19708 31274 19764 31330
rect 19764 31274 19768 31330
rect 19704 31270 19768 31274
rect 19784 31330 19848 31334
rect 19784 31274 19788 31330
rect 19788 31274 19844 31330
rect 19844 31274 19848 31330
rect 19784 31270 19848 31274
rect 19864 31330 19928 31334
rect 19864 31274 19868 31330
rect 19868 31274 19924 31330
rect 19924 31274 19928 31330
rect 19864 31270 19928 31274
rect 50344 31330 50408 31334
rect 50344 31274 50348 31330
rect 50348 31274 50404 31330
rect 50404 31274 50408 31330
rect 50344 31270 50408 31274
rect 50424 31330 50488 31334
rect 50424 31274 50428 31330
rect 50428 31274 50484 31330
rect 50484 31274 50488 31330
rect 50424 31270 50488 31274
rect 50504 31330 50568 31334
rect 50504 31274 50508 31330
rect 50508 31274 50564 31330
rect 50564 31274 50568 31330
rect 50504 31270 50568 31274
rect 50584 31330 50648 31334
rect 50584 31274 50588 31330
rect 50588 31274 50644 31330
rect 50644 31274 50648 31330
rect 50584 31270 50648 31274
rect 4264 30664 4328 30668
rect 4264 30608 4268 30664
rect 4268 30608 4324 30664
rect 4324 30608 4328 30664
rect 4264 30604 4328 30608
rect 4344 30664 4408 30668
rect 4344 30608 4348 30664
rect 4348 30608 4404 30664
rect 4404 30608 4408 30664
rect 4344 30604 4408 30608
rect 4424 30664 4488 30668
rect 4424 30608 4428 30664
rect 4428 30608 4484 30664
rect 4484 30608 4488 30664
rect 4424 30604 4488 30608
rect 4504 30664 4568 30668
rect 4504 30608 4508 30664
rect 4508 30608 4564 30664
rect 4564 30608 4568 30664
rect 4504 30604 4568 30608
rect 34984 30664 35048 30668
rect 34984 30608 34988 30664
rect 34988 30608 35044 30664
rect 35044 30608 35048 30664
rect 34984 30604 35048 30608
rect 35064 30664 35128 30668
rect 35064 30608 35068 30664
rect 35068 30608 35124 30664
rect 35124 30608 35128 30664
rect 35064 30604 35128 30608
rect 35144 30664 35208 30668
rect 35144 30608 35148 30664
rect 35148 30608 35204 30664
rect 35204 30608 35208 30664
rect 35144 30604 35208 30608
rect 35224 30664 35288 30668
rect 35224 30608 35228 30664
rect 35228 30608 35284 30664
rect 35284 30608 35288 30664
rect 35224 30604 35288 30608
rect 19624 29998 19688 30002
rect 19624 29942 19628 29998
rect 19628 29942 19684 29998
rect 19684 29942 19688 29998
rect 19624 29938 19688 29942
rect 19704 29998 19768 30002
rect 19704 29942 19708 29998
rect 19708 29942 19764 29998
rect 19764 29942 19768 29998
rect 19704 29938 19768 29942
rect 19784 29998 19848 30002
rect 19784 29942 19788 29998
rect 19788 29942 19844 29998
rect 19844 29942 19848 29998
rect 19784 29938 19848 29942
rect 19864 29998 19928 30002
rect 19864 29942 19868 29998
rect 19868 29942 19924 29998
rect 19924 29942 19928 29998
rect 19864 29938 19928 29942
rect 50344 29998 50408 30002
rect 50344 29942 50348 29998
rect 50348 29942 50404 29998
rect 50404 29942 50408 29998
rect 50344 29938 50408 29942
rect 50424 29998 50488 30002
rect 50424 29942 50428 29998
rect 50428 29942 50484 29998
rect 50484 29942 50488 29998
rect 50424 29938 50488 29942
rect 50504 29998 50568 30002
rect 50504 29942 50508 29998
rect 50508 29942 50564 29998
rect 50564 29942 50568 29998
rect 50504 29938 50568 29942
rect 50584 29998 50648 30002
rect 50584 29942 50588 29998
rect 50588 29942 50644 29998
rect 50644 29942 50648 29998
rect 50584 29938 50648 29942
rect 4264 29332 4328 29336
rect 4264 29276 4268 29332
rect 4268 29276 4324 29332
rect 4324 29276 4328 29332
rect 4264 29272 4328 29276
rect 4344 29332 4408 29336
rect 4344 29276 4348 29332
rect 4348 29276 4404 29332
rect 4404 29276 4408 29332
rect 4344 29272 4408 29276
rect 4424 29332 4488 29336
rect 4424 29276 4428 29332
rect 4428 29276 4484 29332
rect 4484 29276 4488 29332
rect 4424 29272 4488 29276
rect 4504 29332 4568 29336
rect 4504 29276 4508 29332
rect 4508 29276 4564 29332
rect 4564 29276 4568 29332
rect 4504 29272 4568 29276
rect 34984 29332 35048 29336
rect 34984 29276 34988 29332
rect 34988 29276 35044 29332
rect 35044 29276 35048 29332
rect 34984 29272 35048 29276
rect 35064 29332 35128 29336
rect 35064 29276 35068 29332
rect 35068 29276 35124 29332
rect 35124 29276 35128 29332
rect 35064 29272 35128 29276
rect 35144 29332 35208 29336
rect 35144 29276 35148 29332
rect 35148 29276 35204 29332
rect 35204 29276 35208 29332
rect 35144 29272 35208 29276
rect 35224 29332 35288 29336
rect 35224 29276 35228 29332
rect 35228 29276 35284 29332
rect 35284 29276 35288 29332
rect 35224 29272 35288 29276
rect 19624 28666 19688 28670
rect 19624 28610 19628 28666
rect 19628 28610 19684 28666
rect 19684 28610 19688 28666
rect 19624 28606 19688 28610
rect 19704 28666 19768 28670
rect 19704 28610 19708 28666
rect 19708 28610 19764 28666
rect 19764 28610 19768 28666
rect 19704 28606 19768 28610
rect 19784 28666 19848 28670
rect 19784 28610 19788 28666
rect 19788 28610 19844 28666
rect 19844 28610 19848 28666
rect 19784 28606 19848 28610
rect 19864 28666 19928 28670
rect 19864 28610 19868 28666
rect 19868 28610 19924 28666
rect 19924 28610 19928 28666
rect 19864 28606 19928 28610
rect 50344 28666 50408 28670
rect 50344 28610 50348 28666
rect 50348 28610 50404 28666
rect 50404 28610 50408 28666
rect 50344 28606 50408 28610
rect 50424 28666 50488 28670
rect 50424 28610 50428 28666
rect 50428 28610 50484 28666
rect 50484 28610 50488 28666
rect 50424 28606 50488 28610
rect 50504 28666 50568 28670
rect 50504 28610 50508 28666
rect 50508 28610 50564 28666
rect 50564 28610 50568 28666
rect 50504 28606 50568 28610
rect 50584 28666 50648 28670
rect 50584 28610 50588 28666
rect 50588 28610 50644 28666
rect 50644 28610 50648 28666
rect 50584 28606 50648 28610
rect 4264 28000 4328 28004
rect 4264 27944 4268 28000
rect 4268 27944 4324 28000
rect 4324 27944 4328 28000
rect 4264 27940 4328 27944
rect 4344 28000 4408 28004
rect 4344 27944 4348 28000
rect 4348 27944 4404 28000
rect 4404 27944 4408 28000
rect 4344 27940 4408 27944
rect 4424 28000 4488 28004
rect 4424 27944 4428 28000
rect 4428 27944 4484 28000
rect 4484 27944 4488 28000
rect 4424 27940 4488 27944
rect 4504 28000 4568 28004
rect 4504 27944 4508 28000
rect 4508 27944 4564 28000
rect 4564 27944 4568 28000
rect 4504 27940 4568 27944
rect 34984 28000 35048 28004
rect 34984 27944 34988 28000
rect 34988 27944 35044 28000
rect 35044 27944 35048 28000
rect 34984 27940 35048 27944
rect 35064 28000 35128 28004
rect 35064 27944 35068 28000
rect 35068 27944 35124 28000
rect 35124 27944 35128 28000
rect 35064 27940 35128 27944
rect 35144 28000 35208 28004
rect 35144 27944 35148 28000
rect 35148 27944 35204 28000
rect 35204 27944 35208 28000
rect 35144 27940 35208 27944
rect 35224 28000 35288 28004
rect 35224 27944 35228 28000
rect 35228 27944 35284 28000
rect 35284 27944 35288 28000
rect 35224 27940 35288 27944
rect 19624 27334 19688 27338
rect 19624 27278 19628 27334
rect 19628 27278 19684 27334
rect 19684 27278 19688 27334
rect 19624 27274 19688 27278
rect 19704 27334 19768 27338
rect 19704 27278 19708 27334
rect 19708 27278 19764 27334
rect 19764 27278 19768 27334
rect 19704 27274 19768 27278
rect 19784 27334 19848 27338
rect 19784 27278 19788 27334
rect 19788 27278 19844 27334
rect 19844 27278 19848 27334
rect 19784 27274 19848 27278
rect 19864 27334 19928 27338
rect 19864 27278 19868 27334
rect 19868 27278 19924 27334
rect 19924 27278 19928 27334
rect 19864 27274 19928 27278
rect 50344 27334 50408 27338
rect 50344 27278 50348 27334
rect 50348 27278 50404 27334
rect 50404 27278 50408 27334
rect 50344 27274 50408 27278
rect 50424 27334 50488 27338
rect 50424 27278 50428 27334
rect 50428 27278 50484 27334
rect 50484 27278 50488 27334
rect 50424 27274 50488 27278
rect 50504 27334 50568 27338
rect 50504 27278 50508 27334
rect 50508 27278 50564 27334
rect 50564 27278 50568 27334
rect 50504 27274 50568 27278
rect 50584 27334 50648 27338
rect 50584 27278 50588 27334
rect 50588 27278 50644 27334
rect 50644 27278 50648 27334
rect 50584 27274 50648 27278
rect 4264 26668 4328 26672
rect 4264 26612 4268 26668
rect 4268 26612 4324 26668
rect 4324 26612 4328 26668
rect 4264 26608 4328 26612
rect 4344 26668 4408 26672
rect 4344 26612 4348 26668
rect 4348 26612 4404 26668
rect 4404 26612 4408 26668
rect 4344 26608 4408 26612
rect 4424 26668 4488 26672
rect 4424 26612 4428 26668
rect 4428 26612 4484 26668
rect 4484 26612 4488 26668
rect 4424 26608 4488 26612
rect 4504 26668 4568 26672
rect 4504 26612 4508 26668
rect 4508 26612 4564 26668
rect 4564 26612 4568 26668
rect 4504 26608 4568 26612
rect 34984 26668 35048 26672
rect 34984 26612 34988 26668
rect 34988 26612 35044 26668
rect 35044 26612 35048 26668
rect 34984 26608 35048 26612
rect 35064 26668 35128 26672
rect 35064 26612 35068 26668
rect 35068 26612 35124 26668
rect 35124 26612 35128 26668
rect 35064 26608 35128 26612
rect 35144 26668 35208 26672
rect 35144 26612 35148 26668
rect 35148 26612 35204 26668
rect 35204 26612 35208 26668
rect 35144 26608 35208 26612
rect 35224 26668 35288 26672
rect 35224 26612 35228 26668
rect 35228 26612 35284 26668
rect 35284 26612 35288 26668
rect 35224 26608 35288 26612
rect 19624 26002 19688 26006
rect 19624 25946 19628 26002
rect 19628 25946 19684 26002
rect 19684 25946 19688 26002
rect 19624 25942 19688 25946
rect 19704 26002 19768 26006
rect 19704 25946 19708 26002
rect 19708 25946 19764 26002
rect 19764 25946 19768 26002
rect 19704 25942 19768 25946
rect 19784 26002 19848 26006
rect 19784 25946 19788 26002
rect 19788 25946 19844 26002
rect 19844 25946 19848 26002
rect 19784 25942 19848 25946
rect 19864 26002 19928 26006
rect 19864 25946 19868 26002
rect 19868 25946 19924 26002
rect 19924 25946 19928 26002
rect 19864 25942 19928 25946
rect 50344 26002 50408 26006
rect 50344 25946 50348 26002
rect 50348 25946 50404 26002
rect 50404 25946 50408 26002
rect 50344 25942 50408 25946
rect 50424 26002 50488 26006
rect 50424 25946 50428 26002
rect 50428 25946 50484 26002
rect 50484 25946 50488 26002
rect 50424 25942 50488 25946
rect 50504 26002 50568 26006
rect 50504 25946 50508 26002
rect 50508 25946 50564 26002
rect 50564 25946 50568 26002
rect 50504 25942 50568 25946
rect 50584 26002 50648 26006
rect 50584 25946 50588 26002
rect 50588 25946 50644 26002
rect 50644 25946 50648 26002
rect 50584 25942 50648 25946
rect 4264 25336 4328 25340
rect 4264 25280 4268 25336
rect 4268 25280 4324 25336
rect 4324 25280 4328 25336
rect 4264 25276 4328 25280
rect 4344 25336 4408 25340
rect 4344 25280 4348 25336
rect 4348 25280 4404 25336
rect 4404 25280 4408 25336
rect 4344 25276 4408 25280
rect 4424 25336 4488 25340
rect 4424 25280 4428 25336
rect 4428 25280 4484 25336
rect 4484 25280 4488 25336
rect 4424 25276 4488 25280
rect 4504 25336 4568 25340
rect 4504 25280 4508 25336
rect 4508 25280 4564 25336
rect 4564 25280 4568 25336
rect 4504 25276 4568 25280
rect 34984 25336 35048 25340
rect 34984 25280 34988 25336
rect 34988 25280 35044 25336
rect 35044 25280 35048 25336
rect 34984 25276 35048 25280
rect 35064 25336 35128 25340
rect 35064 25280 35068 25336
rect 35068 25280 35124 25336
rect 35124 25280 35128 25336
rect 35064 25276 35128 25280
rect 35144 25336 35208 25340
rect 35144 25280 35148 25336
rect 35148 25280 35204 25336
rect 35204 25280 35208 25336
rect 35144 25276 35208 25280
rect 35224 25336 35288 25340
rect 35224 25280 35228 25336
rect 35228 25280 35284 25336
rect 35284 25280 35288 25336
rect 35224 25276 35288 25280
rect 19624 24670 19688 24674
rect 19624 24614 19628 24670
rect 19628 24614 19684 24670
rect 19684 24614 19688 24670
rect 19624 24610 19688 24614
rect 19704 24670 19768 24674
rect 19704 24614 19708 24670
rect 19708 24614 19764 24670
rect 19764 24614 19768 24670
rect 19704 24610 19768 24614
rect 19784 24670 19848 24674
rect 19784 24614 19788 24670
rect 19788 24614 19844 24670
rect 19844 24614 19848 24670
rect 19784 24610 19848 24614
rect 19864 24670 19928 24674
rect 19864 24614 19868 24670
rect 19868 24614 19924 24670
rect 19924 24614 19928 24670
rect 19864 24610 19928 24614
rect 50344 24670 50408 24674
rect 50344 24614 50348 24670
rect 50348 24614 50404 24670
rect 50404 24614 50408 24670
rect 50344 24610 50408 24614
rect 50424 24670 50488 24674
rect 50424 24614 50428 24670
rect 50428 24614 50484 24670
rect 50484 24614 50488 24670
rect 50424 24610 50488 24614
rect 50504 24670 50568 24674
rect 50504 24614 50508 24670
rect 50508 24614 50564 24670
rect 50564 24614 50568 24670
rect 50504 24610 50568 24614
rect 50584 24670 50648 24674
rect 50584 24614 50588 24670
rect 50588 24614 50644 24670
rect 50644 24614 50648 24670
rect 50584 24610 50648 24614
rect 4264 24004 4328 24008
rect 4264 23948 4268 24004
rect 4268 23948 4324 24004
rect 4324 23948 4328 24004
rect 4264 23944 4328 23948
rect 4344 24004 4408 24008
rect 4344 23948 4348 24004
rect 4348 23948 4404 24004
rect 4404 23948 4408 24004
rect 4344 23944 4408 23948
rect 4424 24004 4488 24008
rect 4424 23948 4428 24004
rect 4428 23948 4484 24004
rect 4484 23948 4488 24004
rect 4424 23944 4488 23948
rect 4504 24004 4568 24008
rect 4504 23948 4508 24004
rect 4508 23948 4564 24004
rect 4564 23948 4568 24004
rect 4504 23944 4568 23948
rect 34984 24004 35048 24008
rect 34984 23948 34988 24004
rect 34988 23948 35044 24004
rect 35044 23948 35048 24004
rect 34984 23944 35048 23948
rect 35064 24004 35128 24008
rect 35064 23948 35068 24004
rect 35068 23948 35124 24004
rect 35124 23948 35128 24004
rect 35064 23944 35128 23948
rect 35144 24004 35208 24008
rect 35144 23948 35148 24004
rect 35148 23948 35204 24004
rect 35204 23948 35208 24004
rect 35144 23944 35208 23948
rect 35224 24004 35288 24008
rect 35224 23948 35228 24004
rect 35228 23948 35284 24004
rect 35284 23948 35288 24004
rect 35224 23944 35288 23948
rect 19624 23338 19688 23342
rect 19624 23282 19628 23338
rect 19628 23282 19684 23338
rect 19684 23282 19688 23338
rect 19624 23278 19688 23282
rect 19704 23338 19768 23342
rect 19704 23282 19708 23338
rect 19708 23282 19764 23338
rect 19764 23282 19768 23338
rect 19704 23278 19768 23282
rect 19784 23338 19848 23342
rect 19784 23282 19788 23338
rect 19788 23282 19844 23338
rect 19844 23282 19848 23338
rect 19784 23278 19848 23282
rect 19864 23338 19928 23342
rect 19864 23282 19868 23338
rect 19868 23282 19924 23338
rect 19924 23282 19928 23338
rect 19864 23278 19928 23282
rect 50344 23338 50408 23342
rect 50344 23282 50348 23338
rect 50348 23282 50404 23338
rect 50404 23282 50408 23338
rect 50344 23278 50408 23282
rect 50424 23338 50488 23342
rect 50424 23282 50428 23338
rect 50428 23282 50484 23338
rect 50484 23282 50488 23338
rect 50424 23278 50488 23282
rect 50504 23338 50568 23342
rect 50504 23282 50508 23338
rect 50508 23282 50564 23338
rect 50564 23282 50568 23338
rect 50504 23278 50568 23282
rect 50584 23338 50648 23342
rect 50584 23282 50588 23338
rect 50588 23282 50644 23338
rect 50644 23282 50648 23338
rect 50584 23278 50648 23282
rect 4264 22672 4328 22676
rect 4264 22616 4268 22672
rect 4268 22616 4324 22672
rect 4324 22616 4328 22672
rect 4264 22612 4328 22616
rect 4344 22672 4408 22676
rect 4344 22616 4348 22672
rect 4348 22616 4404 22672
rect 4404 22616 4408 22672
rect 4344 22612 4408 22616
rect 4424 22672 4488 22676
rect 4424 22616 4428 22672
rect 4428 22616 4484 22672
rect 4484 22616 4488 22672
rect 4424 22612 4488 22616
rect 4504 22672 4568 22676
rect 4504 22616 4508 22672
rect 4508 22616 4564 22672
rect 4564 22616 4568 22672
rect 4504 22612 4568 22616
rect 34984 22672 35048 22676
rect 34984 22616 34988 22672
rect 34988 22616 35044 22672
rect 35044 22616 35048 22672
rect 34984 22612 35048 22616
rect 35064 22672 35128 22676
rect 35064 22616 35068 22672
rect 35068 22616 35124 22672
rect 35124 22616 35128 22672
rect 35064 22612 35128 22616
rect 35144 22672 35208 22676
rect 35144 22616 35148 22672
rect 35148 22616 35204 22672
rect 35204 22616 35208 22672
rect 35144 22612 35208 22616
rect 35224 22672 35288 22676
rect 35224 22616 35228 22672
rect 35228 22616 35284 22672
rect 35284 22616 35288 22672
rect 35224 22612 35288 22616
rect 19624 22006 19688 22010
rect 19624 21950 19628 22006
rect 19628 21950 19684 22006
rect 19684 21950 19688 22006
rect 19624 21946 19688 21950
rect 19704 22006 19768 22010
rect 19704 21950 19708 22006
rect 19708 21950 19764 22006
rect 19764 21950 19768 22006
rect 19704 21946 19768 21950
rect 19784 22006 19848 22010
rect 19784 21950 19788 22006
rect 19788 21950 19844 22006
rect 19844 21950 19848 22006
rect 19784 21946 19848 21950
rect 19864 22006 19928 22010
rect 19864 21950 19868 22006
rect 19868 21950 19924 22006
rect 19924 21950 19928 22006
rect 19864 21946 19928 21950
rect 50344 22006 50408 22010
rect 50344 21950 50348 22006
rect 50348 21950 50404 22006
rect 50404 21950 50408 22006
rect 50344 21946 50408 21950
rect 50424 22006 50488 22010
rect 50424 21950 50428 22006
rect 50428 21950 50484 22006
rect 50484 21950 50488 22006
rect 50424 21946 50488 21950
rect 50504 22006 50568 22010
rect 50504 21950 50508 22006
rect 50508 21950 50564 22006
rect 50564 21950 50568 22006
rect 50504 21946 50568 21950
rect 50584 22006 50648 22010
rect 50584 21950 50588 22006
rect 50588 21950 50644 22006
rect 50644 21950 50648 22006
rect 50584 21946 50648 21950
rect 4264 21340 4328 21344
rect 4264 21284 4268 21340
rect 4268 21284 4324 21340
rect 4324 21284 4328 21340
rect 4264 21280 4328 21284
rect 4344 21340 4408 21344
rect 4344 21284 4348 21340
rect 4348 21284 4404 21340
rect 4404 21284 4408 21340
rect 4344 21280 4408 21284
rect 4424 21340 4488 21344
rect 4424 21284 4428 21340
rect 4428 21284 4484 21340
rect 4484 21284 4488 21340
rect 4424 21280 4488 21284
rect 4504 21340 4568 21344
rect 4504 21284 4508 21340
rect 4508 21284 4564 21340
rect 4564 21284 4568 21340
rect 4504 21280 4568 21284
rect 34984 21340 35048 21344
rect 34984 21284 34988 21340
rect 34988 21284 35044 21340
rect 35044 21284 35048 21340
rect 34984 21280 35048 21284
rect 35064 21340 35128 21344
rect 35064 21284 35068 21340
rect 35068 21284 35124 21340
rect 35124 21284 35128 21340
rect 35064 21280 35128 21284
rect 35144 21340 35208 21344
rect 35144 21284 35148 21340
rect 35148 21284 35204 21340
rect 35204 21284 35208 21340
rect 35144 21280 35208 21284
rect 35224 21340 35288 21344
rect 35224 21284 35228 21340
rect 35228 21284 35284 21340
rect 35284 21284 35288 21340
rect 35224 21280 35288 21284
rect 19624 20674 19688 20678
rect 19624 20618 19628 20674
rect 19628 20618 19684 20674
rect 19684 20618 19688 20674
rect 19624 20614 19688 20618
rect 19704 20674 19768 20678
rect 19704 20618 19708 20674
rect 19708 20618 19764 20674
rect 19764 20618 19768 20674
rect 19704 20614 19768 20618
rect 19784 20674 19848 20678
rect 19784 20618 19788 20674
rect 19788 20618 19844 20674
rect 19844 20618 19848 20674
rect 19784 20614 19848 20618
rect 19864 20674 19928 20678
rect 19864 20618 19868 20674
rect 19868 20618 19924 20674
rect 19924 20618 19928 20674
rect 19864 20614 19928 20618
rect 50344 20674 50408 20678
rect 50344 20618 50348 20674
rect 50348 20618 50404 20674
rect 50404 20618 50408 20674
rect 50344 20614 50408 20618
rect 50424 20674 50488 20678
rect 50424 20618 50428 20674
rect 50428 20618 50484 20674
rect 50484 20618 50488 20674
rect 50424 20614 50488 20618
rect 50504 20674 50568 20678
rect 50504 20618 50508 20674
rect 50508 20618 50564 20674
rect 50564 20618 50568 20674
rect 50504 20614 50568 20618
rect 50584 20674 50648 20678
rect 50584 20618 50588 20674
rect 50588 20618 50644 20674
rect 50644 20618 50648 20674
rect 50584 20614 50648 20618
rect 4264 20008 4328 20012
rect 4264 19952 4268 20008
rect 4268 19952 4324 20008
rect 4324 19952 4328 20008
rect 4264 19948 4328 19952
rect 4344 20008 4408 20012
rect 4344 19952 4348 20008
rect 4348 19952 4404 20008
rect 4404 19952 4408 20008
rect 4344 19948 4408 19952
rect 4424 20008 4488 20012
rect 4424 19952 4428 20008
rect 4428 19952 4484 20008
rect 4484 19952 4488 20008
rect 4424 19948 4488 19952
rect 4504 20008 4568 20012
rect 4504 19952 4508 20008
rect 4508 19952 4564 20008
rect 4564 19952 4568 20008
rect 4504 19948 4568 19952
rect 34984 20008 35048 20012
rect 34984 19952 34988 20008
rect 34988 19952 35044 20008
rect 35044 19952 35048 20008
rect 34984 19948 35048 19952
rect 35064 20008 35128 20012
rect 35064 19952 35068 20008
rect 35068 19952 35124 20008
rect 35124 19952 35128 20008
rect 35064 19948 35128 19952
rect 35144 20008 35208 20012
rect 35144 19952 35148 20008
rect 35148 19952 35204 20008
rect 35204 19952 35208 20008
rect 35144 19948 35208 19952
rect 35224 20008 35288 20012
rect 35224 19952 35228 20008
rect 35228 19952 35284 20008
rect 35284 19952 35288 20008
rect 35224 19948 35288 19952
rect 19624 19342 19688 19346
rect 19624 19286 19628 19342
rect 19628 19286 19684 19342
rect 19684 19286 19688 19342
rect 19624 19282 19688 19286
rect 19704 19342 19768 19346
rect 19704 19286 19708 19342
rect 19708 19286 19764 19342
rect 19764 19286 19768 19342
rect 19704 19282 19768 19286
rect 19784 19342 19848 19346
rect 19784 19286 19788 19342
rect 19788 19286 19844 19342
rect 19844 19286 19848 19342
rect 19784 19282 19848 19286
rect 19864 19342 19928 19346
rect 19864 19286 19868 19342
rect 19868 19286 19924 19342
rect 19924 19286 19928 19342
rect 19864 19282 19928 19286
rect 50344 19342 50408 19346
rect 50344 19286 50348 19342
rect 50348 19286 50404 19342
rect 50404 19286 50408 19342
rect 50344 19282 50408 19286
rect 50424 19342 50488 19346
rect 50424 19286 50428 19342
rect 50428 19286 50484 19342
rect 50484 19286 50488 19342
rect 50424 19282 50488 19286
rect 50504 19342 50568 19346
rect 50504 19286 50508 19342
rect 50508 19286 50564 19342
rect 50564 19286 50568 19342
rect 50504 19282 50568 19286
rect 50584 19342 50648 19346
rect 50584 19286 50588 19342
rect 50588 19286 50644 19342
rect 50644 19286 50648 19342
rect 50584 19282 50648 19286
rect 4264 18676 4328 18680
rect 4264 18620 4268 18676
rect 4268 18620 4324 18676
rect 4324 18620 4328 18676
rect 4264 18616 4328 18620
rect 4344 18676 4408 18680
rect 4344 18620 4348 18676
rect 4348 18620 4404 18676
rect 4404 18620 4408 18676
rect 4344 18616 4408 18620
rect 4424 18676 4488 18680
rect 4424 18620 4428 18676
rect 4428 18620 4484 18676
rect 4484 18620 4488 18676
rect 4424 18616 4488 18620
rect 4504 18676 4568 18680
rect 4504 18620 4508 18676
rect 4508 18620 4564 18676
rect 4564 18620 4568 18676
rect 4504 18616 4568 18620
rect 34984 18676 35048 18680
rect 34984 18620 34988 18676
rect 34988 18620 35044 18676
rect 35044 18620 35048 18676
rect 34984 18616 35048 18620
rect 35064 18676 35128 18680
rect 35064 18620 35068 18676
rect 35068 18620 35124 18676
rect 35124 18620 35128 18676
rect 35064 18616 35128 18620
rect 35144 18676 35208 18680
rect 35144 18620 35148 18676
rect 35148 18620 35204 18676
rect 35204 18620 35208 18676
rect 35144 18616 35208 18620
rect 35224 18676 35288 18680
rect 35224 18620 35228 18676
rect 35228 18620 35284 18676
rect 35284 18620 35288 18676
rect 35224 18616 35288 18620
rect 19624 18010 19688 18014
rect 19624 17954 19628 18010
rect 19628 17954 19684 18010
rect 19684 17954 19688 18010
rect 19624 17950 19688 17954
rect 19704 18010 19768 18014
rect 19704 17954 19708 18010
rect 19708 17954 19764 18010
rect 19764 17954 19768 18010
rect 19704 17950 19768 17954
rect 19784 18010 19848 18014
rect 19784 17954 19788 18010
rect 19788 17954 19844 18010
rect 19844 17954 19848 18010
rect 19784 17950 19848 17954
rect 19864 18010 19928 18014
rect 19864 17954 19868 18010
rect 19868 17954 19924 18010
rect 19924 17954 19928 18010
rect 19864 17950 19928 17954
rect 50344 18010 50408 18014
rect 50344 17954 50348 18010
rect 50348 17954 50404 18010
rect 50404 17954 50408 18010
rect 50344 17950 50408 17954
rect 50424 18010 50488 18014
rect 50424 17954 50428 18010
rect 50428 17954 50484 18010
rect 50484 17954 50488 18010
rect 50424 17950 50488 17954
rect 50504 18010 50568 18014
rect 50504 17954 50508 18010
rect 50508 17954 50564 18010
rect 50564 17954 50568 18010
rect 50504 17950 50568 17954
rect 50584 18010 50648 18014
rect 50584 17954 50588 18010
rect 50588 17954 50644 18010
rect 50644 17954 50648 18010
rect 50584 17950 50648 17954
rect 4264 17344 4328 17348
rect 4264 17288 4268 17344
rect 4268 17288 4324 17344
rect 4324 17288 4328 17344
rect 4264 17284 4328 17288
rect 4344 17344 4408 17348
rect 4344 17288 4348 17344
rect 4348 17288 4404 17344
rect 4404 17288 4408 17344
rect 4344 17284 4408 17288
rect 4424 17344 4488 17348
rect 4424 17288 4428 17344
rect 4428 17288 4484 17344
rect 4484 17288 4488 17344
rect 4424 17284 4488 17288
rect 4504 17344 4568 17348
rect 4504 17288 4508 17344
rect 4508 17288 4564 17344
rect 4564 17288 4568 17344
rect 4504 17284 4568 17288
rect 34984 17344 35048 17348
rect 34984 17288 34988 17344
rect 34988 17288 35044 17344
rect 35044 17288 35048 17344
rect 34984 17284 35048 17288
rect 35064 17344 35128 17348
rect 35064 17288 35068 17344
rect 35068 17288 35124 17344
rect 35124 17288 35128 17344
rect 35064 17284 35128 17288
rect 35144 17344 35208 17348
rect 35144 17288 35148 17344
rect 35148 17288 35204 17344
rect 35204 17288 35208 17344
rect 35144 17284 35208 17288
rect 35224 17344 35288 17348
rect 35224 17288 35228 17344
rect 35228 17288 35284 17344
rect 35284 17288 35288 17344
rect 35224 17284 35288 17288
rect 19624 16678 19688 16682
rect 19624 16622 19628 16678
rect 19628 16622 19684 16678
rect 19684 16622 19688 16678
rect 19624 16618 19688 16622
rect 19704 16678 19768 16682
rect 19704 16622 19708 16678
rect 19708 16622 19764 16678
rect 19764 16622 19768 16678
rect 19704 16618 19768 16622
rect 19784 16678 19848 16682
rect 19784 16622 19788 16678
rect 19788 16622 19844 16678
rect 19844 16622 19848 16678
rect 19784 16618 19848 16622
rect 19864 16678 19928 16682
rect 19864 16622 19868 16678
rect 19868 16622 19924 16678
rect 19924 16622 19928 16678
rect 19864 16618 19928 16622
rect 50344 16678 50408 16682
rect 50344 16622 50348 16678
rect 50348 16622 50404 16678
rect 50404 16622 50408 16678
rect 50344 16618 50408 16622
rect 50424 16678 50488 16682
rect 50424 16622 50428 16678
rect 50428 16622 50484 16678
rect 50484 16622 50488 16678
rect 50424 16618 50488 16622
rect 50504 16678 50568 16682
rect 50504 16622 50508 16678
rect 50508 16622 50564 16678
rect 50564 16622 50568 16678
rect 50504 16618 50568 16622
rect 50584 16678 50648 16682
rect 50584 16622 50588 16678
rect 50588 16622 50644 16678
rect 50644 16622 50648 16678
rect 50584 16618 50648 16622
rect 4264 16012 4328 16016
rect 4264 15956 4268 16012
rect 4268 15956 4324 16012
rect 4324 15956 4328 16012
rect 4264 15952 4328 15956
rect 4344 16012 4408 16016
rect 4344 15956 4348 16012
rect 4348 15956 4404 16012
rect 4404 15956 4408 16012
rect 4344 15952 4408 15956
rect 4424 16012 4488 16016
rect 4424 15956 4428 16012
rect 4428 15956 4484 16012
rect 4484 15956 4488 16012
rect 4424 15952 4488 15956
rect 4504 16012 4568 16016
rect 4504 15956 4508 16012
rect 4508 15956 4564 16012
rect 4564 15956 4568 16012
rect 4504 15952 4568 15956
rect 34984 16012 35048 16016
rect 34984 15956 34988 16012
rect 34988 15956 35044 16012
rect 35044 15956 35048 16012
rect 34984 15952 35048 15956
rect 35064 16012 35128 16016
rect 35064 15956 35068 16012
rect 35068 15956 35124 16012
rect 35124 15956 35128 16012
rect 35064 15952 35128 15956
rect 35144 16012 35208 16016
rect 35144 15956 35148 16012
rect 35148 15956 35204 16012
rect 35204 15956 35208 16012
rect 35144 15952 35208 15956
rect 35224 16012 35288 16016
rect 35224 15956 35228 16012
rect 35228 15956 35284 16012
rect 35284 15956 35288 16012
rect 35224 15952 35288 15956
rect 19624 15346 19688 15350
rect 19624 15290 19628 15346
rect 19628 15290 19684 15346
rect 19684 15290 19688 15346
rect 19624 15286 19688 15290
rect 19704 15346 19768 15350
rect 19704 15290 19708 15346
rect 19708 15290 19764 15346
rect 19764 15290 19768 15346
rect 19704 15286 19768 15290
rect 19784 15346 19848 15350
rect 19784 15290 19788 15346
rect 19788 15290 19844 15346
rect 19844 15290 19848 15346
rect 19784 15286 19848 15290
rect 19864 15346 19928 15350
rect 19864 15290 19868 15346
rect 19868 15290 19924 15346
rect 19924 15290 19928 15346
rect 19864 15286 19928 15290
rect 50344 15346 50408 15350
rect 50344 15290 50348 15346
rect 50348 15290 50404 15346
rect 50404 15290 50408 15346
rect 50344 15286 50408 15290
rect 50424 15346 50488 15350
rect 50424 15290 50428 15346
rect 50428 15290 50484 15346
rect 50484 15290 50488 15346
rect 50424 15286 50488 15290
rect 50504 15346 50568 15350
rect 50504 15290 50508 15346
rect 50508 15290 50564 15346
rect 50564 15290 50568 15346
rect 50504 15286 50568 15290
rect 50584 15346 50648 15350
rect 50584 15290 50588 15346
rect 50588 15290 50644 15346
rect 50644 15290 50648 15346
rect 50584 15286 50648 15290
rect 4264 14680 4328 14684
rect 4264 14624 4268 14680
rect 4268 14624 4324 14680
rect 4324 14624 4328 14680
rect 4264 14620 4328 14624
rect 4344 14680 4408 14684
rect 4344 14624 4348 14680
rect 4348 14624 4404 14680
rect 4404 14624 4408 14680
rect 4344 14620 4408 14624
rect 4424 14680 4488 14684
rect 4424 14624 4428 14680
rect 4428 14624 4484 14680
rect 4484 14624 4488 14680
rect 4424 14620 4488 14624
rect 4504 14680 4568 14684
rect 4504 14624 4508 14680
rect 4508 14624 4564 14680
rect 4564 14624 4568 14680
rect 4504 14620 4568 14624
rect 34984 14680 35048 14684
rect 34984 14624 34988 14680
rect 34988 14624 35044 14680
rect 35044 14624 35048 14680
rect 34984 14620 35048 14624
rect 35064 14680 35128 14684
rect 35064 14624 35068 14680
rect 35068 14624 35124 14680
rect 35124 14624 35128 14680
rect 35064 14620 35128 14624
rect 35144 14680 35208 14684
rect 35144 14624 35148 14680
rect 35148 14624 35204 14680
rect 35204 14624 35208 14680
rect 35144 14620 35208 14624
rect 35224 14680 35288 14684
rect 35224 14624 35228 14680
rect 35228 14624 35284 14680
rect 35284 14624 35288 14680
rect 35224 14620 35288 14624
rect 19624 14014 19688 14018
rect 19624 13958 19628 14014
rect 19628 13958 19684 14014
rect 19684 13958 19688 14014
rect 19624 13954 19688 13958
rect 19704 14014 19768 14018
rect 19704 13958 19708 14014
rect 19708 13958 19764 14014
rect 19764 13958 19768 14014
rect 19704 13954 19768 13958
rect 19784 14014 19848 14018
rect 19784 13958 19788 14014
rect 19788 13958 19844 14014
rect 19844 13958 19848 14014
rect 19784 13954 19848 13958
rect 19864 14014 19928 14018
rect 19864 13958 19868 14014
rect 19868 13958 19924 14014
rect 19924 13958 19928 14014
rect 19864 13954 19928 13958
rect 50344 14014 50408 14018
rect 50344 13958 50348 14014
rect 50348 13958 50404 14014
rect 50404 13958 50408 14014
rect 50344 13954 50408 13958
rect 50424 14014 50488 14018
rect 50424 13958 50428 14014
rect 50428 13958 50484 14014
rect 50484 13958 50488 14014
rect 50424 13954 50488 13958
rect 50504 14014 50568 14018
rect 50504 13958 50508 14014
rect 50508 13958 50564 14014
rect 50564 13958 50568 14014
rect 50504 13954 50568 13958
rect 50584 14014 50648 14018
rect 50584 13958 50588 14014
rect 50588 13958 50644 14014
rect 50644 13958 50648 14014
rect 50584 13954 50648 13958
rect 4264 13348 4328 13352
rect 4264 13292 4268 13348
rect 4268 13292 4324 13348
rect 4324 13292 4328 13348
rect 4264 13288 4328 13292
rect 4344 13348 4408 13352
rect 4344 13292 4348 13348
rect 4348 13292 4404 13348
rect 4404 13292 4408 13348
rect 4344 13288 4408 13292
rect 4424 13348 4488 13352
rect 4424 13292 4428 13348
rect 4428 13292 4484 13348
rect 4484 13292 4488 13348
rect 4424 13288 4488 13292
rect 4504 13348 4568 13352
rect 4504 13292 4508 13348
rect 4508 13292 4564 13348
rect 4564 13292 4568 13348
rect 4504 13288 4568 13292
rect 34984 13348 35048 13352
rect 34984 13292 34988 13348
rect 34988 13292 35044 13348
rect 35044 13292 35048 13348
rect 34984 13288 35048 13292
rect 35064 13348 35128 13352
rect 35064 13292 35068 13348
rect 35068 13292 35124 13348
rect 35124 13292 35128 13348
rect 35064 13288 35128 13292
rect 35144 13348 35208 13352
rect 35144 13292 35148 13348
rect 35148 13292 35204 13348
rect 35204 13292 35208 13348
rect 35144 13288 35208 13292
rect 35224 13348 35288 13352
rect 35224 13292 35228 13348
rect 35228 13292 35284 13348
rect 35284 13292 35288 13348
rect 35224 13288 35288 13292
rect 19624 12682 19688 12686
rect 19624 12626 19628 12682
rect 19628 12626 19684 12682
rect 19684 12626 19688 12682
rect 19624 12622 19688 12626
rect 19704 12682 19768 12686
rect 19704 12626 19708 12682
rect 19708 12626 19764 12682
rect 19764 12626 19768 12682
rect 19704 12622 19768 12626
rect 19784 12682 19848 12686
rect 19784 12626 19788 12682
rect 19788 12626 19844 12682
rect 19844 12626 19848 12682
rect 19784 12622 19848 12626
rect 19864 12682 19928 12686
rect 19864 12626 19868 12682
rect 19868 12626 19924 12682
rect 19924 12626 19928 12682
rect 19864 12622 19928 12626
rect 50344 12682 50408 12686
rect 50344 12626 50348 12682
rect 50348 12626 50404 12682
rect 50404 12626 50408 12682
rect 50344 12622 50408 12626
rect 50424 12682 50488 12686
rect 50424 12626 50428 12682
rect 50428 12626 50484 12682
rect 50484 12626 50488 12682
rect 50424 12622 50488 12626
rect 50504 12682 50568 12686
rect 50504 12626 50508 12682
rect 50508 12626 50564 12682
rect 50564 12626 50568 12682
rect 50504 12622 50568 12626
rect 50584 12682 50648 12686
rect 50584 12626 50588 12682
rect 50588 12626 50644 12682
rect 50644 12626 50648 12682
rect 50584 12622 50648 12626
rect 4264 12016 4328 12020
rect 4264 11960 4268 12016
rect 4268 11960 4324 12016
rect 4324 11960 4328 12016
rect 4264 11956 4328 11960
rect 4344 12016 4408 12020
rect 4344 11960 4348 12016
rect 4348 11960 4404 12016
rect 4404 11960 4408 12016
rect 4344 11956 4408 11960
rect 4424 12016 4488 12020
rect 4424 11960 4428 12016
rect 4428 11960 4484 12016
rect 4484 11960 4488 12016
rect 4424 11956 4488 11960
rect 4504 12016 4568 12020
rect 4504 11960 4508 12016
rect 4508 11960 4564 12016
rect 4564 11960 4568 12016
rect 4504 11956 4568 11960
rect 34984 12016 35048 12020
rect 34984 11960 34988 12016
rect 34988 11960 35044 12016
rect 35044 11960 35048 12016
rect 34984 11956 35048 11960
rect 35064 12016 35128 12020
rect 35064 11960 35068 12016
rect 35068 11960 35124 12016
rect 35124 11960 35128 12016
rect 35064 11956 35128 11960
rect 35144 12016 35208 12020
rect 35144 11960 35148 12016
rect 35148 11960 35204 12016
rect 35204 11960 35208 12016
rect 35144 11956 35208 11960
rect 35224 12016 35288 12020
rect 35224 11960 35228 12016
rect 35228 11960 35284 12016
rect 35284 11960 35288 12016
rect 35224 11956 35288 11960
rect 19624 11350 19688 11354
rect 19624 11294 19628 11350
rect 19628 11294 19684 11350
rect 19684 11294 19688 11350
rect 19624 11290 19688 11294
rect 19704 11350 19768 11354
rect 19704 11294 19708 11350
rect 19708 11294 19764 11350
rect 19764 11294 19768 11350
rect 19704 11290 19768 11294
rect 19784 11350 19848 11354
rect 19784 11294 19788 11350
rect 19788 11294 19844 11350
rect 19844 11294 19848 11350
rect 19784 11290 19848 11294
rect 19864 11350 19928 11354
rect 19864 11294 19868 11350
rect 19868 11294 19924 11350
rect 19924 11294 19928 11350
rect 19864 11290 19928 11294
rect 50344 11350 50408 11354
rect 50344 11294 50348 11350
rect 50348 11294 50404 11350
rect 50404 11294 50408 11350
rect 50344 11290 50408 11294
rect 50424 11350 50488 11354
rect 50424 11294 50428 11350
rect 50428 11294 50484 11350
rect 50484 11294 50488 11350
rect 50424 11290 50488 11294
rect 50504 11350 50568 11354
rect 50504 11294 50508 11350
rect 50508 11294 50564 11350
rect 50564 11294 50568 11350
rect 50504 11290 50568 11294
rect 50584 11350 50648 11354
rect 50584 11294 50588 11350
rect 50588 11294 50644 11350
rect 50644 11294 50648 11350
rect 50584 11290 50648 11294
rect 4264 10684 4328 10688
rect 4264 10628 4268 10684
rect 4268 10628 4324 10684
rect 4324 10628 4328 10684
rect 4264 10624 4328 10628
rect 4344 10684 4408 10688
rect 4344 10628 4348 10684
rect 4348 10628 4404 10684
rect 4404 10628 4408 10684
rect 4344 10624 4408 10628
rect 4424 10684 4488 10688
rect 4424 10628 4428 10684
rect 4428 10628 4484 10684
rect 4484 10628 4488 10684
rect 4424 10624 4488 10628
rect 4504 10684 4568 10688
rect 4504 10628 4508 10684
rect 4508 10628 4564 10684
rect 4564 10628 4568 10684
rect 4504 10624 4568 10628
rect 34984 10684 35048 10688
rect 34984 10628 34988 10684
rect 34988 10628 35044 10684
rect 35044 10628 35048 10684
rect 34984 10624 35048 10628
rect 35064 10684 35128 10688
rect 35064 10628 35068 10684
rect 35068 10628 35124 10684
rect 35124 10628 35128 10684
rect 35064 10624 35128 10628
rect 35144 10684 35208 10688
rect 35144 10628 35148 10684
rect 35148 10628 35204 10684
rect 35204 10628 35208 10684
rect 35144 10624 35208 10628
rect 35224 10684 35288 10688
rect 35224 10628 35228 10684
rect 35228 10628 35284 10684
rect 35284 10628 35288 10684
rect 35224 10624 35288 10628
rect 19624 10018 19688 10022
rect 19624 9962 19628 10018
rect 19628 9962 19684 10018
rect 19684 9962 19688 10018
rect 19624 9958 19688 9962
rect 19704 10018 19768 10022
rect 19704 9962 19708 10018
rect 19708 9962 19764 10018
rect 19764 9962 19768 10018
rect 19704 9958 19768 9962
rect 19784 10018 19848 10022
rect 19784 9962 19788 10018
rect 19788 9962 19844 10018
rect 19844 9962 19848 10018
rect 19784 9958 19848 9962
rect 19864 10018 19928 10022
rect 19864 9962 19868 10018
rect 19868 9962 19924 10018
rect 19924 9962 19928 10018
rect 19864 9958 19928 9962
rect 50344 10018 50408 10022
rect 50344 9962 50348 10018
rect 50348 9962 50404 10018
rect 50404 9962 50408 10018
rect 50344 9958 50408 9962
rect 50424 10018 50488 10022
rect 50424 9962 50428 10018
rect 50428 9962 50484 10018
rect 50484 9962 50488 10018
rect 50424 9958 50488 9962
rect 50504 10018 50568 10022
rect 50504 9962 50508 10018
rect 50508 9962 50564 10018
rect 50564 9962 50568 10018
rect 50504 9958 50568 9962
rect 50584 10018 50648 10022
rect 50584 9962 50588 10018
rect 50588 9962 50644 10018
rect 50644 9962 50648 10018
rect 50584 9958 50648 9962
rect 4264 9352 4328 9356
rect 4264 9296 4268 9352
rect 4268 9296 4324 9352
rect 4324 9296 4328 9352
rect 4264 9292 4328 9296
rect 4344 9352 4408 9356
rect 4344 9296 4348 9352
rect 4348 9296 4404 9352
rect 4404 9296 4408 9352
rect 4344 9292 4408 9296
rect 4424 9352 4488 9356
rect 4424 9296 4428 9352
rect 4428 9296 4484 9352
rect 4484 9296 4488 9352
rect 4424 9292 4488 9296
rect 4504 9352 4568 9356
rect 4504 9296 4508 9352
rect 4508 9296 4564 9352
rect 4564 9296 4568 9352
rect 4504 9292 4568 9296
rect 34984 9352 35048 9356
rect 34984 9296 34988 9352
rect 34988 9296 35044 9352
rect 35044 9296 35048 9352
rect 34984 9292 35048 9296
rect 35064 9352 35128 9356
rect 35064 9296 35068 9352
rect 35068 9296 35124 9352
rect 35124 9296 35128 9352
rect 35064 9292 35128 9296
rect 35144 9352 35208 9356
rect 35144 9296 35148 9352
rect 35148 9296 35204 9352
rect 35204 9296 35208 9352
rect 35144 9292 35208 9296
rect 35224 9352 35288 9356
rect 35224 9296 35228 9352
rect 35228 9296 35284 9352
rect 35284 9296 35288 9352
rect 35224 9292 35288 9296
rect 19624 8686 19688 8690
rect 19624 8630 19628 8686
rect 19628 8630 19684 8686
rect 19684 8630 19688 8686
rect 19624 8626 19688 8630
rect 19704 8686 19768 8690
rect 19704 8630 19708 8686
rect 19708 8630 19764 8686
rect 19764 8630 19768 8686
rect 19704 8626 19768 8630
rect 19784 8686 19848 8690
rect 19784 8630 19788 8686
rect 19788 8630 19844 8686
rect 19844 8630 19848 8686
rect 19784 8626 19848 8630
rect 19864 8686 19928 8690
rect 19864 8630 19868 8686
rect 19868 8630 19924 8686
rect 19924 8630 19928 8686
rect 19864 8626 19928 8630
rect 50344 8686 50408 8690
rect 50344 8630 50348 8686
rect 50348 8630 50404 8686
rect 50404 8630 50408 8686
rect 50344 8626 50408 8630
rect 50424 8686 50488 8690
rect 50424 8630 50428 8686
rect 50428 8630 50484 8686
rect 50484 8630 50488 8686
rect 50424 8626 50488 8630
rect 50504 8686 50568 8690
rect 50504 8630 50508 8686
rect 50508 8630 50564 8686
rect 50564 8630 50568 8686
rect 50504 8626 50568 8630
rect 50584 8686 50648 8690
rect 50584 8630 50588 8686
rect 50588 8630 50644 8686
rect 50644 8630 50648 8686
rect 50584 8626 50648 8630
rect 4264 8020 4328 8024
rect 4264 7964 4268 8020
rect 4268 7964 4324 8020
rect 4324 7964 4328 8020
rect 4264 7960 4328 7964
rect 4344 8020 4408 8024
rect 4344 7964 4348 8020
rect 4348 7964 4404 8020
rect 4404 7964 4408 8020
rect 4344 7960 4408 7964
rect 4424 8020 4488 8024
rect 4424 7964 4428 8020
rect 4428 7964 4484 8020
rect 4484 7964 4488 8020
rect 4424 7960 4488 7964
rect 4504 8020 4568 8024
rect 4504 7964 4508 8020
rect 4508 7964 4564 8020
rect 4564 7964 4568 8020
rect 4504 7960 4568 7964
rect 34984 8020 35048 8024
rect 34984 7964 34988 8020
rect 34988 7964 35044 8020
rect 35044 7964 35048 8020
rect 34984 7960 35048 7964
rect 35064 8020 35128 8024
rect 35064 7964 35068 8020
rect 35068 7964 35124 8020
rect 35124 7964 35128 8020
rect 35064 7960 35128 7964
rect 35144 8020 35208 8024
rect 35144 7964 35148 8020
rect 35148 7964 35204 8020
rect 35204 7964 35208 8020
rect 35144 7960 35208 7964
rect 35224 8020 35288 8024
rect 35224 7964 35228 8020
rect 35228 7964 35284 8020
rect 35284 7964 35288 8020
rect 35224 7960 35288 7964
rect 19624 7354 19688 7358
rect 19624 7298 19628 7354
rect 19628 7298 19684 7354
rect 19684 7298 19688 7354
rect 19624 7294 19688 7298
rect 19704 7354 19768 7358
rect 19704 7298 19708 7354
rect 19708 7298 19764 7354
rect 19764 7298 19768 7354
rect 19704 7294 19768 7298
rect 19784 7354 19848 7358
rect 19784 7298 19788 7354
rect 19788 7298 19844 7354
rect 19844 7298 19848 7354
rect 19784 7294 19848 7298
rect 19864 7354 19928 7358
rect 19864 7298 19868 7354
rect 19868 7298 19924 7354
rect 19924 7298 19928 7354
rect 19864 7294 19928 7298
rect 50344 7354 50408 7358
rect 50344 7298 50348 7354
rect 50348 7298 50404 7354
rect 50404 7298 50408 7354
rect 50344 7294 50408 7298
rect 50424 7354 50488 7358
rect 50424 7298 50428 7354
rect 50428 7298 50484 7354
rect 50484 7298 50488 7354
rect 50424 7294 50488 7298
rect 50504 7354 50568 7358
rect 50504 7298 50508 7354
rect 50508 7298 50564 7354
rect 50564 7298 50568 7354
rect 50504 7294 50568 7298
rect 50584 7354 50648 7358
rect 50584 7298 50588 7354
rect 50588 7298 50644 7354
rect 50644 7298 50648 7354
rect 50584 7294 50648 7298
rect 4264 6688 4328 6692
rect 4264 6632 4268 6688
rect 4268 6632 4324 6688
rect 4324 6632 4328 6688
rect 4264 6628 4328 6632
rect 4344 6688 4408 6692
rect 4344 6632 4348 6688
rect 4348 6632 4404 6688
rect 4404 6632 4408 6688
rect 4344 6628 4408 6632
rect 4424 6688 4488 6692
rect 4424 6632 4428 6688
rect 4428 6632 4484 6688
rect 4484 6632 4488 6688
rect 4424 6628 4488 6632
rect 4504 6688 4568 6692
rect 4504 6632 4508 6688
rect 4508 6632 4564 6688
rect 4564 6632 4568 6688
rect 4504 6628 4568 6632
rect 34984 6688 35048 6692
rect 34984 6632 34988 6688
rect 34988 6632 35044 6688
rect 35044 6632 35048 6688
rect 34984 6628 35048 6632
rect 35064 6688 35128 6692
rect 35064 6632 35068 6688
rect 35068 6632 35124 6688
rect 35124 6632 35128 6688
rect 35064 6628 35128 6632
rect 35144 6688 35208 6692
rect 35144 6632 35148 6688
rect 35148 6632 35204 6688
rect 35204 6632 35208 6688
rect 35144 6628 35208 6632
rect 35224 6688 35288 6692
rect 35224 6632 35228 6688
rect 35228 6632 35284 6688
rect 35284 6632 35288 6688
rect 35224 6628 35288 6632
rect 19624 6022 19688 6026
rect 19624 5966 19628 6022
rect 19628 5966 19684 6022
rect 19684 5966 19688 6022
rect 19624 5962 19688 5966
rect 19704 6022 19768 6026
rect 19704 5966 19708 6022
rect 19708 5966 19764 6022
rect 19764 5966 19768 6022
rect 19704 5962 19768 5966
rect 19784 6022 19848 6026
rect 19784 5966 19788 6022
rect 19788 5966 19844 6022
rect 19844 5966 19848 6022
rect 19784 5962 19848 5966
rect 19864 6022 19928 6026
rect 19864 5966 19868 6022
rect 19868 5966 19924 6022
rect 19924 5966 19928 6022
rect 19864 5962 19928 5966
rect 50344 6022 50408 6026
rect 50344 5966 50348 6022
rect 50348 5966 50404 6022
rect 50404 5966 50408 6022
rect 50344 5962 50408 5966
rect 50424 6022 50488 6026
rect 50424 5966 50428 6022
rect 50428 5966 50484 6022
rect 50484 5966 50488 6022
rect 50424 5962 50488 5966
rect 50504 6022 50568 6026
rect 50504 5966 50508 6022
rect 50508 5966 50564 6022
rect 50564 5966 50568 6022
rect 50504 5962 50568 5966
rect 50584 6022 50648 6026
rect 50584 5966 50588 6022
rect 50588 5966 50644 6022
rect 50644 5966 50648 6022
rect 50584 5962 50648 5966
rect 4264 5356 4328 5360
rect 4264 5300 4268 5356
rect 4268 5300 4324 5356
rect 4324 5300 4328 5356
rect 4264 5296 4328 5300
rect 4344 5356 4408 5360
rect 4344 5300 4348 5356
rect 4348 5300 4404 5356
rect 4404 5300 4408 5356
rect 4344 5296 4408 5300
rect 4424 5356 4488 5360
rect 4424 5300 4428 5356
rect 4428 5300 4484 5356
rect 4484 5300 4488 5356
rect 4424 5296 4488 5300
rect 4504 5356 4568 5360
rect 4504 5300 4508 5356
rect 4508 5300 4564 5356
rect 4564 5300 4568 5356
rect 4504 5296 4568 5300
rect 34984 5356 35048 5360
rect 34984 5300 34988 5356
rect 34988 5300 35044 5356
rect 35044 5300 35048 5356
rect 34984 5296 35048 5300
rect 35064 5356 35128 5360
rect 35064 5300 35068 5356
rect 35068 5300 35124 5356
rect 35124 5300 35128 5356
rect 35064 5296 35128 5300
rect 35144 5356 35208 5360
rect 35144 5300 35148 5356
rect 35148 5300 35204 5356
rect 35204 5300 35208 5356
rect 35144 5296 35208 5300
rect 35224 5356 35288 5360
rect 35224 5300 35228 5356
rect 35228 5300 35284 5356
rect 35284 5300 35288 5356
rect 35224 5296 35288 5300
rect 19624 4690 19688 4694
rect 19624 4634 19628 4690
rect 19628 4634 19684 4690
rect 19684 4634 19688 4690
rect 19624 4630 19688 4634
rect 19704 4690 19768 4694
rect 19704 4634 19708 4690
rect 19708 4634 19764 4690
rect 19764 4634 19768 4690
rect 19704 4630 19768 4634
rect 19784 4690 19848 4694
rect 19784 4634 19788 4690
rect 19788 4634 19844 4690
rect 19844 4634 19848 4690
rect 19784 4630 19848 4634
rect 19864 4690 19928 4694
rect 19864 4634 19868 4690
rect 19868 4634 19924 4690
rect 19924 4634 19928 4690
rect 19864 4630 19928 4634
rect 50344 4690 50408 4694
rect 50344 4634 50348 4690
rect 50348 4634 50404 4690
rect 50404 4634 50408 4690
rect 50344 4630 50408 4634
rect 50424 4690 50488 4694
rect 50424 4634 50428 4690
rect 50428 4634 50484 4690
rect 50484 4634 50488 4690
rect 50424 4630 50488 4634
rect 50504 4690 50568 4694
rect 50504 4634 50508 4690
rect 50508 4634 50564 4690
rect 50564 4634 50568 4690
rect 50504 4630 50568 4634
rect 50584 4690 50648 4694
rect 50584 4634 50588 4690
rect 50588 4634 50644 4690
rect 50644 4634 50648 4690
rect 50584 4630 50648 4634
rect 4264 4024 4328 4028
rect 4264 3968 4268 4024
rect 4268 3968 4324 4024
rect 4324 3968 4328 4024
rect 4264 3964 4328 3968
rect 4344 4024 4408 4028
rect 4344 3968 4348 4024
rect 4348 3968 4404 4024
rect 4404 3968 4408 4024
rect 4344 3964 4408 3968
rect 4424 4024 4488 4028
rect 4424 3968 4428 4024
rect 4428 3968 4484 4024
rect 4484 3968 4488 4024
rect 4424 3964 4488 3968
rect 4504 4024 4568 4028
rect 4504 3968 4508 4024
rect 4508 3968 4564 4024
rect 4564 3968 4568 4024
rect 4504 3964 4568 3968
rect 34984 4024 35048 4028
rect 34984 3968 34988 4024
rect 34988 3968 35044 4024
rect 35044 3968 35048 4024
rect 34984 3964 35048 3968
rect 35064 4024 35128 4028
rect 35064 3968 35068 4024
rect 35068 3968 35124 4024
rect 35124 3968 35128 4024
rect 35064 3964 35128 3968
rect 35144 4024 35208 4028
rect 35144 3968 35148 4024
rect 35148 3968 35204 4024
rect 35204 3968 35208 4024
rect 35144 3964 35208 3968
rect 35224 4024 35288 4028
rect 35224 3968 35228 4024
rect 35228 3968 35284 4024
rect 35284 3968 35288 4024
rect 35224 3964 35288 3968
rect 19624 3358 19688 3362
rect 19624 3302 19628 3358
rect 19628 3302 19684 3358
rect 19684 3302 19688 3358
rect 19624 3298 19688 3302
rect 19704 3358 19768 3362
rect 19704 3302 19708 3358
rect 19708 3302 19764 3358
rect 19764 3302 19768 3358
rect 19704 3298 19768 3302
rect 19784 3358 19848 3362
rect 19784 3302 19788 3358
rect 19788 3302 19844 3358
rect 19844 3302 19848 3358
rect 19784 3298 19848 3302
rect 19864 3358 19928 3362
rect 19864 3302 19868 3358
rect 19868 3302 19924 3358
rect 19924 3302 19928 3358
rect 19864 3298 19928 3302
rect 50344 3358 50408 3362
rect 50344 3302 50348 3358
rect 50348 3302 50404 3358
rect 50404 3302 50408 3358
rect 50344 3298 50408 3302
rect 50424 3358 50488 3362
rect 50424 3302 50428 3358
rect 50428 3302 50484 3358
rect 50484 3302 50488 3358
rect 50424 3298 50488 3302
rect 50504 3358 50568 3362
rect 50504 3302 50508 3358
rect 50508 3302 50564 3358
rect 50564 3302 50568 3358
rect 50504 3298 50568 3302
rect 50584 3358 50648 3362
rect 50584 3302 50588 3358
rect 50588 3302 50644 3358
rect 50644 3302 50648 3358
rect 50584 3298 50648 3302
rect 4264 2692 4328 2696
rect 4264 2636 4268 2692
rect 4268 2636 4324 2692
rect 4324 2636 4328 2692
rect 4264 2632 4328 2636
rect 4344 2692 4408 2696
rect 4344 2636 4348 2692
rect 4348 2636 4404 2692
rect 4404 2636 4408 2692
rect 4344 2632 4408 2636
rect 4424 2692 4488 2696
rect 4424 2636 4428 2692
rect 4428 2636 4484 2692
rect 4484 2636 4488 2692
rect 4424 2632 4488 2636
rect 4504 2692 4568 2696
rect 4504 2636 4508 2692
rect 4508 2636 4564 2692
rect 4564 2636 4568 2692
rect 4504 2632 4568 2636
rect 34984 2692 35048 2696
rect 34984 2636 34988 2692
rect 34988 2636 35044 2692
rect 35044 2636 35048 2692
rect 34984 2632 35048 2636
rect 35064 2692 35128 2696
rect 35064 2636 35068 2692
rect 35068 2636 35124 2692
rect 35124 2636 35128 2692
rect 35064 2632 35128 2636
rect 35144 2692 35208 2696
rect 35144 2636 35148 2692
rect 35148 2636 35204 2692
rect 35204 2636 35208 2692
rect 35144 2632 35208 2636
rect 35224 2692 35288 2696
rect 35224 2636 35228 2692
rect 35228 2636 35284 2692
rect 35284 2636 35288 2692
rect 35224 2632 35288 2636
<< metal4 >>
rect 4256 57308 4576 57324
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 55976 4576 57244
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 54644 4576 55912
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 53312 4576 54580
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 51980 4576 53248
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 50648 4576 51916
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 49316 4576 50584
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 47984 4576 49252
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 46652 4576 47920
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 45320 4576 46588
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 43988 4576 45256
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 42656 4576 43924
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 41324 4576 42592
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 39992 4576 41260
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 38660 4576 39928
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 37328 4576 38596
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 35996 4576 37264
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 34664 4576 35932
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 33332 4576 34600
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 32000 4576 33268
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 30668 4576 31936
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 29336 4576 30604
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 28004 4576 29272
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 26672 4576 27940
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 25340 4576 26608
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 24008 4576 25276
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 22676 4576 23944
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 21344 4576 22612
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 20012 4576 21280
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 18680 4576 19948
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 17348 4576 18616
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 16016 4576 17284
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 14684 4576 15952
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 13352 4576 14620
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 12020 4576 13288
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 10688 4576 11956
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 9356 4576 10624
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 8024 4576 9292
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 6692 4576 7960
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 5360 4576 6628
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 4028 4576 5296
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 2696 4576 3964
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 56642 19936 57324
rect 34976 57308 35296 57324
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 55310 19936 56578
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 53978 19936 55246
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 52646 19936 53914
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 51314 19936 52582
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 49982 19936 51250
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 48650 19936 49918
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 47318 19936 48586
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 45986 19936 47254
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 44654 19936 45922
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 43322 19936 44590
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 41990 19936 43258
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 40658 19936 41926
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 39326 19936 40594
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 37994 19936 39262
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 36662 19936 37930
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 35330 19936 36598
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 33998 19936 35266
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 32666 19936 33934
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 31334 19936 32602
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 30002 19936 31270
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 28670 19936 29938
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 27338 19936 28606
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 26006 19936 27274
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 24674 19936 25942
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 23342 19936 24610
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 22010 19936 23278
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 20678 19936 21946
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 19346 19936 20614
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 18014 19936 19282
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 16682 19936 17950
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 15350 19936 16618
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 14018 19936 15286
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 12686 19936 13954
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 11354 19936 12622
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 10022 19936 11290
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 8690 19936 9958
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 7358 19936 8626
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 6026 19936 7294
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 4694 19936 5962
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 3362 19936 4630
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 4256 2616 4576 2632
rect 19616 2616 19936 3298
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 55976 35296 57244
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 54644 35296 55912
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 53312 35296 54580
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 51980 35296 53248
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 50648 35296 51916
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 49316 35296 50584
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 47984 35296 49252
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 46652 35296 47920
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 45320 35296 46588
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 43988 35296 45256
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 42656 35296 43924
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 41324 35296 42592
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 39992 35296 41260
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 38660 35296 39928
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 37328 35296 38596
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 35996 35296 37264
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 34664 35296 35932
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 33332 35296 34600
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 32000 35296 33268
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 30668 35296 31936
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 29336 35296 30604
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 28004 35296 29272
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 26672 35296 27940
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 25340 35296 26608
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 24008 35296 25276
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 22676 35296 23944
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 21344 35296 22612
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 20012 35296 21280
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 18680 35296 19948
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 17348 35296 18616
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 16016 35296 17284
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 14684 35296 15952
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 13352 35296 14620
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 12020 35296 13288
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 10688 35296 11956
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 9356 35296 10624
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 8024 35296 9292
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 6692 35296 7960
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 5360 35296 6628
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 4028 35296 5296
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 2696 35296 3964
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 56642 50656 57324
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 55310 50656 56578
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 53978 50656 55246
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 52646 50656 53914
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 51314 50656 52582
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 49982 50656 51250
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 48650 50656 49918
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 47318 50656 48586
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 45986 50656 47254
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 44654 50656 45922
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 43322 50656 44590
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 41990 50656 43258
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 40658 50656 41926
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 39326 50656 40594
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 37994 50656 39262
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 36662 50656 37930
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 35330 50656 36598
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 33998 50656 35266
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 32666 50656 33934
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 31334 50656 32602
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 30002 50656 31270
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 28670 50656 29938
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 27338 50656 28606
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 26006 50656 27274
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 24674 50656 25942
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 23342 50656 24610
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 22010 50656 23278
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 20678 50656 21946
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 19346 50656 20614
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 18014 50656 19282
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 16682 50656 17950
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 15350 50656 16618
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 14018 50656 15286
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 12686 50656 13954
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 11354 50656 12622
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 10022 50656 11290
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 8690 50656 9958
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 7358 50656 8626
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 6026 50656 7294
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 4694 50656 5962
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 3362 50656 4630
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 34976 2616 35296 2632
rect 50336 2616 50656 3298
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
use sky130_fd_sc_ls__clkbuf_1  input296 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input295
timestamp 1621261055
transform 1 0 1536 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_0
timestamp 1621261055
transform 1 0 1152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_8
timestamp 1621261055
transform 1 0 1920 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_8
timestamp 1621261055
transform 1 0 1920 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input319
timestamp 1621261055
transform 1 0 2304 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input297
timestamp 1621261055
transform 1 0 2304 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_16
timestamp 1621261055
transform 1 0 2688 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_16
timestamp 1621261055
transform 1 0 2688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_24
timestamp 1621261055
transform 1 0 3456 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_24
timestamp 1621261055
transform 1 0 3456 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input323
timestamp 1621261055
transform 1 0 3072 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input322
timestamp 1621261055
transform 1 0 3072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_32
timestamp 1621261055
transform 1 0 4224 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3936 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input324
timestamp 1621261055
transform 1 0 3840 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_164 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3840 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_44 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 5376 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_40
timestamp 1621261055
transform 1 0 4992 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_43
timestamp 1621261055
transform 1 0 5280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_37
timestamp 1621261055
transform 1 0 4704 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input325
timestamp 1621261055
transform 1 0 4608 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input298
timestamp 1621261055
transform 1 0 4896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_50
timestamp 1621261055
transform 1 0 5952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_51
timestamp 1621261055
transform 1 0 6048 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input300
timestamp 1621261055
transform 1 0 5568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input299
timestamp 1621261055
transform 1 0 5664 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 6336 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_56
timestamp 1621261055
transform 1 0 6528 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_57
timestamp 1621261055
transform 1 0 6624 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_55
timestamp 1621261055
transform 1 0 6432 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_185
timestamp 1621261055
transform 1 0 6432 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_165
timestamp 1621261055
transform 1 0 6528 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input302
timestamp 1621261055
transform 1 0 6912 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input301
timestamp 1621261055
transform 1 0 7008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_64
timestamp 1621261055
transform 1 0 7296 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_65
timestamp 1621261055
transform 1 0 7392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input304
timestamp 1621261055
transform 1 0 7680 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_72
timestamp 1621261055
transform 1 0 8064 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_73
timestamp 1621261055
transform 1 0 8160 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input303
timestamp 1621261055
transform 1 0 7776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_12 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 8352 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input306
timestamp 1621261055
transform 1 0 8448 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _029_ $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 8544 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_80
timestamp 1621261055
transform 1 0 8832 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_80
timestamp 1621261055
transform 1 0 8832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_85
timestamp 1621261055
transform 1 0 9312 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input309
timestamp 1621261055
transform 1 0 9216 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_166
timestamp 1621261055
transform 1 0 9216 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_88
timestamp 1621261055
transform 1 0 9600 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input307
timestamp 1621261055
transform 1 0 9696 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_93
timestamp 1621261055
transform 1 0 10080 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input311
timestamp 1621261055
transform 1 0 9984 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_96
timestamp 1621261055
transform 1 0 10368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input313
timestamp 1621261055
transform 1 0 10752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input310
timestamp 1621261055
transform 1 0 10464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_104
timestamp 1621261055
transform 1 0 11136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_101
timestamp 1621261055
transform 1 0 10848 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _076_
timestamp 1621261055
transform 1 0 11232 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_108
timestamp 1621261055
transform 1 0 11520 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_108
timestamp 1621261055
transform 1 0 11520 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_111
timestamp 1621261055
transform 1 0 11808 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_113
timestamp 1621261055
transform 1 0 12000 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_186
timestamp 1621261055
transform 1 0 11712 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_167
timestamp 1621261055
transform 1 0 11904 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _172_
timestamp 1621261055
transform 1 0 12192 0 1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_118
timestamp 1621261055
transform 1 0 12480 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_121
timestamp 1621261055
transform 1 0 12768 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input167
timestamp 1621261055
transform 1 0 12864 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input39
timestamp 1621261055
transform 1 0 12960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_134
timestamp 1621261055
transform 1 0 14016 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_126
timestamp 1621261055
transform 1 0 13248 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_127
timestamp 1621261055
transform 1 0 13344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input89
timestamp 1621261055
transform 1 0 13632 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input78
timestamp 1621261055
transform 1 0 13728 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_135
timestamp 1621261055
transform 1 0 14112 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_142
timestamp 1621261055
transform 1 0 14784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_141
timestamp 1621261055
transform 1 0 14688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_139
timestamp 1621261055
transform 1 0 14496 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input100
timestamp 1621261055
transform 1 0 14400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_168
timestamp 1621261055
transform 1 0 14592 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_150
timestamp 1621261055
transform 1 0 15552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_149
timestamp 1621261055
transform 1 0 15456 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__buf_1  input122 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 15168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input111
timestamp 1621261055
transform 1 0 15072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_158
timestamp 1621261055
transform 1 0 16320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_159
timestamp 1621261055
transform 1 0 16416 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_157
timestamp 1621261055
transform 1 0 16224 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input133
timestamp 1621261055
transform 1 0 15936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input50
timestamp 1621261055
transform 1 0 16512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_162
timestamp 1621261055
transform 1 0 16704 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_166
timestamp 1621261055
transform 1 0 17088 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_164
timestamp 1621261055
transform 1 0 16896 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_169
timestamp 1621261055
transform 1 0 17376 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_164
timestamp 1621261055
transform 1 0 16896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input70
timestamp 1621261055
transform 1 0 17472 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_187
timestamp 1621261055
transform 1 0 16992 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_169
timestamp 1621261055
transform 1 0 17280 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_174
timestamp 1621261055
transform 1 0 17856 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_177
timestamp 1621261055
transform 1 0 18144 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input72
timestamp 1621261055
transform 1 0 18240 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input61
timestamp 1621261055
transform 1 0 17760 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_182
timestamp 1621261055
transform 1 0 18624 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_185
timestamp 1621261055
transform 1 0 18912 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input73
timestamp 1621261055
transform 1 0 19008 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input71
timestamp 1621261055
transform 1 0 18528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_190
timestamp 1621261055
transform 1 0 19392 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_197
timestamp 1621261055
transform 1 0 20064 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_195
timestamp 1621261055
transform 1 0 19872 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_193
timestamp 1621261055
transform 1 0 19680 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input75
timestamp 1621261055
transform 1 0 19776 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_170
timestamp 1621261055
transform 1 0 19968 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_206
timestamp 1621261055
transform 1 0 20928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_198
timestamp 1621261055
transform 1 0 20160 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_205
timestamp 1621261055
transform 1 0 20832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input77
timestamp 1621261055
transform 1 0 20544 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input74
timestamp 1621261055
transform 1 0 20448 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_214
timestamp 1621261055
transform 1 0 21696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_213
timestamp 1621261055
transform 1 0 21600 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input80
timestamp 1621261055
transform 1 0 21312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input76
timestamp 1621261055
transform 1 0 21216 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_218
timestamp 1621261055
transform 1 0 22080 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_188
timestamp 1621261055
transform 1 0 22272 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_221
timestamp 1621261055
transform 1 0 22368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_225
timestamp 1621261055
transform 1 0 22752 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_223
timestamp 1621261055
transform 1 0 22560 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_221
timestamp 1621261055
transform 1 0 22368 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input84
timestamp 1621261055
transform 1 0 22752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_171
timestamp 1621261055
transform 1 0 22656 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_229
timestamp 1621261055
transform 1 0 23136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input82
timestamp 1621261055
transform 1 0 23136 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_233
timestamp 1621261055
transform 1 0 23520 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input86
timestamp 1621261055
transform 1 0 23520 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_237
timestamp 1621261055
transform 1 0 23904 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input85
timestamp 1621261055
transform 1 0 23904 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_241
timestamp 1621261055
transform 1 0 24288 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_41
timestamp 1621261055
transform 1 0 24480 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input88
timestamp 1621261055
transform 1 0 24288 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_245
timestamp 1621261055
transform 1 0 24672 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _046_
timestamp 1621261055
transform 1 0 24672 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_248
timestamp 1621261055
transform 1 0 24960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input91
timestamp 1621261055
transform 1 0 25056 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_172
timestamp 1621261055
transform 1 0 25344 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_253
timestamp 1621261055
transform 1 0 25440 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_253
timestamp 1621261055
transform 1 0 25440 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input92
timestamp 1621261055
transform 1 0 25824 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input90
timestamp 1621261055
transform 1 0 25824 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_261
timestamp 1621261055
transform 1 0 26208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_261
timestamp 1621261055
transform 1 0 26208 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input95
timestamp 1621261055
transform 1 0 26592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input93
timestamp 1621261055
transform 1 0 26592 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_269
timestamp 1621261055
transform 1 0 26976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_269
timestamp 1621261055
transform 1 0 26976 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_273
timestamp 1621261055
transform 1 0 27360 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_45
timestamp 1621261055
transform 1 0 27168 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _047_
timestamp 1621261055
transform 1 0 27360 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_276
timestamp 1621261055
transform 1 0 27648 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_276
timestamp 1621261055
transform 1 0 27648 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_189
timestamp 1621261055
transform 1 0 27552 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_284
timestamp 1621261055
transform 1 0 28416 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_281
timestamp 1621261055
transform 1 0 28128 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input99
timestamp 1621261055
transform 1 0 28032 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_173
timestamp 1621261055
transform 1 0 28032 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_289
timestamp 1621261055
transform 1 0 28896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input102
timestamp 1621261055
transform 1 0 28800 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input98
timestamp 1621261055
transform 1 0 28512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_292
timestamp 1621261055
transform 1 0 29184 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input101
timestamp 1621261055
transform 1 0 29280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_297
timestamp 1621261055
transform 1 0 29664 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input104
timestamp 1621261055
transform 1 0 29568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_300
timestamp 1621261055
transform 1 0 29952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _111_
timestamp 1621261055
transform 1 0 30048 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_304
timestamp 1621261055
transform 1 0 30336 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input106
timestamp 1621261055
transform 1 0 30336 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_308
timestamp 1621261055
transform 1 0 30720 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_309
timestamp 1621261055
transform 1 0 30816 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_174
timestamp 1621261055
transform 1 0 30720 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_316
timestamp 1621261055
transform 1 0 31488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input108
timestamp 1621261055
transform 1 0 31104 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input107
timestamp 1621261055
transform 1 0 31200 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_317
timestamp 1621261055
transform 1 0 31584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input112
timestamp 1621261055
transform 1 0 31872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input109
timestamp 1621261055
transform 1 0 31968 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_324
timestamp 1621261055
transform 1 0 32256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_331
timestamp 1621261055
transform 1 0 32928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_328
timestamp 1621261055
transform 1 0 32640 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_325
timestamp 1621261055
transform 1 0 32352 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_190
timestamp 1621261055
transform 1 0 32832 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_339
timestamp 1621261055
transform 1 0 33696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_337
timestamp 1621261055
transform 1 0 33504 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_335
timestamp 1621261055
transform 1 0 33312 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_333
timestamp 1621261055
transform 1 0 33120 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input115
timestamp 1621261055
transform 1 0 33312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input114
timestamp 1621261055
transform 1 0 33888 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_175
timestamp 1621261055
transform 1 0 33408 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_347
timestamp 1621261055
transform 1 0 34464 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_345
timestamp 1621261055
transform 1 0 34272 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input118
timestamp 1621261055
transform 1 0 34080 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input117
timestamp 1621261055
transform 1 0 34656 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input120
timestamp 1621261055
transform 1 0 34848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_355
timestamp 1621261055
transform 1 0 35232 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_353
timestamp 1621261055
transform 1 0 35040 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input123
timestamp 1621261055
transform 1 0 35616 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_363
timestamp 1621261055
transform 1 0 36000 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_365
timestamp 1621261055
transform 1 0 36192 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_363
timestamp 1621261055
transform 1 0 36000 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_361
timestamp 1621261055
transform 1 0 35808 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input125
timestamp 1621261055
transform 1 0 36384 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_176
timestamp 1621261055
transform 1 0 36096 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_371
timestamp 1621261055
transform 1 0 36768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_373
timestamp 1621261055
transform 1 0 36960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input127
timestamp 1621261055
transform 1 0 37152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input126
timestamp 1621261055
transform 1 0 37344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input124
timestamp 1621261055
transform 1 0 36576 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_379
timestamp 1621261055
transform 1 0 37536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_381
timestamp 1621261055
transform 1 0 37728 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_386
timestamp 1621261055
transform 1 0 38208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_383
timestamp 1621261055
transform 1 0 37920 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_191
timestamp 1621261055
transform 1 0 38112 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _110_
timestamp 1621261055
transform 1 0 38112 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_388
timestamp 1621261055
transform 1 0 38400 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input131
timestamp 1621261055
transform 1 0 38592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_177
timestamp 1621261055
transform 1 0 38784 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_394
timestamp 1621261055
transform 1 0 38976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_393
timestamp 1621261055
transform 1 0 38880 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input130
timestamp 1621261055
transform 1 0 39264 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_402
timestamp 1621261055
transform 1 0 39744 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_401
timestamp 1621261055
transform 1 0 39648 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input134
timestamp 1621261055
transform 1 0 39360 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input132
timestamp 1621261055
transform 1 0 40032 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_409
timestamp 1621261055
transform 1 0 40416 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input136
timestamp 1621261055
transform 1 0 40128 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_410
timestamp 1621261055
transform 1 0 40512 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input138
timestamp 1621261055
transform 1 0 40896 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _180_
timestamp 1621261055
transform 1 0 40800 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_418
timestamp 1621261055
transform 1 0 41280 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_416
timestamp 1621261055
transform 1 0 41088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_421
timestamp 1621261055
transform 1 0 41568 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input140
timestamp 1621261055
transform 1 0 41664 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_178
timestamp 1621261055
transform 1 0 41472 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_426
timestamp 1621261055
transform 1 0 42048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_429
timestamp 1621261055
transform 1 0 42336 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input139
timestamp 1621261055
transform 1 0 41952 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input142
timestamp 1621261055
transform 1 0 42432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_438
timestamp 1621261055
transform 1 0 43200 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_434
timestamp 1621261055
transform 1 0 42816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_437
timestamp 1621261055
transform 1 0 43104 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input141
timestamp 1621261055
transform 1 0 42720 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_192
timestamp 1621261055
transform 1 0 43392 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_449
timestamp 1621261055
transform 1 0 44256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_441
timestamp 1621261055
transform 1 0 43488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_449
timestamp 1621261055
transform 1 0 44256 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_447
timestamp 1621261055
transform 1 0 44064 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_445
timestamp 1621261055
transform 1 0 43872 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input146
timestamp 1621261055
transform 1 0 43872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_179
timestamp 1621261055
transform 1 0 44160 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_457
timestamp 1621261055
transform 1 0 45024 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_457
timestamp 1621261055
transform 1 0 45024 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input149
timestamp 1621261055
transform 1 0 44640 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input147
timestamp 1621261055
transform 1 0 44640 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input151
timestamp 1621261055
transform 1 0 45408 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input150
timestamp 1621261055
transform 1 0 45408 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_465
timestamp 1621261055
transform 1 0 45792 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_465
timestamp 1621261055
transform 1 0 45792 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_473
timestamp 1621261055
transform 1 0 46560 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_472
timestamp 1621261055
transform 1 0 46464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input153
timestamp 1621261055
transform 1 0 46176 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _060_
timestamp 1621261055
transform 1 0 46176 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_477
timestamp 1621261055
transform 1 0 46944 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input156
timestamp 1621261055
transform 1 0 46944 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_180
timestamp 1621261055
transform 1 0 46848 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_481
timestamp 1621261055
transform 1 0 47328 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input154
timestamp 1621261055
transform 1 0 47328 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_485
timestamp 1621261055
transform 1 0 47712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input159
timestamp 1621261055
transform 1 0 47712 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_493
timestamp 1621261055
transform 1 0 48480 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_489
timestamp 1621261055
transform 1 0 48096 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_493
timestamp 1621261055
transform 1 0 48480 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input157
timestamp 1621261055
transform 1 0 48096 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_496
timestamp 1621261055
transform 1 0 48768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_500
timestamp 1621261055
transform 1 0 49152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input162
timestamp 1621261055
transform 1 0 49152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_193
timestamp 1621261055
transform 1 0 48672 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _181_
timestamp 1621261055
transform 1 0 48864 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_1_512
timestamp 1621261055
transform 1 0 50304 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_504
timestamp 1621261055
transform 1 0 49536 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_505
timestamp 1621261055
transform 1 0 49632 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input40
timestamp 1621261055
transform 1 0 50016 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_181
timestamp 1621261055
transform 1 0 49536 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_513
timestamp 1621261055
transform 1 0 50400 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input42
timestamp 1621261055
transform 1 0 50400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_517
timestamp 1621261055
transform 1 0 50784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_521
timestamp 1621261055
transform 1 0 51168 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input43
timestamp 1621261055
transform 1 0 51168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input41
timestamp 1621261055
transform 1 0 50784 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_525
timestamp 1621261055
transform 1 0 51552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_529
timestamp 1621261055
transform 1 0 51936 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input44
timestamp 1621261055
transform 1 0 51936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_533
timestamp 1621261055
transform 1 0 52320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_533
timestamp 1621261055
transform 1 0 52320 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_531
timestamp 1621261055
transform 1 0 52128 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input46
timestamp 1621261055
transform 1 0 52704 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input45
timestamp 1621261055
transform 1 0 52704 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_182
timestamp 1621261055
transform 1 0 52224 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_1_549
timestamp 1621261055
transform 1 0 53856 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_541
timestamp 1621261055
transform 1 0 53088 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_0_549
timestamp 1621261055
transform 1 0 53856 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_541
timestamp 1621261055
transform 1 0 53088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input47
timestamp 1621261055
transform 1 0 53472 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_551
timestamp 1621261055
transform 1 0 54048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_557
timestamp 1621261055
transform 1 0 54624 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input51
timestamp 1621261055
transform 1 0 54432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_194
timestamp 1621261055
transform 1 0 53952 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_559
timestamp 1621261055
transform 1 0 54816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_561
timestamp 1621261055
transform 1 0 55008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_559
timestamp 1621261055
transform 1 0 54816 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input54
timestamp 1621261055
transform 1 0 55200 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input52
timestamp 1621261055
transform 1 0 55392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_183
timestamp 1621261055
transform 1 0 54912 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_567
timestamp 1621261055
transform 1 0 55584 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_575
timestamp 1621261055
transform 1 0 56352 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_569
timestamp 1621261055
transform 1 0 55776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input56
timestamp 1621261055
transform 1 0 55968 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input55
timestamp 1621261055
transform 1 0 56160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_583
timestamp 1621261055
transform 1 0 57120 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_577
timestamp 1621261055
transform 1 0 56544 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input58
timestamp 1621261055
transform 1 0 56736 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_591
timestamp 1621261055
transform 1 0 57888 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_589
timestamp 1621261055
transform 1 0 57696 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_0_587
timestamp 1621261055
transform 1 0 57504 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_585
timestamp 1621261055
transform 1 0 57312 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input59
timestamp 1621261055
transform 1 0 57504 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_184
timestamp 1621261055
transform 1 0 57600 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_1
timestamp 1621261055
transform -1 0 58848 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_3
timestamp 1621261055
transform -1 0 58848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_595
timestamp 1621261055
transform 1 0 58272 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_4
timestamp 1621261055
transform 1 0 1152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input308
timestamp 1621261055
transform 1 0 1536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input330
timestamp 1621261055
transform 1 0 2304 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input341
timestamp 1621261055
transform 1 0 3072 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_8
timestamp 1621261055
transform 1 0 1920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_16
timestamp 1621261055
transform 1 0 2688 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_24
timestamp 1621261055
transform 1 0 3456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_195
timestamp 1621261055
transform 1 0 3840 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input326
timestamp 1621261055
transform 1 0 4320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input328
timestamp 1621261055
transform 1 0 5088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input331
timestamp 1621261055
transform 1 0 5856 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_29
timestamp 1621261055
transform 1 0 3936 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_37
timestamp 1621261055
transform 1 0 4704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_45
timestamp 1621261055
transform 1 0 5472 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_53
timestamp 1621261055
transform 1 0 6240 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input305
timestamp 1621261055
transform 1 0 7392 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input333
timestamp 1621261055
transform 1 0 6624 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input335
timestamp 1621261055
transform 1 0 8160 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_61
timestamp 1621261055
transform 1 0 7008 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_69
timestamp 1621261055
transform 1 0 7776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_77
timestamp 1621261055
transform 1 0 8544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_81
timestamp 1621261055
transform 1 0 8928 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_196
timestamp 1621261055
transform 1 0 9120 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input312
timestamp 1621261055
transform 1 0 9600 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input314
timestamp 1621261055
transform 1 0 10368 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input315
timestamp 1621261055
transform 1 0 11136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_84
timestamp 1621261055
transform 1 0 9216 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_92
timestamp 1621261055
transform 1 0 9984 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_100
timestamp 1621261055
transform 1 0 10752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_108
timestamp 1621261055
transform 1 0 11520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input206
timestamp 1621261055
transform 1 0 13536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input316
timestamp 1621261055
transform 1 0 11904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input317
timestamp 1621261055
transform 1 0 12672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_116
timestamp 1621261055
transform 1 0 12288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_124
timestamp 1621261055
transform 1 0 13056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_128
timestamp 1621261055
transform 1 0 13440 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_133
timestamp 1621261055
transform 1 0 13920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_197
timestamp 1621261055
transform 1 0 14400 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__buf_1  input144
timestamp 1621261055
transform 1 0 15456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input155
timestamp 1621261055
transform 1 0 16224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_137
timestamp 1621261055
transform 1 0 14304 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_139
timestamp 1621261055
transform 1 0 14496 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_147
timestamp 1621261055
transform 1 0 15264 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_153
timestamp 1621261055
transform 1 0 15840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_161
timestamp 1621261055
transform 1 0 16608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input166
timestamp 1621261055
transform 1 0 16992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input178
timestamp 1621261055
transform 1 0 17760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input198
timestamp 1621261055
transform 1 0 18528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_169
timestamp 1621261055
transform 1 0 17376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_177
timestamp 1621261055
transform 1 0 18144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_185
timestamp 1621261055
transform 1 0 18912 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_198
timestamp 1621261055
transform 1 0 19680 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input79
timestamp 1621261055
transform 1 0 20256 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input81
timestamp 1621261055
transform 1 0 21024 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input83
timestamp 1621261055
transform 1 0 21792 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_194
timestamp 1621261055
transform 1 0 19776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_198
timestamp 1621261055
transform 1 0 20160 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_203
timestamp 1621261055
transform 1 0 20640 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_211
timestamp 1621261055
transform 1 0 21408 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input87
timestamp 1621261055
transform 1 0 23232 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input211
timestamp 1621261055
transform 1 0 24000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_219
timestamp 1621261055
transform 1 0 22176 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_227
timestamp 1621261055
transform 1 0 22944 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_229
timestamp 1621261055
transform 1 0 23136 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_234
timestamp 1621261055
transform 1 0 23616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_242
timestamp 1621261055
transform 1 0 24384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_199
timestamp 1621261055
transform 1 0 24960 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input94
timestamp 1621261055
transform 1 0 25440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input96
timestamp 1621261055
transform 1 0 26208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input97
timestamp 1621261055
transform 1 0 26976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_246
timestamp 1621261055
transform 1 0 24768 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_249
timestamp 1621261055
transform 1 0 25056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_257
timestamp 1621261055
transform 1 0 25824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_265
timestamp 1621261055
transform 1 0 26592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input103
timestamp 1621261055
transform 1 0 28320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input105
timestamp 1621261055
transform 1 0 29088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_273
timestamp 1621261055
transform 1 0 27360 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_281
timestamp 1621261055
transform 1 0 28128 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_287
timestamp 1621261055
transform 1 0 28704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_295
timestamp 1621261055
transform 1 0 29472 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_200
timestamp 1621261055
transform 1 0 30240 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input110
timestamp 1621261055
transform 1 0 30912 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input113
timestamp 1621261055
transform 1 0 31680 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_304
timestamp 1621261055
transform 1 0 30336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_308
timestamp 1621261055
transform 1 0 30720 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_314
timestamp 1621261055
transform 1 0 31296 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_322
timestamp 1621261055
transform 1 0 32064 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input116
timestamp 1621261055
transform 1 0 32736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input119
timestamp 1621261055
transform 1 0 33888 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input121
timestamp 1621261055
transform 1 0 34656 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_326
timestamp 1621261055
transform 1 0 32448 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_328
timestamp 1621261055
transform 1 0 32640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_333
timestamp 1621261055
transform 1 0 33120 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_345
timestamp 1621261055
transform 1 0 34272 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_201
timestamp 1621261055
transform 1 0 35520 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input128
timestamp 1621261055
transform 1 0 36768 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input247
timestamp 1621261055
transform 1 0 36000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_353
timestamp 1621261055
transform 1 0 35040 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_357
timestamp 1621261055
transform 1 0 35424 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_359
timestamp 1621261055
transform 1 0 35616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_367
timestamp 1621261055
transform 1 0 36384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_375
timestamp 1621261055
transform 1 0 37152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input129
timestamp 1621261055
transform 1 0 37536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input135
timestamp 1621261055
transform 1 0 38976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input137
timestamp 1621261055
transform 1 0 39744 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_383
timestamp 1621261055
transform 1 0 37920 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_391
timestamp 1621261055
transform 1 0 38688 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_393
timestamp 1621261055
transform 1 0 38880 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_398
timestamp 1621261055
transform 1 0 39360 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _061_
timestamp 1621261055
transform 1 0 41280 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_202
timestamp 1621261055
transform 1 0 40800 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input143
timestamp 1621261055
transform 1 0 41952 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_406
timestamp 1621261055
transform 1 0 40128 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_410
timestamp 1621261055
transform 1 0 40512 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_412
timestamp 1621261055
transform 1 0 40704 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_414
timestamp 1621261055
transform 1 0 40896 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_421
timestamp 1621261055
transform 1 0 41568 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_429
timestamp 1621261055
transform 1 0 42336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _125_
timestamp 1621261055
transform 1 0 44256 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input145
timestamp 1621261055
transform 1 0 42720 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input148
timestamp 1621261055
transform 1 0 43488 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input152
timestamp 1621261055
transform 1 0 44928 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_437
timestamp 1621261055
transform 1 0 43104 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_445
timestamp 1621261055
transform 1 0 43872 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_452
timestamp 1621261055
transform 1 0 44544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_203
timestamp 1621261055
transform 1 0 46080 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input158
timestamp 1621261055
transform 1 0 46752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input160
timestamp 1621261055
transform 1 0 47520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_460
timestamp 1621261055
transform 1 0 45312 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_469
timestamp 1621261055
transform 1 0 46176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_473
timestamp 1621261055
transform 1 0 46560 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_479
timestamp 1621261055
transform 1 0 47136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input161
timestamp 1621261055
transform 1 0 48288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input163
timestamp 1621261055
transform 1 0 49056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input164
timestamp 1621261055
transform 1 0 49824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_487
timestamp 1621261055
transform 1 0 47904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_495
timestamp 1621261055
transform 1 0 48672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_503
timestamp 1621261055
transform 1 0 49440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_511
timestamp 1621261055
transform 1 0 50208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_204
timestamp 1621261055
transform 1 0 51360 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input48
timestamp 1621261055
transform 1 0 52608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input168
timestamp 1621261055
transform 1 0 50592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input171
timestamp 1621261055
transform 1 0 51840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_519
timestamp 1621261055
transform 1 0 50976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_524
timestamp 1621261055
transform 1 0 51456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_532
timestamp 1621261055
transform 1 0 52224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_540
timestamp 1621261055
transform 1 0 52992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input49
timestamp 1621261055
transform 1 0 53376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input53
timestamp 1621261055
transform 1 0 54144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input57
timestamp 1621261055
transform 1 0 55584 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_548
timestamp 1621261055
transform 1 0 53760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_556
timestamp 1621261055
transform 1 0 54528 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_564
timestamp 1621261055
transform 1 0 55296 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_566
timestamp 1621261055
transform 1 0 55488 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_205
timestamp 1621261055
transform 1 0 56640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input60
timestamp 1621261055
transform 1 0 57120 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_571
timestamp 1621261055
transform 1 0 55968 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_575
timestamp 1621261055
transform 1 0 56352 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_577
timestamp 1621261055
transform 1 0 56544 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_579
timestamp 1621261055
transform 1 0 56736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_587
timestamp 1621261055
transform 1 0 57504 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_5
timestamp 1621261055
transform -1 0 58848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_595
timestamp 1621261055
transform 1 0 58272 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_6
timestamp 1621261055
transform 1 0 1152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input329
timestamp 1621261055
transform 1 0 1536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input352
timestamp 1621261055
transform 1 0 2304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input355
timestamp 1621261055
transform 1 0 3072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_8
timestamp 1621261055
transform 1 0 1920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_16
timestamp 1621261055
transform 1 0 2688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_24
timestamp 1621261055
transform 1 0 3456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input327
timestamp 1621261055
transform 1 0 4128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input332
timestamp 1621261055
transform 1 0 5376 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_28
timestamp 1621261055
transform 1 0 3840 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_30
timestamp 1621261055
transform 1 0 4032 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_3_35
timestamp 1621261055
transform 1 0 4512 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_3_43
timestamp 1621261055
transform 1 0 5280 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_48
timestamp 1621261055
transform 1 0 5760 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_52
timestamp 1621261055
transform 1 0 6144 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_54
timestamp 1621261055
transform 1 0 6336 0 1 4662
box -38 -49 134 715
use AND2X1  AND2X1
timestamp 1624893035
transform 1 0 7680 0 1 4662
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_206
timestamp 1621261055
transform 1 0 6432 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input334
timestamp 1621261055
transform 1 0 6912 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_75
timestamp 1621261055
transform 1 0 7488 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_56
timestamp 1621261055
transform 1 0 6528 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_64
timestamp 1621261055
transform 1 0 7296 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_80
timestamp 1621261055
transform 1 0 8832 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input339
timestamp 1621261055
transform 1 0 9216 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input340
timestamp 1621261055
transform 1 0 9984 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input343
timestamp 1621261055
transform 1 0 10752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_88
timestamp 1621261055
transform 1 0 9600 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_96
timestamp 1621261055
transform 1 0 10368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_104
timestamp 1621261055
transform 1 0 11136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_108
timestamp 1621261055
transform 1 0 11520 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_207
timestamp 1621261055
transform 1 0 11712 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input217
timestamp 1621261055
transform 1 0 13920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input318
timestamp 1621261055
transform 1 0 12192 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input320
timestamp 1621261055
transform 1 0 12960 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_111
timestamp 1621261055
transform 1 0 11808 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_119
timestamp 1621261055
transform 1 0 12576 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_127
timestamp 1621261055
transform 1 0 13344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_131
timestamp 1621261055
transform 1 0 13728 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input228
timestamp 1621261055
transform 1 0 14688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input239
timestamp 1621261055
transform 1 0 15456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input261
timestamp 1621261055
transform 1 0 16224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_137
timestamp 1621261055
transform 1 0 14304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_145
timestamp 1621261055
transform 1 0 15072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_153
timestamp 1621261055
transform 1 0 15840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_161
timestamp 1621261055
transform 1 0 16608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_208
timestamp 1621261055
transform 1 0 16992 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input189
timestamp 1621261055
transform 1 0 17472 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input199
timestamp 1621261055
transform 1 0 18240 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input200
timestamp 1621261055
transform 1 0 19008 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_166
timestamp 1621261055
transform 1 0 17088 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_174
timestamp 1621261055
transform 1 0 17856 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_182
timestamp 1621261055
transform 1 0 18624 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input202
timestamp 1621261055
transform 1 0 19776 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input203
timestamp 1621261055
transform 1 0 20544 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input205
timestamp 1621261055
transform 1 0 21312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_190
timestamp 1621261055
transform 1 0 19392 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_198
timestamp 1621261055
transform 1 0 20160 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_206
timestamp 1621261055
transform 1 0 20928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_214
timestamp 1621261055
transform 1 0 21696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_209
timestamp 1621261055
transform 1 0 22272 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input209
timestamp 1621261055
transform 1 0 22752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input212
timestamp 1621261055
transform 1 0 23520 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input214
timestamp 1621261055
transform 1 0 24288 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_218
timestamp 1621261055
transform 1 0 22080 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_221
timestamp 1621261055
transform 1 0 22368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_229
timestamp 1621261055
transform 1 0 23136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_237
timestamp 1621261055
transform 1 0 23904 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input216
timestamp 1621261055
transform 1 0 25056 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input218
timestamp 1621261055
transform 1 0 25824 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input220
timestamp 1621261055
transform 1 0 26592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_245
timestamp 1621261055
transform 1 0 24672 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_253
timestamp 1621261055
transform 1 0 25440 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_261
timestamp 1621261055
transform 1 0 26208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_269
timestamp 1621261055
transform 1 0 26976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_210
timestamp 1621261055
transform 1 0 27552 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input224
timestamp 1621261055
transform 1 0 28032 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input227
timestamp 1621261055
transform 1 0 28800 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input230
timestamp 1621261055
transform 1 0 29568 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_273
timestamp 1621261055
transform 1 0 27360 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_276
timestamp 1621261055
transform 1 0 27648 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_284
timestamp 1621261055
transform 1 0 28416 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_292
timestamp 1621261055
transform 1 0 29184 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input232
timestamp 1621261055
transform 1 0 30336 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input233
timestamp 1621261055
transform 1 0 31104 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input236
timestamp 1621261055
transform 1 0 31872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_300
timestamp 1621261055
transform 1 0 29952 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_308
timestamp 1621261055
transform 1 0 30720 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_316
timestamp 1621261055
transform 1 0 31488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_324
timestamp 1621261055
transform 1 0 32256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_211
timestamp 1621261055
transform 1 0 32832 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input241
timestamp 1621261055
transform 1 0 33312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input243
timestamp 1621261055
transform 1 0 34080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input245
timestamp 1621261055
transform 1 0 34848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_328
timestamp 1621261055
transform 1 0 32640 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_331
timestamp 1621261055
transform 1 0 32928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_339
timestamp 1621261055
transform 1 0 33696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_347
timestamp 1621261055
transform 1 0 34464 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input248
timestamp 1621261055
transform 1 0 35616 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input249
timestamp 1621261055
transform 1 0 36384 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input252
timestamp 1621261055
transform 1 0 37152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_355
timestamp 1621261055
transform 1 0 35232 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_363
timestamp 1621261055
transform 1 0 36000 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_371
timestamp 1621261055
transform 1 0 36768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_212
timestamp 1621261055
transform 1 0 38112 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input256
timestamp 1621261055
transform 1 0 38592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input258
timestamp 1621261055
transform 1 0 39360 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_379
timestamp 1621261055
transform 1 0 37536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_383
timestamp 1621261055
transform 1 0 37920 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_386
timestamp 1621261055
transform 1 0 38208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_394
timestamp 1621261055
transform 1 0 38976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_402
timestamp 1621261055
transform 1 0 39744 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input260
timestamp 1621261055
transform 1 0 40128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input264
timestamp 1621261055
transform 1 0 40896 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input265
timestamp 1621261055
transform 1 0 41664 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input268
timestamp 1621261055
transform 1 0 42432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_410
timestamp 1621261055
transform 1 0 40512 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_418
timestamp 1621261055
transform 1 0 41280 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_426
timestamp 1621261055
transform 1 0 42048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_213
timestamp 1621261055
transform 1 0 43392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input273
timestamp 1621261055
transform 1 0 43872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input275
timestamp 1621261055
transform 1 0 44640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_434
timestamp 1621261055
transform 1 0 42816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_438
timestamp 1621261055
transform 1 0 43200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_441
timestamp 1621261055
transform 1 0 43488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_449
timestamp 1621261055
transform 1 0 44256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_457
timestamp 1621261055
transform 1 0 45024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input277
timestamp 1621261055
transform 1 0 45408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input279
timestamp 1621261055
transform 1 0 46176 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input280
timestamp 1621261055
transform 1 0 46944 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input284
timestamp 1621261055
transform 1 0 47712 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_465
timestamp 1621261055
transform 1 0 45792 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_473
timestamp 1621261055
transform 1 0 46560 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_481
timestamp 1621261055
transform 1 0 47328 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_214
timestamp 1621261055
transform 1 0 48672 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input165
timestamp 1621261055
transform 1 0 49344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input169
timestamp 1621261055
transform 1 0 50304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_489
timestamp 1621261055
transform 1 0 48096 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_493
timestamp 1621261055
transform 1 0 48480 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_496
timestamp 1621261055
transform 1 0 48768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_500
timestamp 1621261055
transform 1 0 49152 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_506
timestamp 1621261055
transform 1 0 49728 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_510
timestamp 1621261055
transform 1 0 50112 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input170
timestamp 1621261055
transform 1 0 51072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input172
timestamp 1621261055
transform 1 0 51840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input173
timestamp 1621261055
transform 1 0 52608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_516
timestamp 1621261055
transform 1 0 50688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_524
timestamp 1621261055
transform 1 0 51456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_532
timestamp 1621261055
transform 1 0 52224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_540
timestamp 1621261055
transform 1 0 52992 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_215
timestamp 1621261055
transform 1 0 53952 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input68
timestamp 1621261055
transform 1 0 55488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input177
timestamp 1621261055
transform 1 0 54432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_548
timestamp 1621261055
transform 1 0 53760 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_551
timestamp 1621261055
transform 1 0 54048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_559
timestamp 1621261055
transform 1 0 54816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_563
timestamp 1621261055
transform 1 0 55200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_565
timestamp 1621261055
transform 1 0 55392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input62
timestamp 1621261055
transform 1 0 57024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input64
timestamp 1621261055
transform 1 0 56256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_570
timestamp 1621261055
transform 1 0 55872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_578
timestamp 1621261055
transform 1 0 56640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_586
timestamp 1621261055
transform 1 0 57408 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_594
timestamp 1621261055
transform 1 0 58176 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_7
timestamp 1621261055
transform -1 0 58848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_596
timestamp 1621261055
transform 1 0 58368 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_8
timestamp 1621261055
transform 1 0 1152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input356
timestamp 1621261055
transform 1 0 2784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input362
timestamp 1621261055
transform 1 0 1536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_8
timestamp 1621261055
transform 1 0 1920 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_4_16
timestamp 1621261055
transform 1 0 2688 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_21
timestamp 1621261055
transform 1 0 3168 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_25
timestamp 1621261055
transform 1 0 3552 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_27
timestamp 1621261055
transform 1 0 3744 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_216
timestamp 1621261055
transform 1 0 3840 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input358
timestamp 1621261055
transform 1 0 4320 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input360
timestamp 1621261055
transform 1 0 5088 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output574 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 5856 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_223
timestamp 1621261055
transform 1 0 5664 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_29
timestamp 1621261055
transform 1 0 3936 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_37
timestamp 1621261055
transform 1 0 4704 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_45
timestamp 1621261055
transform 1 0 5472 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_53
timestamp 1621261055
transform 1 0 6240 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input336
timestamp 1621261055
transform 1 0 6816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input337
timestamp 1621261055
transform 1 0 7584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input338
timestamp 1621261055
transform 1 0 8352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_57
timestamp 1621261055
transform 1 0 6624 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_63
timestamp 1621261055
transform 1 0 7200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_71
timestamp 1621261055
transform 1 0 7968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_79
timestamp 1621261055
transform 1 0 8736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_217
timestamp 1621261055
transform 1 0 9120 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input342
timestamp 1621261055
transform 1 0 9600 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input345
timestamp 1621261055
transform 1 0 10368 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input347
timestamp 1621261055
transform 1 0 11136 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_84
timestamp 1621261055
transform 1 0 9216 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_92
timestamp 1621261055
transform 1 0 9984 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_100
timestamp 1621261055
transform 1 0 10752 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_108
timestamp 1621261055
transform 1 0 11520 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input321
timestamp 1621261055
transform 1 0 12576 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input351
timestamp 1621261055
transform 1 0 13344 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_116
timestamp 1621261055
transform 1 0 12288 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_118
timestamp 1621261055
transform 1 0 12480 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_123
timestamp 1621261055
transform 1 0 12960 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_131
timestamp 1621261055
transform 1 0 13728 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_135
timestamp 1621261055
transform 1 0 14112 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_218
timestamp 1621261055
transform 1 0 14400 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input250
timestamp 1621261055
transform 1 0 14976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input272
timestamp 1621261055
transform 1 0 15744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input283
timestamp 1621261055
transform 1 0 16512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_137
timestamp 1621261055
transform 1 0 14304 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_139
timestamp 1621261055
transform 1 0 14496 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_143
timestamp 1621261055
transform 1 0 14880 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_148
timestamp 1621261055
transform 1 0 15360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_156
timestamp 1621261055
transform 1 0 16128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input201
timestamp 1621261055
transform 1 0 18720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input294
timestamp 1621261055
transform 1 0 17280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_164
timestamp 1621261055
transform 1 0 16896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_4_172
timestamp 1621261055
transform 1 0 17664 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_180
timestamp 1621261055
transform 1 0 18432 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_182
timestamp 1621261055
transform 1 0 18624 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_187
timestamp 1621261055
transform 1 0 19104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_219
timestamp 1621261055
transform 1 0 19680 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input204
timestamp 1621261055
transform 1 0 20160 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input207
timestamp 1621261055
transform 1 0 20928 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input208
timestamp 1621261055
transform 1 0 21696 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_191
timestamp 1621261055
transform 1 0 19488 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_194
timestamp 1621261055
transform 1 0 19776 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_202
timestamp 1621261055
transform 1 0 20544 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_210
timestamp 1621261055
transform 1 0 21312 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input210
timestamp 1621261055
transform 1 0 22464 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input213
timestamp 1621261055
transform 1 0 23232 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input215
timestamp 1621261055
transform 1 0 24000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_218
timestamp 1621261055
transform 1 0 22080 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_226
timestamp 1621261055
transform 1 0 22848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_234
timestamp 1621261055
transform 1 0 23616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_242
timestamp 1621261055
transform 1 0 24384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_220
timestamp 1621261055
transform 1 0 24960 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input219
timestamp 1621261055
transform 1 0 25440 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input221
timestamp 1621261055
transform 1 0 26208 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input223
timestamp 1621261055
transform 1 0 26976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_246
timestamp 1621261055
transform 1 0 24768 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_249
timestamp 1621261055
transform 1 0 25056 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_257
timestamp 1621261055
transform 1 0 25824 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_265
timestamp 1621261055
transform 1 0 26592 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input226
timestamp 1621261055
transform 1 0 27744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input229
timestamp 1621261055
transform 1 0 28512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input231
timestamp 1621261055
transform 1 0 29280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_273
timestamp 1621261055
transform 1 0 27360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_281
timestamp 1621261055
transform 1 0 28128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_289
timestamp 1621261055
transform 1 0 28896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_297
timestamp 1621261055
transform 1 0 29664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_221
timestamp 1621261055
transform 1 0 30240 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input235
timestamp 1621261055
transform 1 0 30720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input237
timestamp 1621261055
transform 1 0 31488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input240
timestamp 1621261055
transform 1 0 32256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_301
timestamp 1621261055
transform 1 0 30048 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_304
timestamp 1621261055
transform 1 0 30336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_312
timestamp 1621261055
transform 1 0 31104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_320
timestamp 1621261055
transform 1 0 31872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input242
timestamp 1621261055
transform 1 0 33024 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input244
timestamp 1621261055
transform 1 0 33792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input246
timestamp 1621261055
transform 1 0 34560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_328
timestamp 1621261055
transform 1 0 32640 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_336
timestamp 1621261055
transform 1 0 33408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_344
timestamp 1621261055
transform 1 0 34176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_222
timestamp 1621261055
transform 1 0 35520 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input251
timestamp 1621261055
transform 1 0 36000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input253
timestamp 1621261055
transform 1 0 36768 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_352
timestamp 1621261055
transform 1 0 34944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_356
timestamp 1621261055
transform 1 0 35328 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_359
timestamp 1621261055
transform 1 0 35616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_367
timestamp 1621261055
transform 1 0 36384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_375
timestamp 1621261055
transform 1 0 37152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input255
timestamp 1621261055
transform 1 0 37536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input257
timestamp 1621261055
transform 1 0 38304 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input259
timestamp 1621261055
transform 1 0 39072 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input263
timestamp 1621261055
transform 1 0 39840 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_383
timestamp 1621261055
transform 1 0 37920 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_391
timestamp 1621261055
transform 1 0 38688 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_399
timestamp 1621261055
transform 1 0 39456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_223
timestamp 1621261055
transform 1 0 40800 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input267
timestamp 1621261055
transform 1 0 41280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input269
timestamp 1621261055
transform 1 0 42048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_407
timestamp 1621261055
transform 1 0 40224 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_411
timestamp 1621261055
transform 1 0 40608 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_414
timestamp 1621261055
transform 1 0 40896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_422
timestamp 1621261055
transform 1 0 41664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_430
timestamp 1621261055
transform 1 0 42432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input271
timestamp 1621261055
transform 1 0 42816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input274
timestamp 1621261055
transform 1 0 43584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input276
timestamp 1621261055
transform 1 0 44352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input278
timestamp 1621261055
transform 1 0 45120 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_438
timestamp 1621261055
transform 1 0 43200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_446
timestamp 1621261055
transform 1 0 43968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_454
timestamp 1621261055
transform 1 0 44736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_224
timestamp 1621261055
transform 1 0 46080 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input282
timestamp 1621261055
transform 1 0 46560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input285
timestamp 1621261055
transform 1 0 47328 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_462
timestamp 1621261055
transform 1 0 45504 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_466
timestamp 1621261055
transform 1 0 45888 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_469
timestamp 1621261055
transform 1 0 46176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_477
timestamp 1621261055
transform 1 0 46944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_485
timestamp 1621261055
transform 1 0 47712 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input287
timestamp 1621261055
transform 1 0 48096 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input289
timestamp 1621261055
transform 1 0 48864 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input290
timestamp 1621261055
transform 1 0 49632 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input292
timestamp 1621261055
transform 1 0 50400 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_493
timestamp 1621261055
transform 1 0 48480 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_501
timestamp 1621261055
transform 1 0 49248 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_509
timestamp 1621261055
transform 1 0 50016 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_225
timestamp 1621261055
transform 1 0 51360 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input174
timestamp 1621261055
transform 1 0 52128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input175
timestamp 1621261055
transform 1 0 52896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_517
timestamp 1621261055
transform 1 0 50784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_521
timestamp 1621261055
transform 1 0 51168 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_524
timestamp 1621261055
transform 1 0 51456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_528
timestamp 1621261055
transform 1 0 51840 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_530
timestamp 1621261055
transform 1 0 52032 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_535
timestamp 1621261055
transform 1 0 52512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _133_
timestamp 1621261055
transform 1 0 55200 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input176
timestamp 1621261055
transform 1 0 53664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input179
timestamp 1621261055
transform 1 0 54432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_543
timestamp 1621261055
transform 1 0 53280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_551
timestamp 1621261055
transform 1 0 54048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_559
timestamp 1621261055
transform 1 0 54816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_566
timestamp 1621261055
transform 1 0 55488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_226
timestamp 1621261055
transform 1 0 56640 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input63
timestamp 1621261055
transform 1 0 57408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input69
timestamp 1621261055
transform 1 0 55872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_574
timestamp 1621261055
transform 1 0 56256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_579
timestamp 1621261055
transform 1 0 56736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_583
timestamp 1621261055
transform 1 0 57120 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_4_585
timestamp 1621261055
transform 1 0 57312 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_590
timestamp 1621261055
transform 1 0 57792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_594
timestamp 1621261055
transform 1 0 58176 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_9
timestamp 1621261055
transform -1 0 58848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_596
timestamp 1621261055
transform 1 0 58368 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_10
timestamp 1621261055
transform 1 0 1152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input357
timestamp 1621261055
transform 1 0 3168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input363
timestamp 1621261055
transform 1 0 1536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input364
timestamp 1621261055
transform 1 0 2304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_8
timestamp 1621261055
transform 1 0 1920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_16
timestamp 1621261055
transform 1 0 2688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_20
timestamp 1621261055
transform 1 0 3072 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_25
timestamp 1621261055
transform 1 0 3552 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input359
timestamp 1621261055
transform 1 0 3936 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input361
timestamp 1621261055
transform 1 0 4704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output575
timestamp 1621261055
transform 1 0 5472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_225
timestamp 1621261055
transform 1 0 5280 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_33
timestamp 1621261055
transform 1 0 4320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_41
timestamp 1621261055
transform 1 0 5088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_49
timestamp 1621261055
transform 1 0 5856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_53
timestamp 1621261055
transform 1 0 6240 0 1 5994
box -38 -49 230 715
use AND2X2  AND2X2
timestamp 1624893035
transform 1 0 7680 0 1 5994
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_227
timestamp 1621261055
transform 1 0 6432 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output577
timestamp 1621261055
transform 1 0 6912 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_93
timestamp 1621261055
transform 1 0 7488 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_56
timestamp 1621261055
transform 1 0 6528 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_64
timestamp 1621261055
transform 1 0 7296 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_80
timestamp 1621261055
transform 1 0 8832 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input344
timestamp 1621261055
transform 1 0 9408 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input346
timestamp 1621261055
transform 1 0 10176 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input348
timestamp 1621261055
transform 1 0 10944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_84
timestamp 1621261055
transform 1 0 9216 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_90
timestamp 1621261055
transform 1 0 9792 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_98
timestamp 1621261055
transform 1 0 10560 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_106
timestamp 1621261055
transform 1 0 11328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_228
timestamp 1621261055
transform 1 0 11712 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input350
timestamp 1621261055
transform 1 0 12192 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input353
timestamp 1621261055
transform 1 0 12960 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output444
timestamp 1621261055
transform 1 0 13728 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_98
timestamp 1621261055
transform 1 0 13536 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_111
timestamp 1621261055
transform 1 0 11808 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_119
timestamp 1621261055
transform 1 0 12576 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_127
timestamp 1621261055
transform 1 0 13344 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_135
timestamp 1621261055
transform 1 0 14112 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output494
timestamp 1621261055
transform 1 0 14496 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output505
timestamp 1621261055
transform 1 0 15264 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output527
timestamp 1621261055
transform 1 0 16032 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_173
timestamp 1621261055
transform 1 0 15840 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_143
timestamp 1621261055
transform 1 0 14880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_151
timestamp 1621261055
transform 1 0 15648 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_159
timestamp 1621261055
transform 1 0 16416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_166
timestamp 1621261055
transform 1 0 17088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_163
timestamp 1621261055
transform 1 0 16800 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_229
timestamp 1621261055
transform 1 0 16992 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_112
timestamp 1621261055
transform 1 0 17280 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output455
timestamp 1621261055
transform 1 0 17472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_174
timestamp 1621261055
transform 1 0 17856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output475
timestamp 1621261055
transform 1 0 18240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_182
timestamp 1621261055
transform 1 0 18624 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_134
timestamp 1621261055
transform -1 0 19008 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output477
timestamp 1621261055
transform -1 0 19392 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output479
timestamp 1621261055
transform 1 0 19776 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output480
timestamp 1621261055
transform 1 0 20544 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output482
timestamp 1621261055
transform 1 0 21312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_136
timestamp 1621261055
transform 1 0 19584 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_190
timestamp 1621261055
transform 1 0 19392 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_198
timestamp 1621261055
transform 1 0 20160 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_206
timestamp 1621261055
transform 1 0 20928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_214
timestamp 1621261055
transform 1 0 21696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_230
timestamp 1621261055
transform 1 0 22272 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output487
timestamp 1621261055
transform 1 0 22752 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output489
timestamp 1621261055
transform 1 0 23520 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output491
timestamp 1621261055
transform 1 0 24288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_146
timestamp 1621261055
transform 1 0 24096 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_218
timestamp 1621261055
transform 1 0 22080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_221
timestamp 1621261055
transform 1 0 22368 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_229
timestamp 1621261055
transform 1 0 23136 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_237
timestamp 1621261055
transform 1 0 23904 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input222
timestamp 1621261055
transform 1 0 25632 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input225
timestamp 1621261055
transform 1 0 26784 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_245
timestamp 1621261055
transform 1 0 24672 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_253
timestamp 1621261055
transform 1 0 25440 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_259
timestamp 1621261055
transform 1 0 26016 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_231
timestamp 1621261055
transform 1 0 27552 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input234
timestamp 1621261055
transform 1 0 29664 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output501
timestamp 1621261055
transform 1 0 28032 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output504
timestamp 1621261055
transform 1 0 28800 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_271
timestamp 1621261055
transform 1 0 27168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_276
timestamp 1621261055
transform 1 0 27648 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_284
timestamp 1621261055
transform 1 0 28416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_292
timestamp 1621261055
transform 1 0 29184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_296
timestamp 1621261055
transform 1 0 29568 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input238
timestamp 1621261055
transform 1 0 31200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output509
timestamp 1621261055
transform -1 0 30816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output513
timestamp 1621261055
transform 1 0 31968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_160
timestamp 1621261055
transform -1 0 30432 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_164
timestamp 1621261055
transform 1 0 31776 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_301
timestamp 1621261055
transform 1 0 30048 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_309
timestamp 1621261055
transform 1 0 30816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_317
timestamp 1621261055
transform 1 0 31584 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_325
timestamp 1621261055
transform 1 0 32352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_331
timestamp 1621261055
transform 1 0 32928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_329
timestamp 1621261055
transform 1 0 32736 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_232
timestamp 1621261055
transform 1 0 32832 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output518
timestamp 1621261055
transform 1 0 33312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_339
timestamp 1621261055
transform 1 0 33696 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_170
timestamp 1621261055
transform -1 0 34080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output520
timestamp 1621261055
transform -1 0 34464 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_347
timestamp 1621261055
transform 1 0 34464 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_171
timestamp 1621261055
transform -1 0 34848 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output522
timestamp 1621261055
transform -1 0 35232 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input254
timestamp 1621261055
transform 1 0 36288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output529
timestamp 1621261055
transform 1 0 37056 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_175
timestamp 1621261055
transform 1 0 36864 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_355
timestamp 1621261055
transform 1 0 35232 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_363
timestamp 1621261055
transform 1 0 36000 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_365
timestamp 1621261055
transform 1 0 36192 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_370
timestamp 1621261055
transform 1 0 36672 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_378
timestamp 1621261055
transform 1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_382
timestamp 1621261055
transform 1 0 37824 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_386
timestamp 1621261055
transform 1 0 38208 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_384
timestamp 1621261055
transform 1 0 38016 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_233
timestamp 1621261055
transform 1 0 38112 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_5_392
timestamp 1621261055
transform 1 0 38784 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_390
timestamp 1621261055
transform 1 0 38592 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_397
timestamp 1621261055
transform 1 0 39264 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input262
timestamp 1621261055
transform 1 0 38880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _166_
timestamp 1621261055
transform 1 0 39648 0 1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_5_404
timestamp 1621261055
transform 1 0 39936 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input266
timestamp 1621261055
transform 1 0 40320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input270
timestamp 1621261055
transform 1 0 41856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output540
timestamp 1621261055
transform 1 0 41088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output544
timestamp 1621261055
transform -1 0 43008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_189
timestamp 1621261055
transform -1 0 42624 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_412
timestamp 1621261055
transform 1 0 40704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_420
timestamp 1621261055
transform 1 0 41472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_428
timestamp 1621261055
transform 1 0 42240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_234
timestamp 1621261055
transform 1 0 43392 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output548
timestamp 1621261055
transform 1 0 43872 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output552
timestamp 1621261055
transform 1 0 44640 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_436
timestamp 1621261055
transform 1 0 43008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_441
timestamp 1621261055
transform 1 0 43488 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_449
timestamp 1621261055
transform 1 0 44256 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_457
timestamp 1621261055
transform 1 0 45024 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input281
timestamp 1621261055
transform 1 0 45504 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input286
timestamp 1621261055
transform 1 0 46944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input288
timestamp 1621261055
transform 1 0 47712 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_461
timestamp 1621261055
transform 1 0 45408 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_5_466
timestamp 1621261055
transform 1 0 45888 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_474
timestamp 1621261055
transform 1 0 46656 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_476
timestamp 1621261055
transform 1 0 46848 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_481
timestamp 1621261055
transform 1 0 47328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_235
timestamp 1621261055
transform 1 0 48672 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input291
timestamp 1621261055
transform 1 0 49152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input293
timestamp 1621261055
transform 1 0 49920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_489
timestamp 1621261055
transform 1 0 48096 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_493
timestamp 1621261055
transform 1 0 48480 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_496
timestamp 1621261055
transform 1 0 48768 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_504
timestamp 1621261055
transform 1 0 49536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_512
timestamp 1621261055
transform 1 0 50304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output445
timestamp 1621261055
transform 1 0 50688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output447
timestamp 1621261055
transform -1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output448
timestamp 1621261055
transform 1 0 52224 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_102
timestamp 1621261055
transform -1 0 51456 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_520
timestamp 1621261055
transform 1 0 51072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_528
timestamp 1621261055
transform 1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_536
timestamp 1621261055
transform 1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_540
timestamp 1621261055
transform 1 0 52992 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_236
timestamp 1621261055
transform 1 0 53952 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input180
timestamp 1621261055
transform 1 0 54432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input181
timestamp 1621261055
transform 1 0 55200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input192
timestamp 1621261055
transform 1 0 53184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_546
timestamp 1621261055
transform 1 0 53568 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_551
timestamp 1621261055
transform 1 0 54048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_559
timestamp 1621261055
transform 1 0 54816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_567
timestamp 1621261055
transform 1 0 55584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input65
timestamp 1621261055
transform 1 0 57696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input67
timestamp 1621261055
transform 1 0 56928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input183
timestamp 1621261055
transform 1 0 55968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_575
timestamp 1621261055
transform 1 0 56352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_579
timestamp 1621261055
transform 1 0 56736 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_585
timestamp 1621261055
transform 1 0 57312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_593
timestamp 1621261055
transform 1 0 58080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_11
timestamp 1621261055
transform -1 0 58848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_12
timestamp 1621261055
transform 1 0 1152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input365
timestamp 1621261055
transform 1 0 2496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input366
timestamp 1621261055
transform 1 0 1536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_8
timestamp 1621261055
transform 1 0 1920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_12
timestamp 1621261055
transform 1 0 2304 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_18
timestamp 1621261055
transform 1 0 2880 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_26
timestamp 1621261055
transform 1 0 3648 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_29
timestamp 1621261055
transform 1 0 3936 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_237
timestamp 1621261055
transform 1 0 3840 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output598
timestamp 1621261055
transform 1 0 4320 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_37
timestamp 1621261055
transform 1 0 4704 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_250
timestamp 1621261055
transform 1 0 4896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output601
timestamp 1621261055
transform 1 0 5088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_45
timestamp 1621261055
transform 1 0 5472 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_227
timestamp 1621261055
transform 1 0 5664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output576
timestamp 1621261055
transform 1 0 5856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_53
timestamp 1621261055
transform 1 0 6240 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output578
timestamp 1621261055
transform 1 0 6624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output579
timestamp 1621261055
transform 1 0 7392 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output580
timestamp 1621261055
transform 1 0 8160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_228
timestamp 1621261055
transform 1 0 6432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_230
timestamp 1621261055
transform 1 0 7968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_61
timestamp 1621261055
transform 1 0 7008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_69
timestamp 1621261055
transform 1 0 7776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_77
timestamp 1621261055
transform 1 0 8544 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_81
timestamp 1621261055
transform 1 0 8928 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_238
timestamp 1621261055
transform 1 0 9120 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input349
timestamp 1621261055
transform 1 0 11232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output582
timestamp 1621261055
transform 1 0 9600 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output585
timestamp 1621261055
transform 1 0 10368 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_236
timestamp 1621261055
transform 1 0 10176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_84
timestamp 1621261055
transform 1 0 9216 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_92
timestamp 1621261055
transform 1 0 9984 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_100
timestamp 1621261055
transform 1 0 10752 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_104
timestamp 1621261055
transform 1 0 11136 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input354
timestamp 1621261055
transform 1 0 12672 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output483
timestamp 1621261055
transform 1 0 13440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_109
timestamp 1621261055
transform 1 0 11616 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_117
timestamp 1621261055
transform 1 0 12384 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_119
timestamp 1621261055
transform 1 0 12576 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_124
timestamp 1621261055
transform 1 0 13056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_132
timestamp 1621261055
transform 1 0 13824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_239
timestamp 1621261055
transform 1 0 14400 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output516
timestamp 1621261055
transform 1 0 14880 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output538
timestamp 1621261055
transform 1 0 15648 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_136
timestamp 1621261055
transform 1 0 14208 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_139
timestamp 1621261055
transform 1 0 14496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_147
timestamp 1621261055
transform 1 0 15264 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_155
timestamp 1621261055
transform 1 0 16032 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output466
timestamp 1621261055
transform 1 0 17088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output476
timestamp 1621261055
transform 1 0 17856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output478
timestamp 1621261055
transform 1 0 18624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_124
timestamp 1621261055
transform 1 0 16896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_132
timestamp 1621261055
transform 1 0 17664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_163
timestamp 1621261055
transform 1 0 16800 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_170
timestamp 1621261055
transform 1 0 17472 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_178
timestamp 1621261055
transform 1 0 18240 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_186
timestamp 1621261055
transform 1 0 19008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_192
timestamp 1621261055
transform 1 0 19584 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_190
timestamp 1621261055
transform 1 0 19392 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_240
timestamp 1621261055
transform 1 0 19680 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_194
timestamp 1621261055
transform 1 0 19776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_138
timestamp 1621261055
transform 1 0 19968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output481
timestamp 1621261055
transform 1 0 20160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_202
timestamp 1621261055
transform 1 0 20544 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_140
timestamp 1621261055
transform -1 0 20928 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output484
timestamp 1621261055
transform -1 0 21312 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_210
timestamp 1621261055
transform 1 0 21312 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output486
timestamp 1621261055
transform 1 0 21696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output488
timestamp 1621261055
transform 1 0 22464 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output490
timestamp 1621261055
transform 1 0 23232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output492
timestamp 1621261055
transform 1 0 24000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_144
timestamp 1621261055
transform 1 0 22272 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_148
timestamp 1621261055
transform 1 0 23808 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_218
timestamp 1621261055
transform 1 0 22080 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_226
timestamp 1621261055
transform 1 0 22848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_234
timestamp 1621261055
transform 1 0 23616 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_242
timestamp 1621261055
transform 1 0 24384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_241
timestamp 1621261055
transform 1 0 24960 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output496
timestamp 1621261055
transform 1 0 25440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output498
timestamp 1621261055
transform 1 0 26208 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output500
timestamp 1621261055
transform -1 0 27360 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_152
timestamp 1621261055
transform -1 0 26976 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_246
timestamp 1621261055
transform 1 0 24768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_249
timestamp 1621261055
transform 1 0 25056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_257
timestamp 1621261055
transform 1 0 25824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_265
timestamp 1621261055
transform 1 0 26592 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output503
timestamp 1621261055
transform 1 0 27744 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output506
timestamp 1621261055
transform 1 0 28512 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output508
timestamp 1621261055
transform -1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_154
timestamp 1621261055
transform 1 0 27552 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_158
timestamp 1621261055
transform -1 0 29280 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_273
timestamp 1621261055
transform 1 0 27360 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_281
timestamp 1621261055
transform 1 0 28128 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_289
timestamp 1621261055
transform 1 0 28896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_297
timestamp 1621261055
transform 1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_242
timestamp 1621261055
transform 1 0 30240 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output512
timestamp 1621261055
transform 1 0 30720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output514
timestamp 1621261055
transform 1 0 31488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output517
timestamp 1621261055
transform -1 0 32640 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_166
timestamp 1621261055
transform -1 0 32256 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_301
timestamp 1621261055
transform 1 0 30048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_304
timestamp 1621261055
transform 1 0 30336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_312
timestamp 1621261055
transform 1 0 31104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_320
timestamp 1621261055
transform 1 0 31872 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output519
timestamp 1621261055
transform 1 0 33024 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output521
timestamp 1621261055
transform 1 0 33792 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output524
timestamp 1621261055
transform 1 0 34560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_168
timestamp 1621261055
transform 1 0 32832 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_328
timestamp 1621261055
transform 1 0 32640 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_336
timestamp 1621261055
transform 1 0 33408 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_344
timestamp 1621261055
transform 1 0 34176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_352
timestamp 1621261055
transform 1 0 34944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_359
timestamp 1621261055
transform 1 0 35616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_356
timestamp 1621261055
transform 1 0 35328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_243
timestamp 1621261055
transform 1 0 35520 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output528
timestamp 1621261055
transform 1 0 36000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_367
timestamp 1621261055
transform 1 0 36384 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_177
timestamp 1621261055
transform -1 0 36768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_375
timestamp 1621261055
transform 1 0 37152 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output531
timestamp 1621261055
transform -1 0 37152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_181
timestamp 1621261055
transform 1 0 37344 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output533
timestamp 1621261055
transform 1 0 37536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output534
timestamp 1621261055
transform 1 0 38304 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output535
timestamp 1621261055
transform 1 0 39072 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output537
timestamp 1621261055
transform -1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_183
timestamp 1621261055
transform -1 0 39840 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_383
timestamp 1621261055
transform 1 0 37920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_391
timestamp 1621261055
transform 1 0 38688 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_399
timestamp 1621261055
transform 1 0 39456 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_407
timestamp 1621261055
transform 1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_414
timestamp 1621261055
transform 1 0 40896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_411
timestamp 1621261055
transform 1 0 40608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_244
timestamp 1621261055
transform 1 0 40800 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_185
timestamp 1621261055
transform -1 0 41280 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output542
timestamp 1621261055
transform -1 0 41664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_422
timestamp 1621261055
transform 1 0 41664 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_191
timestamp 1621261055
transform -1 0 42048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output545
timestamp 1621261055
transform -1 0 42432 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_430
timestamp 1621261055
transform 1 0 42432 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_192
timestamp 1621261055
transform -1 0 42816 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output547
timestamp 1621261055
transform -1 0 43200 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_438
timestamp 1621261055
transform 1 0 43200 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_196
timestamp 1621261055
transform 1 0 43392 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_446
timestamp 1621261055
transform 1 0 43968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output551
timestamp 1621261055
transform 1 0 43584 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_198
timestamp 1621261055
transform 1 0 44160 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output553
timestamp 1621261055
transform 1 0 44352 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_454
timestamp 1621261055
transform 1 0 44736 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_200
timestamp 1621261055
transform -1 0 45120 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output555
timestamp 1621261055
transform -1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_245
timestamp 1621261055
transform 1 0 46080 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output558
timestamp 1621261055
transform -1 0 46944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output561
timestamp 1621261055
transform 1 0 47328 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_204
timestamp 1621261055
transform -1 0 46560 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_462
timestamp 1621261055
transform 1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_466
timestamp 1621261055
transform 1 0 45888 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_469
timestamp 1621261055
transform 1 0 46176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_477
timestamp 1621261055
transform 1 0 46944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_485
timestamp 1621261055
transform 1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output446
timestamp 1621261055
transform -1 0 50496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output563
timestamp 1621261055
transform 1 0 48096 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output565
timestamp 1621261055
transform -1 0 49248 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_100
timestamp 1621261055
transform -1 0 50112 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_210
timestamp 1621261055
transform -1 0 48864 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_493
timestamp 1621261055
transform 1 0 48480 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_501
timestamp 1621261055
transform 1 0 49248 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_505
timestamp 1621261055
transform 1 0 49632 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_507
timestamp 1621261055
transform 1 0 49824 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_246
timestamp 1621261055
transform 1 0 51360 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output449
timestamp 1621261055
transform 1 0 51840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output451
timestamp 1621261055
transform -1 0 52992 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_106
timestamp 1621261055
transform -1 0 52608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_514
timestamp 1621261055
transform 1 0 50496 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_6_522
timestamp 1621261055
transform 1 0 51264 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_524
timestamp 1621261055
transform 1 0 51456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_532
timestamp 1621261055
transform 1 0 52224 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_540
timestamp 1621261055
transform 1 0 52992 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input182
timestamp 1621261055
transform 1 0 54720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input184
timestamp 1621261055
transform 1 0 55488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input196
timestamp 1621261055
transform 1 0 53952 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_548
timestamp 1621261055
transform 1 0 53760 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_554
timestamp 1621261055
transform 1 0 54336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_562
timestamp 1621261055
transform 1 0 55104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_247
timestamp 1621261055
transform 1 0 56640 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input66
timestamp 1621261055
transform 1 0 57696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_570
timestamp 1621261055
transform 1 0 55872 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_6_579
timestamp 1621261055
transform 1 0 56736 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_587
timestamp 1621261055
transform 1 0 57504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_593
timestamp 1621261055
transform 1 0 58080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_13
timestamp 1621261055
transform -1 0 58848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output572
timestamp 1621261055
transform 1 0 1536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input367
timestamp 1621261055
transform 1 0 1536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_16
timestamp 1621261055
transform 1 0 1152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_14
timestamp 1621261055
transform 1 0 1152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_8
timestamp 1621261055
transform 1 0 1920 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_219
timestamp 1621261055
transform 1 0 1920 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_10
timestamp 1621261055
transform 1 0 2112 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_221
timestamp 1621261055
transform 1 0 2112 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output584
timestamp 1621261055
transform 1 0 2304 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output573
timestamp 1621261055
transform 1 0 2304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_16
timestamp 1621261055
transform 1 0 2688 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_16
timestamp 1621261055
transform 1 0 2688 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_24
timestamp 1621261055
transform 1 0 3456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_24
timestamp 1621261055
transform 1 0 3456 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output599
timestamp 1621261055
transform 1 0 3072 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output595
timestamp 1621261055
transform 1 0 3072 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_248
timestamp 1621261055
transform 1 0 3648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_29
timestamp 1621261055
transform 1 0 3936 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_32
timestamp 1621261055
transform 1 0 4224 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_252
timestamp 1621261055
transform 1 0 4128 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output603
timestamp 1621261055
transform 1 0 4320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output600
timestamp 1621261055
transform 1 0 3840 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_258
timestamp 1621261055
transform 1 0 3840 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_41
timestamp 1621261055
transform 1 0 5088 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_37
timestamp 1621261055
transform 1 0 4704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_40
timestamp 1621261055
transform 1 0 4992 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output604
timestamp 1621261055
transform 1 0 5376 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output602
timestamp 1621261055
transform 1 0 4608 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _185_
timestamp 1621261055
transform 1 0 5280 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_46
timestamp 1621261055
transform 1 0 5568 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_52
timestamp 1621261055
transform 1 0 6144 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_48
timestamp 1621261055
transform 1 0 5760 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_54
timestamp 1621261055
transform 1 0 6336 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_54
timestamp 1621261055
transform 1 0 6336 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_62
timestamp 1621261055
transform 1 0 7104 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_64
timestamp 1621261055
transform 1 0 7296 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_56
timestamp 1621261055
transform 1 0 6528 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_232
timestamp 1621261055
transform 1 0 7488 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_95
timestamp 1621261055
transform 1 0 7488 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_248
timestamp 1621261055
transform 1 0 6432 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_72
timestamp 1621261055
transform 1 0 8064 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output581
timestamp 1621261055
transform 1 0 7680 0 -1 8658
box -38 -49 422 715
use AOI21X1  AOI21X1
timestamp 1624893035
transform 1 0 7680 0 1 7326
box 0 -48 1152 714
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_80
timestamp 1621261055
transform 1 0 8832 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_80
timestamp 1621261055
transform 1 0 8832 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_84
timestamp 1621261055
transform 1 0 9216 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_82
timestamp 1621261055
transform 1 0 9024 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_234
timestamp 1621261055
transform 1 0 9024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output583
timestamp 1621261055
transform 1 0 9216 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_259
timestamp 1621261055
transform 1 0 9120 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_88
timestamp 1621261055
transform 1 0 9600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_238
timestamp 1621261055
transform 1 0 9408 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output587
timestamp 1621261055
transform 1 0 9600 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_92
timestamp 1621261055
transform 1 0 9984 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_242
timestamp 1621261055
transform 1 0 10176 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output586
timestamp 1621261055
transform 1 0 9984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_100
timestamp 1621261055
transform 1 0 10752 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_96
timestamp 1621261055
transform 1 0 10368 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_240
timestamp 1621261055
transform 1 0 10560 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output589
timestamp 1621261055
transform 1 0 10368 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output588
timestamp 1621261055
transform 1 0 10752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_104
timestamp 1621261055
transform 1 0 11136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_244
timestamp 1621261055
transform 1 0 10944 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output590
timestamp 1621261055
transform 1 0 11136 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_108
timestamp 1621261055
transform 1 0 11520 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_108
timestamp 1621261055
transform 1 0 11520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_111
timestamp 1621261055
transform 1 0 11808 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output592
timestamp 1621261055
transform 1 0 11904 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_249
timestamp 1621261055
transform 1 0 11712 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_116
timestamp 1621261055
transform 1 0 12288 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output591
timestamp 1621261055
transform 1 0 12192 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_119
timestamp 1621261055
transform 1 0 12576 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output594
timestamp 1621261055
transform 1 0 12672 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_124
timestamp 1621261055
transform 1 0 13056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_127
timestamp 1621261055
transform 1 0 13344 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output593
timestamp 1621261055
transform 1 0 12960 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_132
timestamp 1621261055
transform 1 0 13824 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_246
timestamp 1621261055
transform 1 0 13536 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output597
timestamp 1621261055
transform 1 0 13440 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output596
timestamp 1621261055
transform 1 0 13728 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_135
timestamp 1621261055
transform 1 0 14112 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_139
timestamp 1621261055
transform 1 0 14496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_136
timestamp 1621261055
transform 1 0 14208 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_139
timestamp 1621261055
transform 1 0 14496 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_16
timestamp 1621261055
transform -1 0 14880 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_260
timestamp 1621261055
transform 1 0 14400 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _008_
timestamp 1621261055
transform -1 0 15168 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_147
timestamp 1621261055
transform 1 0 15264 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_150
timestamp 1621261055
transform 1 0 15552 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_146
timestamp 1621261055
transform 1 0 15168 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output549
timestamp 1621261055
transform 1 0 15648 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_159
timestamp 1621261055
transform 1 0 16416 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_155
timestamp 1621261055
transform 1 0 16032 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output560
timestamp 1621261055
transform 1 0 16032 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_167
timestamp 1621261055
transform 1 0 17184 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_166
timestamp 1621261055
transform 1 0 17088 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_163
timestamp 1621261055
transform 1 0 16800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output571
timestamp 1621261055
transform 1 0 16800 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_250
timestamp 1621261055
transform 1 0 16992 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_175
timestamp 1621261055
transform 1 0 17952 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_174
timestamp 1621261055
transform 1 0 17856 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _196_
timestamp 1621261055
transform 1 0 18144 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_8_188
timestamp 1621261055
transform 1 0 19200 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_180
timestamp 1621261055
transform 1 0 18432 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_182
timestamp 1621261055
transform 1 0 18624 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_194
timestamp 1621261055
transform 1 0 19776 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_192
timestamp 1621261055
transform 1 0 19584 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_7_190
timestamp 1621261055
transform 1 0 19392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_261
timestamp 1621261055
transform 1 0 19680 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_202
timestamp 1621261055
transform 1 0 20544 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_198
timestamp 1621261055
transform 1 0 20160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_142
timestamp 1621261055
transform 1 0 20544 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output485
timestamp 1621261055
transform 1 0 20736 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_210
timestamp 1621261055
transform 1 0 21312 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_208
timestamp 1621261055
transform 1 0 21120 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_216
timestamp 1621261055
transform 1 0 21888 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_218
timestamp 1621261055
transform 1 0 22080 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_221
timestamp 1621261055
transform 1 0 22368 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_251
timestamp 1621261055
transform 1 0 22272 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_226
timestamp 1621261055
transform 1 0 22848 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_229
timestamp 1621261055
transform 1 0 23136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_150
timestamp 1621261055
transform 1 0 23520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_242
timestamp 1621261055
transform 1 0 24384 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_234
timestamp 1621261055
transform 1 0 23616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_239
timestamp 1621261055
transform 1 0 24096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output493
timestamp 1621261055
transform 1 0 23712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output495
timestamp 1621261055
transform 1 0 24480 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_249
timestamp 1621261055
transform 1 0 25056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_246
timestamp 1621261055
transform 1 0 24768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_247
timestamp 1621261055
transform 1 0 24864 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output497
timestamp 1621261055
transform 1 0 25248 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_262
timestamp 1621261055
transform 1 0 24960 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_256
timestamp 1621261055
transform 1 0 25728 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_255
timestamp 1621261055
transform 1 0 25632 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output499
timestamp 1621261055
transform 1 0 26016 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _187_
timestamp 1621261055
transform 1 0 25440 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_264
timestamp 1621261055
transform 1 0 26496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_263
timestamp 1621261055
transform 1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output502
timestamp 1621261055
transform 1 0 26784 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_272
timestamp 1621261055
transform 1 0 27264 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_278
timestamp 1621261055
transform 1 0 27840 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_276
timestamp 1621261055
transform 1 0 27648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_271
timestamp 1621261055
transform 1 0 27168 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_252
timestamp 1621261055
transform 1 0 27552 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_280
timestamp 1621261055
transform 1 0 28032 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_285
timestamp 1621261055
transform 1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_156
timestamp 1621261055
transform 1 0 27936 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output507
timestamp 1621261055
transform 1 0 28128 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_292
timestamp 1621261055
transform 1 0 29184 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_288
timestamp 1621261055
transform 1 0 28800 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_296
timestamp 1621261055
transform 1 0 29568 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_7_291
timestamp 1621261055
transform 1 0 29088 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_289
timestamp 1621261055
transform 1 0 28896 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output510
timestamp 1621261055
transform 1 0 29184 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _103_
timestamp 1621261055
transform 1 0 29376 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_8_297
timestamp 1621261055
transform 1 0 29664 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_304
timestamp 1621261055
transform 1 0 30336 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_301
timestamp 1621261055
transform 1 0 30048 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_304
timestamp 1621261055
transform 1 0 30336 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_162
timestamp 1621261055
transform -1 0 29952 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output511
timestamp 1621261055
transform -1 0 30336 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_263
timestamp 1621261055
transform 1 0 30240 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_312
timestamp 1621261055
transform 1 0 31104 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_310
timestamp 1621261055
transform 1 0 30912 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_308
timestamp 1621261055
transform 1 0 30720 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output515
timestamp 1621261055
transform 1 0 31008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_320
timestamp 1621261055
transform 1 0 31872 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_323
timestamp 1621261055
transform 1 0 32160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_315
timestamp 1621261055
transform 1 0 31392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_328
timestamp 1621261055
transform 1 0 32640 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_331
timestamp 1621261055
transform 1 0 32928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_329
timestamp 1621261055
transform 1 0 32736 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_327
timestamp 1621261055
transform 1 0 32544 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_253
timestamp 1621261055
transform 1 0 32832 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_336
timestamp 1621261055
transform 1 0 33408 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_337
timestamp 1621261055
transform 1 0 33504 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_335
timestamp 1621261055
transform 1 0 33312 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output523
timestamp 1621261055
transform 1 0 33600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_344
timestamp 1621261055
transform 1 0 34176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_350
timestamp 1621261055
transform 1 0 34752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_342
timestamp 1621261055
transform 1 0 33984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output525
timestamp 1621261055
transform 1 0 34368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_359
timestamp 1621261055
transform 1 0 35616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_356
timestamp 1621261055
transform 1 0 35328 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_352
timestamp 1621261055
transform 1 0 34944 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_358
timestamp 1621261055
transform 1 0 35520 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output526
timestamp 1621261055
transform 1 0 35136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_264
timestamp 1621261055
transform 1 0 35520 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_367
timestamp 1621261055
transform 1 0 36384 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_366
timestamp 1621261055
transform 1 0 36288 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_179
timestamp 1621261055
transform -1 0 36672 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output530
timestamp 1621261055
transform 1 0 35904 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_375
timestamp 1621261055
transform 1 0 37152 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_374
timestamp 1621261055
transform 1 0 37056 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output532
timestamp 1621261055
transform -1 0 37056 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_383
timestamp 1621261055
transform 1 0 37920 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_386
timestamp 1621261055
transform 1 0 38208 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_7_384
timestamp 1621261055
transform 1 0 38016 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_382
timestamp 1621261055
transform 1 0 37824 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_254
timestamp 1621261055
transform 1 0 38112 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_393
timestamp 1621261055
transform 1 0 38880 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_387
timestamp 1621261055
transform 1 0 38304 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_394
timestamp 1621261055
transform 1 0 38976 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_241
timestamp 1621261055
transform -1 0 38592 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output536
timestamp 1621261055
transform 1 0 38592 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _207_
timestamp 1621261055
transform -1 0 38880 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_401
timestamp 1621261055
transform 1 0 39648 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_402
timestamp 1621261055
transform 1 0 39744 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output539
timestamp 1621261055
transform 1 0 39360 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_409
timestamp 1621261055
transform 1 0 40416 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_410
timestamp 1621261055
transform 1 0 40512 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_187
timestamp 1621261055
transform 1 0 40704 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output541
timestamp 1621261055
transform 1 0 40128 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_265
timestamp 1621261055
transform 1 0 40800 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_422
timestamp 1621261055
transform 1 0 41664 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_414
timestamp 1621261055
transform 1 0 40896 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_418
timestamp 1621261055
transform 1 0 41280 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output546
timestamp 1621261055
transform 1 0 41664 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output543
timestamp 1621261055
transform 1 0 40896 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_430
timestamp 1621261055
transform 1 0 42432 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_426
timestamp 1621261055
transform 1 0 42048 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_194
timestamp 1621261055
transform -1 0 42432 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output550
timestamp 1621261055
transform -1 0 42816 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_438
timestamp 1621261055
transform 1 0 43200 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_438
timestamp 1621261055
transform 1 0 43200 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_434
timestamp 1621261055
transform 1 0 42816 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_255
timestamp 1621261055
transform 1 0 43392 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_446
timestamp 1621261055
transform 1 0 43968 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_449
timestamp 1621261055
transform 1 0 44256 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_441
timestamp 1621261055
transform 1 0 43488 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output554
timestamp 1621261055
transform 1 0 43872 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_454
timestamp 1621261055
transform 1 0 44736 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_457
timestamp 1621261055
transform 1 0 45024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_202
timestamp 1621261055
transform 1 0 44448 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output556
timestamp 1621261055
transform 1 0 44640 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _197_
timestamp 1621261055
transform 1 0 44928 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_459
timestamp 1621261055
transform 1 0 45216 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_203
timestamp 1621261055
transform -1 0 45408 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_467
timestamp 1621261055
transform 1 0 45984 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_465
timestamp 1621261055
transform 1 0 45792 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_206
timestamp 1621261055
transform -1 0 46176 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output557
timestamp 1621261055
transform -1 0 45792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_469
timestamp 1621261055
transform 1 0 46176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_473
timestamp 1621261055
transform 1 0 46560 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output559
timestamp 1621261055
transform -1 0 46560 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_266
timestamp 1621261055
transform 1 0 46080 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_485
timestamp 1621261055
transform 1 0 47712 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_477
timestamp 1621261055
transform 1 0 46944 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_481
timestamp 1621261055
transform 1 0 47328 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_208
timestamp 1621261055
transform -1 0 47712 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output564
timestamp 1621261055
transform -1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output562
timestamp 1621261055
transform 1 0 46944 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_211
timestamp 1621261055
transform -1 0 48000 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_492
timestamp 1621261055
transform 1 0 48384 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_493
timestamp 1621261055
transform 1 0 48480 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_489
timestamp 1621261055
transform 1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_215
timestamp 1621261055
transform -1 0 48768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output566
timestamp 1621261055
transform -1 0 48384 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_500
timestamp 1621261055
transform 1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_496
timestamp 1621261055
transform 1 0 48768 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_213
timestamp 1621261055
transform -1 0 49152 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output568
timestamp 1621261055
transform -1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output567
timestamp 1621261055
transform -1 0 49536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_256
timestamp 1621261055
transform 1 0 48672 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_508
timestamp 1621261055
transform 1 0 49920 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_512
timestamp 1621261055
transform 1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_504
timestamp 1621261055
transform 1 0 49536 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_217
timestamp 1621261055
transform -1 0 49920 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output570
timestamp 1621261055
transform 1 0 49536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output569
timestamp 1621261055
transform -1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_520
timestamp 1621261055
transform 1 0 51072 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_516
timestamp 1621261055
transform 1 0 50688 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_516
timestamp 1621261055
transform 1 0 50688 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output473
timestamp 1621261055
transform 1 0 50880 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_524
timestamp 1621261055
transform 1 0 51456 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_522
timestamp 1621261055
transform 1 0 51264 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_530
timestamp 1621261055
transform 1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_522
timestamp 1621261055
transform 1 0 51264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_104
timestamp 1621261055
transform -1 0 51648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output450
timestamp 1621261055
transform -1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_267
timestamp 1621261055
transform 1 0 51360 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_537
timestamp 1621261055
transform 1 0 52704 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_532
timestamp 1621261055
transform 1 0 52224 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_538
timestamp 1621261055
transform 1 0 52800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_110
timestamp 1621261055
transform -1 0 53088 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output472
timestamp 1621261055
transform 1 0 52320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output452
timestamp 1621261055
transform 1 0 52416 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_108
timestamp 1621261055
transform -1 0 53184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_545
timestamp 1621261055
transform 1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_546
timestamp 1621261055
transform 1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output456
timestamp 1621261055
transform 1 0 53856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output454
timestamp 1621261055
transform -1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output453
timestamp 1621261055
transform -1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_553
timestamp 1621261055
transform 1 0 54240 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_551
timestamp 1621261055
transform 1 0 54048 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_257
timestamp 1621261055
transform 1 0 53952 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_566
timestamp 1621261055
transform 1 0 55488 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_561
timestamp 1621261055
transform 1 0 55008 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_565
timestamp 1621261055
transform 1 0 55392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_559
timestamp 1621261055
transform 1 0 54816 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input197
timestamp 1621261055
transform 1 0 55104 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input194
timestamp 1621261055
transform 1 0 55008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_574
timestamp 1621261055
transform 1 0 56256 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_573
timestamp 1621261055
transform 1 0 56160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input193
timestamp 1621261055
transform 1 0 55872 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input185
timestamp 1621261055
transform 1 0 55776 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_579
timestamp 1621261055
transform 1 0 56736 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_581
timestamp 1621261055
transform 1 0 56928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input188
timestamp 1621261055
transform 1 0 57120 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input186
timestamp 1621261055
transform 1 0 56544 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_268
timestamp 1621261055
transform 1 0 56640 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_587
timestamp 1621261055
transform 1 0 57504 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_589
timestamp 1621261055
transform 1 0 57696 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input187
timestamp 1621261055
transform 1 0 57312 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_15
timestamp 1621261055
transform -1 0 58848 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_17
timestamp 1621261055
transform -1 0 58848 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_595
timestamp 1621261055
transform 1 0 58272 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_18
timestamp 1621261055
transform 1 0 1152 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_4
timestamp 1621261055
transform 1 0 1536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_12
timestamp 1621261055
transform 1 0 2304 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_20
timestamp 1621261055
transform 1 0 3072 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _216_
timestamp 1621261055
transform 1 0 5376 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_29
timestamp 1621261055
transform 1 0 5184 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_28
timestamp 1621261055
transform 1 0 3840 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_36
timestamp 1621261055
transform 1 0 4608 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_40
timestamp 1621261055
transform 1 0 4992 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_47
timestamp 1621261055
transform 1 0 5664 0 1 8658
box -38 -49 806 715
use AOI22X1  AOI22X1
timestamp 1624893035
transform 1 0 7680 0 1 8658
box 0 -48 1440 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_269
timestamp 1621261055
transform 1 0 6432 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_39
timestamp 1621261055
transform 1 0 7488 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_56
timestamp 1621261055
transform 1 0 6528 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_64
timestamp 1621261055
transform 1 0 7296 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_83
timestamp 1621261055
transform 1 0 9120 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_91
timestamp 1621261055
transform 1 0 9888 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_99
timestamp 1621261055
transform 1 0 10656 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_107
timestamp 1621261055
transform 1 0 11424 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_270
timestamp 1621261055
transform 1 0 11712 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_9_109
timestamp 1621261055
transform 1 0 11616 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_111
timestamp 1621261055
transform 1 0 11808 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_119
timestamp 1621261055
transform 1 0 12576 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_127
timestamp 1621261055
transform 1 0 13344 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_135
timestamp 1621261055
transform 1 0 14112 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_143
timestamp 1621261055
transform 1 0 14880 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_151
timestamp 1621261055
transform 1 0 15648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_159
timestamp 1621261055
transform 1 0 16416 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_271
timestamp 1621261055
transform 1 0 16992 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_163
timestamp 1621261055
transform 1 0 16800 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_166
timestamp 1621261055
transform 1 0 17088 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_174
timestamp 1621261055
transform 1 0 17856 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_182
timestamp 1621261055
transform 1 0 18624 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_190
timestamp 1621261055
transform 1 0 19392 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_198
timestamp 1621261055
transform 1 0 20160 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_206
timestamp 1621261055
transform 1 0 20928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_214
timestamp 1621261055
transform 1 0 21696 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_272
timestamp 1621261055
transform 1 0 22272 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_218
timestamp 1621261055
transform 1 0 22080 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_221
timestamp 1621261055
transform 1 0 22368 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_229
timestamp 1621261055
transform 1 0 23136 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_237
timestamp 1621261055
transform 1 0 23904 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _138_
timestamp 1621261055
transform 1 0 25440 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_9_245
timestamp 1621261055
transform 1 0 24672 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_256
timestamp 1621261055
transform 1 0 25728 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_264
timestamp 1621261055
transform 1 0 26496 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_273
timestamp 1621261055
transform 1 0 27552 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_272
timestamp 1621261055
transform 1 0 27264 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_274
timestamp 1621261055
transform 1 0 27456 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_276
timestamp 1621261055
transform 1 0 27648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_284
timestamp 1621261055
transform 1 0 28416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_292
timestamp 1621261055
transform 1 0 29184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_300
timestamp 1621261055
transform 1 0 29952 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_308
timestamp 1621261055
transform 1 0 30720 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_316
timestamp 1621261055
transform 1 0 31488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_324
timestamp 1621261055
transform 1 0 32256 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_274
timestamp 1621261055
transform 1 0 32832 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_328
timestamp 1621261055
transform 1 0 32640 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_331
timestamp 1621261055
transform 1 0 32928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_339
timestamp 1621261055
transform 1 0 33696 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_347
timestamp 1621261055
transform 1 0 34464 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_355
timestamp 1621261055
transform 1 0 35232 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_363
timestamp 1621261055
transform 1 0 36000 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_371
timestamp 1621261055
transform 1 0 36768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_275
timestamp 1621261055
transform 1 0 38112 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_379
timestamp 1621261055
transform 1 0 37536 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_383
timestamp 1621261055
transform 1 0 37920 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_386
timestamp 1621261055
transform 1 0 38208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_394
timestamp 1621261055
transform 1 0 38976 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_402
timestamp 1621261055
transform 1 0 39744 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_410
timestamp 1621261055
transform 1 0 40512 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_418
timestamp 1621261055
transform 1 0 41280 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_426
timestamp 1621261055
transform 1 0 42048 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_276
timestamp 1621261055
transform 1 0 43392 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_434
timestamp 1621261055
transform 1 0 42816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_438
timestamp 1621261055
transform 1 0 43200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_441
timestamp 1621261055
transform 1 0 43488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_449
timestamp 1621261055
transform 1 0 44256 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_457
timestamp 1621261055
transform 1 0 45024 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_465
timestamp 1621261055
transform 1 0 45792 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_473
timestamp 1621261055
transform 1 0 46560 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_481
timestamp 1621261055
transform 1 0 47328 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_277
timestamp 1621261055
transform 1 0 48672 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_489
timestamp 1621261055
transform 1 0 48096 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_493
timestamp 1621261055
transform 1 0 48480 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_496
timestamp 1621261055
transform 1 0 48768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_504
timestamp 1621261055
transform 1 0 49536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_512
timestamp 1621261055
transform 1 0 50304 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_127
timestamp 1621261055
transform -1 0 53184 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_520
timestamp 1621261055
transform 1 0 51072 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_528
timestamp 1621261055
transform 1 0 51840 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_536
timestamp 1621261055
transform 1 0 52608 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output469
timestamp 1621261055
transform -1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_546
timestamp 1621261055
transform 1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_551
timestamp 1621261055
transform 1 0 54048 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_113
timestamp 1621261055
transform -1 0 54432 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_278
timestamp 1621261055
transform 1 0 53952 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_559
timestamp 1621261055
transform 1 0 54816 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output457
timestamp 1621261055
transform -1 0 54816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_115
timestamp 1621261055
transform -1 0 55200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output459
timestamp 1621261055
transform -1 0 55584 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_116
timestamp 1621261055
transform -1 0 55776 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input190
timestamp 1621261055
transform 1 0 57216 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input195
timestamp 1621261055
transform 1 0 56448 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_569
timestamp 1621261055
transform 1 0 55776 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_573
timestamp 1621261055
transform 1 0 56160 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_575
timestamp 1621261055
transform 1 0 56352 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_580
timestamp 1621261055
transform 1 0 56832 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_588
timestamp 1621261055
transform 1 0 57600 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_19
timestamp 1621261055
transform -1 0 58848 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_596
timestamp 1621261055
transform 1 0 58368 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_20
timestamp 1621261055
transform 1 0 1152 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_10_4
timestamp 1621261055
transform 1 0 1536 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_12
timestamp 1621261055
transform 1 0 2304 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_20
timestamp 1621261055
transform 1 0 3072 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_279
timestamp 1621261055
transform 1 0 3840 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_29
timestamp 1621261055
transform 1 0 3936 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_37
timestamp 1621261055
transform 1 0 4704 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_45
timestamp 1621261055
transform 1 0 5472 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_53
timestamp 1621261055
transform 1 0 6240 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_61
timestamp 1621261055
transform 1 0 7008 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_69
timestamp 1621261055
transform 1 0 7776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_77
timestamp 1621261055
transform 1 0 8544 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_81
timestamp 1621261055
transform 1 0 8928 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_280
timestamp 1621261055
transform 1 0 9120 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_84
timestamp 1621261055
transform 1 0 9216 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_92
timestamp 1621261055
transform 1 0 9984 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_100
timestamp 1621261055
transform 1 0 10752 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_108
timestamp 1621261055
transform 1 0 11520 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_116
timestamp 1621261055
transform 1 0 12288 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_124
timestamp 1621261055
transform 1 0 13056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_132
timestamp 1621261055
transform 1 0 13824 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_281
timestamp 1621261055
transform 1 0 14400 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_136
timestamp 1621261055
transform 1 0 14208 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_139
timestamp 1621261055
transform 1 0 14496 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_147
timestamp 1621261055
transform 1 0 15264 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_155
timestamp 1621261055
transform 1 0 16032 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_163
timestamp 1621261055
transform 1 0 16800 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_171
timestamp 1621261055
transform 1 0 17568 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_179
timestamp 1621261055
transform 1 0 18336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_187
timestamp 1621261055
transform 1 0 19104 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_282
timestamp 1621261055
transform 1 0 19680 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_191
timestamp 1621261055
transform 1 0 19488 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_194
timestamp 1621261055
transform 1 0 19776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_202
timestamp 1621261055
transform 1 0 20544 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_210
timestamp 1621261055
transform 1 0 21312 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_218
timestamp 1621261055
transform 1 0 22080 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_226
timestamp 1621261055
transform 1 0 22848 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_234
timestamp 1621261055
transform 1 0 23616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_242
timestamp 1621261055
transform 1 0 24384 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _192_
timestamp 1621261055
transform 1 0 25632 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_283
timestamp 1621261055
transform 1 0 24960 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_246
timestamp 1621261055
transform 1 0 24768 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_10_249
timestamp 1621261055
transform 1 0 25056 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_253
timestamp 1621261055
transform 1 0 25440 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_258
timestamp 1621261055
transform 1 0 25920 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_266
timestamp 1621261055
transform 1 0 26688 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_274
timestamp 1621261055
transform 1 0 27456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_282
timestamp 1621261055
transform 1 0 28224 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_290
timestamp 1621261055
transform 1 0 28992 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _122_
timestamp 1621261055
transform 1 0 32160 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_284
timestamp 1621261055
transform 1 0 30240 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_298
timestamp 1621261055
transform 1 0 29760 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_302
timestamp 1621261055
transform 1 0 30144 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_304
timestamp 1621261055
transform 1 0 30336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_312
timestamp 1621261055
transform 1 0 31104 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_320
timestamp 1621261055
transform 1 0 31872 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_322
timestamp 1621261055
transform 1 0 32064 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_326
timestamp 1621261055
transform 1 0 32448 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_334
timestamp 1621261055
transform 1 0 33216 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_342
timestamp 1621261055
transform 1 0 33984 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_350
timestamp 1621261055
transform 1 0 34752 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_285
timestamp 1621261055
transform 1 0 35520 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_359
timestamp 1621261055
transform 1 0 35616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_367
timestamp 1621261055
transform 1 0 36384 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_375
timestamp 1621261055
transform 1 0 37152 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_383
timestamp 1621261055
transform 1 0 37920 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_391
timestamp 1621261055
transform 1 0 38688 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_399
timestamp 1621261055
transform 1 0 39456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_286
timestamp 1621261055
transform 1 0 40800 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_407
timestamp 1621261055
transform 1 0 40224 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_411
timestamp 1621261055
transform 1 0 40608 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_414
timestamp 1621261055
transform 1 0 40896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_422
timestamp 1621261055
transform 1 0 41664 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_430
timestamp 1621261055
transform 1 0 42432 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_438
timestamp 1621261055
transform 1 0 43200 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_446
timestamp 1621261055
transform 1 0 43968 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_454
timestamp 1621261055
transform 1 0 44736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_287
timestamp 1621261055
transform 1 0 46080 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_462
timestamp 1621261055
transform 1 0 45504 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_466
timestamp 1621261055
transform 1 0 45888 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_469
timestamp 1621261055
transform 1 0 46176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_477
timestamp 1621261055
transform 1 0 46944 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_485
timestamp 1621261055
transform 1 0 47712 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_493
timestamp 1621261055
transform 1 0 48480 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_501
timestamp 1621261055
transform 1 0 49248 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_509
timestamp 1621261055
transform 1 0 50016 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_288
timestamp 1621261055
transform 1 0 51360 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_517
timestamp 1621261055
transform 1 0 50784 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_521
timestamp 1621261055
transform 1 0 51168 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_524
timestamp 1621261055
transform 1 0 51456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_532
timestamp 1621261055
transform 1 0 52224 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_540
timestamp 1621261055
transform 1 0 52992 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output458
timestamp 1621261055
transform 1 0 54240 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output460
timestamp 1621261055
transform 1 0 55008 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_548
timestamp 1621261055
transform 1 0 53760 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_552
timestamp 1621261055
transform 1 0 54144 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_557
timestamp 1621261055
transform 1 0 54624 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_565
timestamp 1621261055
transform 1 0 55392 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_289
timestamp 1621261055
transform 1 0 56640 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input191
timestamp 1621261055
transform 1 0 57600 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output461
timestamp 1621261055
transform 1 0 55776 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_10_573
timestamp 1621261055
transform 1 0 56160 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_577
timestamp 1621261055
transform 1 0 56544 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_579
timestamp 1621261055
transform 1 0 56736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_10_587
timestamp 1621261055
transform 1 0 57504 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_592
timestamp 1621261055
transform 1 0 57984 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_21
timestamp 1621261055
transform -1 0 58848 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_596
timestamp 1621261055
transform 1 0 58368 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_22
timestamp 1621261055
transform 1 0 1152 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_4
timestamp 1621261055
transform 1 0 1536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_12
timestamp 1621261055
transform 1 0 2304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_20
timestamp 1621261055
transform 1 0 3072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_28
timestamp 1621261055
transform 1 0 3840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_36
timestamp 1621261055
transform 1 0 4608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_44
timestamp 1621261055
transform 1 0 5376 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_52
timestamp 1621261055
transform 1 0 6144 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_54
timestamp 1621261055
transform 1 0 6336 0 1 9990
box -38 -49 134 715
use BUFX2  BUFX2
timestamp 1624893035
transform 1 0 7680 0 1 9990
box 0 -48 864 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_290
timestamp 1621261055
transform 1 0 6432 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_43
timestamp 1621261055
transform 1 0 7488 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_56
timestamp 1621261055
transform 1 0 6528 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_64
timestamp 1621261055
transform 1 0 7296 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_77
timestamp 1621261055
transform 1 0 8544 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_85
timestamp 1621261055
transform 1 0 9312 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_93
timestamp 1621261055
transform 1 0 10080 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_101
timestamp 1621261055
transform 1 0 10848 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_291
timestamp 1621261055
transform 1 0 11712 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_11_109
timestamp 1621261055
transform 1 0 11616 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_111
timestamp 1621261055
transform 1 0 11808 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_119
timestamp 1621261055
transform 1 0 12576 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_127
timestamp 1621261055
transform 1 0 13344 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_135
timestamp 1621261055
transform 1 0 14112 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_143
timestamp 1621261055
transform 1 0 14880 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_151
timestamp 1621261055
transform 1 0 15648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_159
timestamp 1621261055
transform 1 0 16416 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_292
timestamp 1621261055
transform 1 0 16992 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_163
timestamp 1621261055
transform 1 0 16800 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_166
timestamp 1621261055
transform 1 0 17088 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_174
timestamp 1621261055
transform 1 0 17856 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_182
timestamp 1621261055
transform 1 0 18624 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_190
timestamp 1621261055
transform 1 0 19392 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_198
timestamp 1621261055
transform 1 0 20160 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_206
timestamp 1621261055
transform 1 0 20928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_214
timestamp 1621261055
transform 1 0 21696 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_293
timestamp 1621261055
transform 1 0 22272 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_218
timestamp 1621261055
transform 1 0 22080 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_221
timestamp 1621261055
transform 1 0 22368 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_229
timestamp 1621261055
transform 1 0 23136 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_237
timestamp 1621261055
transform 1 0 23904 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_245
timestamp 1621261055
transform 1 0 24672 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_253
timestamp 1621261055
transform 1 0 25440 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_261
timestamp 1621261055
transform 1 0 26208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_269
timestamp 1621261055
transform 1 0 26976 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _062_
timestamp 1621261055
transform 1 0 28224 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _080_
timestamp 1621261055
transform 1 0 28992 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_294
timestamp 1621261055
transform 1 0 27552 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_273
timestamp 1621261055
transform 1 0 27360 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_276
timestamp 1621261055
transform 1 0 27648 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_280
timestamp 1621261055
transform 1 0 28032 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_285
timestamp 1621261055
transform 1 0 28512 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_289
timestamp 1621261055
transform 1 0 28896 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_293
timestamp 1621261055
transform 1 0 29280 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_301
timestamp 1621261055
transform 1 0 30048 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_309
timestamp 1621261055
transform 1 0 30816 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_317
timestamp 1621261055
transform 1 0 31584 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_295
timestamp 1621261055
transform 1 0 32832 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_325
timestamp 1621261055
transform 1 0 32352 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_329
timestamp 1621261055
transform 1 0 32736 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_331
timestamp 1621261055
transform 1 0 32928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_339
timestamp 1621261055
transform 1 0 33696 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_347
timestamp 1621261055
transform 1 0 34464 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_355
timestamp 1621261055
transform 1 0 35232 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_363
timestamp 1621261055
transform 1 0 36000 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_371
timestamp 1621261055
transform 1 0 36768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_296
timestamp 1621261055
transform 1 0 38112 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_379
timestamp 1621261055
transform 1 0 37536 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_383
timestamp 1621261055
transform 1 0 37920 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_386
timestamp 1621261055
transform 1 0 38208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_394
timestamp 1621261055
transform 1 0 38976 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_402
timestamp 1621261055
transform 1 0 39744 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _179_
timestamp 1621261055
transform 1 0 41280 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_11_410
timestamp 1621261055
transform 1 0 40512 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_421
timestamp 1621261055
transform 1 0 41568 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_429
timestamp 1621261055
transform 1 0 42336 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_297
timestamp 1621261055
transform 1 0 43392 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_437
timestamp 1621261055
transform 1 0 43104 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_439
timestamp 1621261055
transform 1 0 43296 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_441
timestamp 1621261055
transform 1 0 43488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_449
timestamp 1621261055
transform 1 0 44256 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_457
timestamp 1621261055
transform 1 0 45024 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_465
timestamp 1621261055
transform 1 0 45792 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_473
timestamp 1621261055
transform 1 0 46560 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_481
timestamp 1621261055
transform 1 0 47328 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_298
timestamp 1621261055
transform 1 0 48672 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_489
timestamp 1621261055
transform 1 0 48096 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_493
timestamp 1621261055
transform 1 0 48480 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_496
timestamp 1621261055
transform 1 0 48768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_504
timestamp 1621261055
transform 1 0 49536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_512
timestamp 1621261055
transform 1 0 50304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_520
timestamp 1621261055
transform 1 0 51072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_528
timestamp 1621261055
transform 1 0 51840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_536
timestamp 1621261055
transform 1 0 52608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_299
timestamp 1621261055
transform 1 0 53952 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output471
timestamp 1621261055
transform 1 0 54912 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_117
timestamp 1621261055
transform -1 0 55680 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_544
timestamp 1621261055
transform 1 0 53376 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_548
timestamp 1621261055
transform 1 0 53760 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_551
timestamp 1621261055
transform 1 0 54048 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_11_559
timestamp 1621261055
transform 1 0 54816 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_564
timestamp 1621261055
transform 1 0 55296 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output462
timestamp 1621261055
transform -1 0 56064 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output463
timestamp 1621261055
transform -1 0 56832 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output464
timestamp 1621261055
transform -1 0 57600 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_119
timestamp 1621261055
transform -1 0 56448 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_120
timestamp 1621261055
transform -1 0 57024 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_121
timestamp 1621261055
transform -1 0 57216 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_572
timestamp 1621261055
transform 1 0 56064 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_588
timestamp 1621261055
transform 1 0 57600 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_23
timestamp 1621261055
transform -1 0 58848 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_596
timestamp 1621261055
transform 1 0 58368 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_24
timestamp 1621261055
transform 1 0 1152 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_4
timestamp 1621261055
transform 1 0 1536 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_12
timestamp 1621261055
transform 1 0 2304 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_20
timestamp 1621261055
transform 1 0 3072 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_300
timestamp 1621261055
transform 1 0 3840 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_29
timestamp 1621261055
transform 1 0 3936 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_37
timestamp 1621261055
transform 1 0 4704 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_45
timestamp 1621261055
transform 1 0 5472 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_53
timestamp 1621261055
transform 1 0 6240 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_61
timestamp 1621261055
transform 1 0 7008 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_69
timestamp 1621261055
transform 1 0 7776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_77
timestamp 1621261055
transform 1 0 8544 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_81
timestamp 1621261055
transform 1 0 8928 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_301
timestamp 1621261055
transform 1 0 9120 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_84
timestamp 1621261055
transform 1 0 9216 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_92
timestamp 1621261055
transform 1 0 9984 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_100
timestamp 1621261055
transform 1 0 10752 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_108
timestamp 1621261055
transform 1 0 11520 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _114_
timestamp 1621261055
transform 1 0 11904 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_115
timestamp 1621261055
transform 1 0 12192 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_123
timestamp 1621261055
transform 1 0 12960 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_131
timestamp 1621261055
transform 1 0 13728 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_135
timestamp 1621261055
transform 1 0 14112 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_302
timestamp 1621261055
transform 1 0 14400 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_12_137
timestamp 1621261055
transform 1 0 14304 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_139
timestamp 1621261055
transform 1 0 14496 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_147
timestamp 1621261055
transform 1 0 15264 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_155
timestamp 1621261055
transform 1 0 16032 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_163
timestamp 1621261055
transform 1 0 16800 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_171
timestamp 1621261055
transform 1 0 17568 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_179
timestamp 1621261055
transform 1 0 18336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_187
timestamp 1621261055
transform 1 0 19104 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_303
timestamp 1621261055
transform 1 0 19680 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_191
timestamp 1621261055
transform 1 0 19488 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_194
timestamp 1621261055
transform 1 0 19776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_202
timestamp 1621261055
transform 1 0 20544 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_210
timestamp 1621261055
transform 1 0 21312 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_218
timestamp 1621261055
transform 1 0 22080 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_226
timestamp 1621261055
transform 1 0 22848 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_234
timestamp 1621261055
transform 1 0 23616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_242
timestamp 1621261055
transform 1 0 24384 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_304
timestamp 1621261055
transform 1 0 24960 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_246
timestamp 1621261055
transform 1 0 24768 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_249
timestamp 1621261055
transform 1 0 25056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_257
timestamp 1621261055
transform 1 0 25824 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_265
timestamp 1621261055
transform 1 0 26592 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_273
timestamp 1621261055
transform 1 0 27360 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_281
timestamp 1621261055
transform 1 0 28128 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_289
timestamp 1621261055
transform 1 0 28896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_297
timestamp 1621261055
transform 1 0 29664 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_305
timestamp 1621261055
transform 1 0 30240 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_301
timestamp 1621261055
transform 1 0 30048 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_304
timestamp 1621261055
transform 1 0 30336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_312
timestamp 1621261055
transform 1 0 31104 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_320
timestamp 1621261055
transform 1 0 31872 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_328
timestamp 1621261055
transform 1 0 32640 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_336
timestamp 1621261055
transform 1 0 33408 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_344
timestamp 1621261055
transform 1 0 34176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_306
timestamp 1621261055
transform 1 0 35520 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_352
timestamp 1621261055
transform 1 0 34944 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_356
timestamp 1621261055
transform 1 0 35328 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_359
timestamp 1621261055
transform 1 0 35616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_367
timestamp 1621261055
transform 1 0 36384 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_375
timestamp 1621261055
transform 1 0 37152 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_383
timestamp 1621261055
transform 1 0 37920 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_391
timestamp 1621261055
transform 1 0 38688 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_399
timestamp 1621261055
transform 1 0 39456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_307
timestamp 1621261055
transform 1 0 40800 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_407
timestamp 1621261055
transform 1 0 40224 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_411
timestamp 1621261055
transform 1 0 40608 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_414
timestamp 1621261055
transform 1 0 40896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_422
timestamp 1621261055
transform 1 0 41664 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_430
timestamp 1621261055
transform 1 0 42432 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_438
timestamp 1621261055
transform 1 0 43200 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_446
timestamp 1621261055
transform 1 0 43968 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_454
timestamp 1621261055
transform 1 0 44736 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_308
timestamp 1621261055
transform 1 0 46080 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_462
timestamp 1621261055
transform 1 0 45504 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_466
timestamp 1621261055
transform 1 0 45888 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_469
timestamp 1621261055
transform 1 0 46176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_477
timestamp 1621261055
transform 1 0 46944 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_485
timestamp 1621261055
transform 1 0 47712 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_493
timestamp 1621261055
transform 1 0 48480 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_501
timestamp 1621261055
transform 1 0 49248 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_509
timestamp 1621261055
transform 1 0 50016 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_309
timestamp 1621261055
transform 1 0 51360 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_517
timestamp 1621261055
transform 1 0 50784 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_521
timestamp 1621261055
transform 1 0 51168 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_524
timestamp 1621261055
transform 1 0 51456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_532
timestamp 1621261055
transform 1 0 52224 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_540
timestamp 1621261055
transform 1 0 52992 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_548
timestamp 1621261055
transform 1 0 53760 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_556
timestamp 1621261055
transform 1 0 54528 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_564
timestamp 1621261055
transform 1 0 55296 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_310
timestamp 1621261055
transform 1 0 56640 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output465
timestamp 1621261055
transform -1 0 57504 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output470
timestamp 1621261055
transform -1 0 56256 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_122
timestamp 1621261055
transform -1 0 57120 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_129
timestamp 1621261055
transform -1 0 55872 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_130
timestamp 1621261055
transform -1 0 56448 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_576
timestamp 1621261055
transform 1 0 56448 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_579
timestamp 1621261055
transform 1 0 56736 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_587
timestamp 1621261055
transform 1 0 57504 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_25
timestamp 1621261055
transform -1 0 58848 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_595
timestamp 1621261055
transform 1 0 58272 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _035_
timestamp 1621261055
transform 1 0 1536 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_26
timestamp 1621261055
transform 1 0 1152 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_35
timestamp 1621261055
transform 1 0 1824 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_9
timestamp 1621261055
transform 1 0 2016 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_17
timestamp 1621261055
transform 1 0 2784 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_25
timestamp 1621261055
transform 1 0 3552 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _209_
timestamp 1621261055
transform 1 0 4992 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_13_33
timestamp 1621261055
transform 1 0 4320 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_37
timestamp 1621261055
transform 1 0 4704 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_39
timestamp 1621261055
transform 1 0 4896 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_43
timestamp 1621261055
transform 1 0 5280 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_51
timestamp 1621261055
transform 1 0 6048 0 1 11322
box -38 -49 422 715
use BUFX4  BUFX4
timestamp 1624893035
transform 1 0 7680 0 1 11322
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_311
timestamp 1621261055
transform 1 0 6432 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_47
timestamp 1621261055
transform 1 0 7488 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_56
timestamp 1621261055
transform 1 0 6528 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_64
timestamp 1621261055
transform 1 0 7296 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_80
timestamp 1621261055
transform 1 0 8832 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _051_
timestamp 1621261055
transform 1 0 9312 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_63
timestamp 1621261055
transform 1 0 9120 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_82
timestamp 1621261055
transform 1 0 9024 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_88
timestamp 1621261055
transform 1 0 9600 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_96
timestamp 1621261055
transform 1 0 10368 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_104
timestamp 1621261055
transform 1 0 11136 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_108
timestamp 1621261055
transform 1 0 11520 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_312
timestamp 1621261055
transform 1 0 11712 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_111
timestamp 1621261055
transform 1 0 11808 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_119
timestamp 1621261055
transform 1 0 12576 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_127
timestamp 1621261055
transform 1 0 13344 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_135
timestamp 1621261055
transform 1 0 14112 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_143
timestamp 1621261055
transform 1 0 14880 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_151
timestamp 1621261055
transform 1 0 15648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_159
timestamp 1621261055
transform 1 0 16416 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_313
timestamp 1621261055
transform 1 0 16992 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_163
timestamp 1621261055
transform 1 0 16800 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_166
timestamp 1621261055
transform 1 0 17088 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_174
timestamp 1621261055
transform 1 0 17856 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_182
timestamp 1621261055
transform 1 0 18624 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_190
timestamp 1621261055
transform 1 0 19392 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_198
timestamp 1621261055
transform 1 0 20160 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_206
timestamp 1621261055
transform 1 0 20928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_214
timestamp 1621261055
transform 1 0 21696 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_314
timestamp 1621261055
transform 1 0 22272 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_218
timestamp 1621261055
transform 1 0 22080 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_221
timestamp 1621261055
transform 1 0 22368 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_229
timestamp 1621261055
transform 1 0 23136 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_237
timestamp 1621261055
transform 1 0 23904 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_245
timestamp 1621261055
transform 1 0 24672 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_253
timestamp 1621261055
transform 1 0 25440 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_261
timestamp 1621261055
transform 1 0 26208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_269
timestamp 1621261055
transform 1 0 26976 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_315
timestamp 1621261055
transform 1 0 27552 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_273
timestamp 1621261055
transform 1 0 27360 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_276
timestamp 1621261055
transform 1 0 27648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_284
timestamp 1621261055
transform 1 0 28416 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_292
timestamp 1621261055
transform 1 0 29184 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_300
timestamp 1621261055
transform 1 0 29952 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_308
timestamp 1621261055
transform 1 0 30720 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_316
timestamp 1621261055
transform 1 0 31488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_324
timestamp 1621261055
transform 1 0 32256 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_316
timestamp 1621261055
transform 1 0 32832 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_328
timestamp 1621261055
transform 1 0 32640 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_331
timestamp 1621261055
transform 1 0 32928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_339
timestamp 1621261055
transform 1 0 33696 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_347
timestamp 1621261055
transform 1 0 34464 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _120_
timestamp 1621261055
transform 1 0 37440 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_13_355
timestamp 1621261055
transform 1 0 35232 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_363
timestamp 1621261055
transform 1 0 36000 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_371
timestamp 1621261055
transform 1 0 36768 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_375
timestamp 1621261055
transform 1 0 37152 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_377
timestamp 1621261055
transform 1 0 37344 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_317
timestamp 1621261055
transform 1 0 38112 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_381
timestamp 1621261055
transform 1 0 37728 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_386
timestamp 1621261055
transform 1 0 38208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_394
timestamp 1621261055
transform 1 0 38976 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_402
timestamp 1621261055
transform 1 0 39744 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_410
timestamp 1621261055
transform 1 0 40512 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_418
timestamp 1621261055
transform 1 0 41280 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_426
timestamp 1621261055
transform 1 0 42048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_318
timestamp 1621261055
transform 1 0 43392 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_434
timestamp 1621261055
transform 1 0 42816 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_438
timestamp 1621261055
transform 1 0 43200 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_441
timestamp 1621261055
transform 1 0 43488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_449
timestamp 1621261055
transform 1 0 44256 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_457
timestamp 1621261055
transform 1 0 45024 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_465
timestamp 1621261055
transform 1 0 45792 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_473
timestamp 1621261055
transform 1 0 46560 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_481
timestamp 1621261055
transform 1 0 47328 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_319
timestamp 1621261055
transform 1 0 48672 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_489
timestamp 1621261055
transform 1 0 48096 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_493
timestamp 1621261055
transform 1 0 48480 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_496
timestamp 1621261055
transform 1 0 48768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_504
timestamp 1621261055
transform 1 0 49536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_512
timestamp 1621261055
transform 1 0 50304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_520
timestamp 1621261055
transform 1 0 51072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_528
timestamp 1621261055
transform 1 0 51840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_536
timestamp 1621261055
transform 1 0 52608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _071_
timestamp 1621261055
transform 1 0 54432 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_320
timestamp 1621261055
transform 1 0 53952 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_544
timestamp 1621261055
transform 1 0 53376 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_548
timestamp 1621261055
transform 1 0 53760 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_551
timestamp 1621261055
transform 1 0 54048 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_558
timestamp 1621261055
transform 1 0 54720 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_566
timestamp 1621261055
transform 1 0 55488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output467
timestamp 1621261055
transform -1 0 57504 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output474
timestamp 1621261055
transform 1 0 56352 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_125
timestamp 1621261055
transform -1 0 57120 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_574
timestamp 1621261055
transform 1 0 56256 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_579
timestamp 1621261055
transform 1 0 56736 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_587
timestamp 1621261055
transform 1 0 57504 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_27
timestamp 1621261055
transform -1 0 58848 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_595
timestamp 1621261055
transform 1 0 58272 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_28
timestamp 1621261055
transform 1 0 1152 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_14_4
timestamp 1621261055
transform 1 0 1536 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_12
timestamp 1621261055
transform 1 0 2304 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_20
timestamp 1621261055
transform 1 0 3072 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _064_
timestamp 1621261055
transform 1 0 4800 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_321
timestamp 1621261055
transform 1 0 3840 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_29
timestamp 1621261055
transform 1 0 3936 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_14_37
timestamp 1621261055
transform 1 0 4704 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_41
timestamp 1621261055
transform 1 0 5088 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_49
timestamp 1621261055
transform 1 0 5856 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_57
timestamp 1621261055
transform 1 0 6624 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_65
timestamp 1621261055
transform 1 0 7392 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_73
timestamp 1621261055
transform 1 0 8160 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_81
timestamp 1621261055
transform 1 0 8928 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_322
timestamp 1621261055
transform 1 0 9120 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_84
timestamp 1621261055
transform 1 0 9216 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_92
timestamp 1621261055
transform 1 0 9984 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_100
timestamp 1621261055
transform 1 0 10752 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_108
timestamp 1621261055
transform 1 0 11520 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_116
timestamp 1621261055
transform 1 0 12288 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_124
timestamp 1621261055
transform 1 0 13056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_132
timestamp 1621261055
transform 1 0 13824 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _132_
timestamp 1621261055
transform 1 0 14976 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_323
timestamp 1621261055
transform 1 0 14400 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_136
timestamp 1621261055
transform 1 0 14208 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_139
timestamp 1621261055
transform 1 0 14496 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_14_143
timestamp 1621261055
transform 1 0 14880 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_147
timestamp 1621261055
transform 1 0 15264 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_155
timestamp 1621261055
transform 1 0 16032 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _077_
timestamp 1621261055
transform 1 0 18528 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_14_163
timestamp 1621261055
transform 1 0 16800 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_171
timestamp 1621261055
transform 1 0 17568 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_179
timestamp 1621261055
transform 1 0 18336 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_184
timestamp 1621261055
transform 1 0 18816 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_324
timestamp 1621261055
transform 1 0 19680 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_14_192
timestamp 1621261055
transform 1 0 19584 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_194
timestamp 1621261055
transform 1 0 19776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_202
timestamp 1621261055
transform 1 0 20544 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_210
timestamp 1621261055
transform 1 0 21312 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_218
timestamp 1621261055
transform 1 0 22080 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_226
timestamp 1621261055
transform 1 0 22848 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_234
timestamp 1621261055
transform 1 0 23616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_242
timestamp 1621261055
transform 1 0 24384 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_325
timestamp 1621261055
transform 1 0 24960 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_246
timestamp 1621261055
transform 1 0 24768 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_249
timestamp 1621261055
transform 1 0 25056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_257
timestamp 1621261055
transform 1 0 25824 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_265
timestamp 1621261055
transform 1 0 26592 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _105_
timestamp 1621261055
transform 1 0 29376 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_14_273
timestamp 1621261055
transform 1 0 27360 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_281
timestamp 1621261055
transform 1 0 28128 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_289
timestamp 1621261055
transform 1 0 28896 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_14_293
timestamp 1621261055
transform 1 0 29280 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_297
timestamp 1621261055
transform 1 0 29664 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _012_
timestamp 1621261055
transform -1 0 31392 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_326
timestamp 1621261055
transform 1 0 30240 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_22
timestamp 1621261055
transform -1 0 31104 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_301
timestamp 1621261055
transform 1 0 30048 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_304
timestamp 1621261055
transform 1 0 30336 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_308
timestamp 1621261055
transform 1 0 30720 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_315
timestamp 1621261055
transform 1 0 31392 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_323
timestamp 1621261055
transform 1 0 32160 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_331
timestamp 1621261055
transform 1 0 32928 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_339
timestamp 1621261055
transform 1 0 33696 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_347
timestamp 1621261055
transform 1 0 34464 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_327
timestamp 1621261055
transform 1 0 35520 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_355
timestamp 1621261055
transform 1 0 35232 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_14_357
timestamp 1621261055
transform 1 0 35424 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_359
timestamp 1621261055
transform 1 0 35616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_367
timestamp 1621261055
transform 1 0 36384 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_375
timestamp 1621261055
transform 1 0 37152 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_383
timestamp 1621261055
transform 1 0 37920 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_391
timestamp 1621261055
transform 1 0 38688 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_399
timestamp 1621261055
transform 1 0 39456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_328
timestamp 1621261055
transform 1 0 40800 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_407
timestamp 1621261055
transform 1 0 40224 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_411
timestamp 1621261055
transform 1 0 40608 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_414
timestamp 1621261055
transform 1 0 40896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_422
timestamp 1621261055
transform 1 0 41664 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_430
timestamp 1621261055
transform 1 0 42432 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_438
timestamp 1621261055
transform 1 0 43200 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_446
timestamp 1621261055
transform 1 0 43968 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_454
timestamp 1621261055
transform 1 0 44736 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_329
timestamp 1621261055
transform 1 0 46080 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_462
timestamp 1621261055
transform 1 0 45504 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_466
timestamp 1621261055
transform 1 0 45888 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_469
timestamp 1621261055
transform 1 0 46176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_477
timestamp 1621261055
transform 1 0 46944 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_485
timestamp 1621261055
transform 1 0 47712 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_493
timestamp 1621261055
transform 1 0 48480 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_501
timestamp 1621261055
transform 1 0 49248 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_509
timestamp 1621261055
transform 1 0 50016 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_330
timestamp 1621261055
transform 1 0 51360 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_14_517
timestamp 1621261055
transform 1 0 50784 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_521
timestamp 1621261055
transform 1 0 51168 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_524
timestamp 1621261055
transform 1 0 51456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_532
timestamp 1621261055
transform 1 0 52224 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_540
timestamp 1621261055
transform 1 0 52992 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_548
timestamp 1621261055
transform 1 0 53760 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_556
timestamp 1621261055
transform 1 0 54528 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_564
timestamp 1621261055
transform 1 0 55296 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_331
timestamp 1621261055
transform 1 0 56640 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output468
timestamp 1621261055
transform 1 0 57504 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_14_572
timestamp 1621261055
transform 1 0 56064 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_576
timestamp 1621261055
transform 1 0 56448 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_579
timestamp 1621261055
transform 1 0 56736 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_591
timestamp 1621261055
transform 1 0 57888 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_29
timestamp 1621261055
transform -1 0 58848 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_595
timestamp 1621261055
transform 1 0 58272 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_30
timestamp 1621261055
transform 1 0 1152 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_32
timestamp 1621261055
transform 1 0 1152 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_4
timestamp 1621261055
transform 1 0 1536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_12
timestamp 1621261055
transform 1 0 2304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_20
timestamp 1621261055
transform 1 0 3072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_4
timestamp 1621261055
transform 1 0 1536 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_12
timestamp 1621261055
transform 1 0 2304 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_20
timestamp 1621261055
transform 1 0 3072 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_29
timestamp 1621261055
transform 1 0 3936 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_28
timestamp 1621261055
transform 1 0 3840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_342
timestamp 1621261055
transform 1 0 3840 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_37
timestamp 1621261055
transform 1 0 4704 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_44
timestamp 1621261055
transform 1 0 5376 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_36
timestamp 1621261055
transform 1 0 4608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_53
timestamp 1621261055
transform 1 0 6240 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_45
timestamp 1621261055
transform 1 0 5472 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_52
timestamp 1621261055
transform 1 0 6144 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_15_54
timestamp 1621261055
transform 1 0 6336 0 1 12654
box -38 -49 134 715
use CLKBUF1  CLKBUF1
timestamp 1624893035
transform 1 0 7680 0 1 12654
box 0 -48 2592 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_332
timestamp 1621261055
transform 1 0 6432 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_53
timestamp 1621261055
transform 1 0 7488 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_56
timestamp 1621261055
transform 1 0 6528 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_64
timestamp 1621261055
transform 1 0 7296 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_61
timestamp 1621261055
transform 1 0 7008 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_69
timestamp 1621261055
transform 1 0 7776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_77
timestamp 1621261055
transform 1 0 8544 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_81
timestamp 1621261055
transform 1 0 8928 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_343
timestamp 1621261055
transform 1 0 9120 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_95
timestamp 1621261055
transform 1 0 10272 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_103
timestamp 1621261055
transform 1 0 11040 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_107
timestamp 1621261055
transform 1 0 11424 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_84
timestamp 1621261055
transform 1 0 9216 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_92
timestamp 1621261055
transform 1 0 9984 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_100
timestamp 1621261055
transform 1 0 10752 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_108
timestamp 1621261055
transform 1 0 11520 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_333
timestamp 1621261055
transform 1 0 11712 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_15_109
timestamp 1621261055
transform 1 0 11616 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_111
timestamp 1621261055
transform 1 0 11808 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_119
timestamp 1621261055
transform 1 0 12576 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_127
timestamp 1621261055
transform 1 0 13344 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_135
timestamp 1621261055
transform 1 0 14112 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_116
timestamp 1621261055
transform 1 0 12288 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_124
timestamp 1621261055
transform 1 0 13056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_132
timestamp 1621261055
transform 1 0 13824 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_16_139
timestamp 1621261055
transform 1 0 14496 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_136
timestamp 1621261055
transform 1 0 14208 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_143
timestamp 1621261055
transform 1 0 14880 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_344
timestamp 1621261055
transform 1 0 14400 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _146_
timestamp 1621261055
transform 1 0 14880 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_146
timestamp 1621261055
transform 1 0 15168 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_151
timestamp 1621261055
transform 1 0 15648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_154
timestamp 1621261055
transform 1 0 15936 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_159
timestamp 1621261055
transform 1 0 16416 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_162
timestamp 1621261055
transform 1 0 16704 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_334
timestamp 1621261055
transform 1 0 16992 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_163
timestamp 1621261055
transform 1 0 16800 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_166
timestamp 1621261055
transform 1 0 17088 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_174
timestamp 1621261055
transform 1 0 17856 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_182
timestamp 1621261055
transform 1 0 18624 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_170
timestamp 1621261055
transform 1 0 17472 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_178
timestamp 1621261055
transform 1 0 18240 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_186
timestamp 1621261055
transform 1 0 19008 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_194
timestamp 1621261055
transform 1 0 19776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_192
timestamp 1621261055
transform 1 0 19584 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_190
timestamp 1621261055
transform 1 0 19392 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_190
timestamp 1621261055
transform 1 0 19392 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_345
timestamp 1621261055
transform 1 0 19680 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_202
timestamp 1621261055
transform 1 0 20544 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_206
timestamp 1621261055
transform 1 0 20928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_198
timestamp 1621261055
transform 1 0 20160 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_210
timestamp 1621261055
transform 1 0 21312 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_214
timestamp 1621261055
transform 1 0 21696 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_335
timestamp 1621261055
transform 1 0 22272 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_218
timestamp 1621261055
transform 1 0 22080 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_221
timestamp 1621261055
transform 1 0 22368 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_229
timestamp 1621261055
transform 1 0 23136 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_237
timestamp 1621261055
transform 1 0 23904 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_218
timestamp 1621261055
transform 1 0 22080 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_226
timestamp 1621261055
transform 1 0 22848 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_234
timestamp 1621261055
transform 1 0 23616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_242
timestamp 1621261055
transform 1 0 24384 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_249
timestamp 1621261055
transform 1 0 25056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_246
timestamp 1621261055
transform 1 0 24768 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_245
timestamp 1621261055
transform 1 0 24672 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_346
timestamp 1621261055
transform 1 0 24960 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_257
timestamp 1621261055
transform 1 0 25824 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_253
timestamp 1621261055
transform 1 0 25440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_265
timestamp 1621261055
transform 1 0 26592 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_267
timestamp 1621261055
transform 1 0 26784 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_263
timestamp 1621261055
transform 1 0 26400 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_261
timestamp 1621261055
transform 1 0 26208 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _124_
timestamp 1621261055
transform 1 0 26496 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_336
timestamp 1621261055
transform 1 0 27552 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_276
timestamp 1621261055
transform 1 0 27648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_284
timestamp 1621261055
transform 1 0 28416 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_292
timestamp 1621261055
transform 1 0 29184 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_273
timestamp 1621261055
transform 1 0 27360 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_281
timestamp 1621261055
transform 1 0 28128 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_289
timestamp 1621261055
transform 1 0 28896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_297
timestamp 1621261055
transform 1 0 29664 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_347
timestamp 1621261055
transform 1 0 30240 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_300
timestamp 1621261055
transform 1 0 29952 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_308
timestamp 1621261055
transform 1 0 30720 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_316
timestamp 1621261055
transform 1 0 31488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_324
timestamp 1621261055
transform 1 0 32256 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_301
timestamp 1621261055
transform 1 0 30048 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_304
timestamp 1621261055
transform 1 0 30336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_312
timestamp 1621261055
transform 1 0 31104 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_320
timestamp 1621261055
transform 1 0 31872 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_337
timestamp 1621261055
transform 1 0 32832 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_328
timestamp 1621261055
transform 1 0 32640 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_331
timestamp 1621261055
transform 1 0 32928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_339
timestamp 1621261055
transform 1 0 33696 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_347
timestamp 1621261055
transform 1 0 34464 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_328
timestamp 1621261055
transform 1 0 32640 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_336
timestamp 1621261055
transform 1 0 33408 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_344
timestamp 1621261055
transform 1 0 34176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_348
timestamp 1621261055
transform 1 0 35520 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_355
timestamp 1621261055
transform 1 0 35232 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_363
timestamp 1621261055
transform 1 0 36000 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_371
timestamp 1621261055
transform 1 0 36768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_352
timestamp 1621261055
transform 1 0 34944 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_356
timestamp 1621261055
transform 1 0 35328 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_359
timestamp 1621261055
transform 1 0 35616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_367
timestamp 1621261055
transform 1 0 36384 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_375
timestamp 1621261055
transform 1 0 37152 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_338
timestamp 1621261055
transform 1 0 38112 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_379
timestamp 1621261055
transform 1 0 37536 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_383
timestamp 1621261055
transform 1 0 37920 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_386
timestamp 1621261055
transform 1 0 38208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_394
timestamp 1621261055
transform 1 0 38976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_402
timestamp 1621261055
transform 1 0 39744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_383
timestamp 1621261055
transform 1 0 37920 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_391
timestamp 1621261055
transform 1 0 38688 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_399
timestamp 1621261055
transform 1 0 39456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_349
timestamp 1621261055
transform 1 0 40800 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_410
timestamp 1621261055
transform 1 0 40512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_418
timestamp 1621261055
transform 1 0 41280 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_426
timestamp 1621261055
transform 1 0 42048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_407
timestamp 1621261055
transform 1 0 40224 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_411
timestamp 1621261055
transform 1 0 40608 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_414
timestamp 1621261055
transform 1 0 40896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_422
timestamp 1621261055
transform 1 0 41664 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_430
timestamp 1621261055
transform 1 0 42432 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_339
timestamp 1621261055
transform 1 0 43392 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_15_434
timestamp 1621261055
transform 1 0 42816 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_438
timestamp 1621261055
transform 1 0 43200 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_441
timestamp 1621261055
transform 1 0 43488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_449
timestamp 1621261055
transform 1 0 44256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_457
timestamp 1621261055
transform 1 0 45024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_438
timestamp 1621261055
transform 1 0 43200 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_446
timestamp 1621261055
transform 1 0 43968 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_454
timestamp 1621261055
transform 1 0 44736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_466
timestamp 1621261055
transform 1 0 45888 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_462
timestamp 1621261055
transform 1 0 45504 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_465
timestamp 1621261055
transform 1 0 45792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_469
timestamp 1621261055
transform 1 0 46176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_473
timestamp 1621261055
transform 1 0 46560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_350
timestamp 1621261055
transform 1 0 46080 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_485
timestamp 1621261055
transform 1 0 47712 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_479
timestamp 1621261055
transform 1 0 47136 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_477
timestamp 1621261055
transform 1 0 46944 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_481
timestamp 1621261055
transform 1 0 47328 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_79
timestamp 1621261055
transform 1 0 47232 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _055_
timestamp 1621261055
transform 1 0 47424 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_493
timestamp 1621261055
transform 1 0 48480 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_493
timestamp 1621261055
transform 1 0 48480 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_489
timestamp 1621261055
transform 1 0 48096 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_501
timestamp 1621261055
transform 1 0 49248 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_503
timestamp 1621261055
transform 1 0 49440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_496
timestamp 1621261055
transform 1 0 48768 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_6
timestamp 1621261055
transform 1 0 48960 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_340
timestamp 1621261055
transform 1 0 48672 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _005_
timestamp 1621261055
transform 1 0 49152 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_509
timestamp 1621261055
transform 1 0 50016 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_511
timestamp 1621261055
transform 1 0 50208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_351
timestamp 1621261055
transform 1 0 51360 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_15_519
timestamp 1621261055
transform 1 0 50976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_527
timestamp 1621261055
transform 1 0 51744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_535
timestamp 1621261055
transform 1 0 52512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_517
timestamp 1621261055
transform 1 0 50784 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_521
timestamp 1621261055
transform 1 0 51168 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_524
timestamp 1621261055
transform 1 0 51456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_532
timestamp 1621261055
transform 1 0 52224 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_540
timestamp 1621261055
transform 1 0 52992 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_548
timestamp 1621261055
transform 1 0 53760 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_549
timestamp 1621261055
transform 1 0 53856 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_547
timestamp 1621261055
transform 1 0 53664 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_543
timestamp 1621261055
transform 1 0 53280 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_556
timestamp 1621261055
transform 1 0 54528 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_551
timestamp 1621261055
transform 1 0 54048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_341
timestamp 1621261055
transform 1 0 53952 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_564
timestamp 1621261055
transform 1 0 55296 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_559
timestamp 1621261055
transform 1 0 54816 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_567
timestamp 1621261055
transform 1 0 55584 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_576
timestamp 1621261055
transform 1 0 56448 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_572
timestamp 1621261055
transform 1 0 56064 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_575
timestamp 1621261055
transform 1 0 56352 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_579
timestamp 1621261055
transform 1 0 56736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_583
timestamp 1621261055
transform 1 0 57120 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_352
timestamp 1621261055
transform 1 0 56640 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_587
timestamp 1621261055
transform 1 0 57504 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_593
timestamp 1621261055
transform 1 0 58080 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_15_589
timestamp 1621261055
transform 1 0 57696 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_587
timestamp 1621261055
transform 1 0 57504 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _090_
timestamp 1621261055
transform 1 0 57792 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_31
timestamp 1621261055
transform -1 0 58848 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_33
timestamp 1621261055
transform -1 0 58848 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_595
timestamp 1621261055
transform 1 0 58272 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _031_
timestamp 1621261055
transform 1 0 3648 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_34
timestamp 1621261055
transform 1 0 1152 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_18
timestamp 1621261055
transform 1 0 3456 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_4
timestamp 1621261055
transform 1 0 1536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_12
timestamp 1621261055
transform 1 0 2304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_20
timestamp 1621261055
transform 1 0 3072 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _003_
timestamp 1621261055
transform -1 0 4800 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_4
timestamp 1621261055
transform -1 0 4512 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_17_29
timestamp 1621261055
transform 1 0 3936 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_38
timestamp 1621261055
transform 1 0 4800 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_46
timestamp 1621261055
transform 1 0 5568 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_17_54
timestamp 1621261055
transform 1 0 6336 0 1 13986
box -38 -49 134 715
use INV  INV
timestamp 1624893035
transform 1 0 7680 0 1 13986
box 0 -48 576 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_353
timestamp 1621261055
transform 1 0 6432 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_57
timestamp 1621261055
transform 1 0 7488 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_56
timestamp 1621261055
transform 1 0 6528 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_64
timestamp 1621261055
transform 1 0 7296 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_74
timestamp 1621261055
transform 1 0 8256 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_82
timestamp 1621261055
transform 1 0 9024 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_90
timestamp 1621261055
transform 1 0 9792 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_98
timestamp 1621261055
transform 1 0 10560 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_106
timestamp 1621261055
transform 1 0 11328 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _141_
timestamp 1621261055
transform 1 0 12480 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_354
timestamp 1621261055
transform 1 0 11712 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_111
timestamp 1621261055
transform 1 0 11808 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_115
timestamp 1621261055
transform 1 0 12192 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_117
timestamp 1621261055
transform 1 0 12384 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_121
timestamp 1621261055
transform 1 0 12768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_129
timestamp 1621261055
transform 1 0 13536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_137
timestamp 1621261055
transform 1 0 14304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_145
timestamp 1621261055
transform 1 0 15072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_153
timestamp 1621261055
transform 1 0 15840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_161
timestamp 1621261055
transform 1 0 16608 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _053_
timestamp 1621261055
transform 1 0 17568 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_355
timestamp 1621261055
transform 1 0 16992 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_72
timestamp 1621261055
transform 1 0 17376 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_166
timestamp 1621261055
transform 1 0 17088 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_168
timestamp 1621261055
transform 1 0 17280 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_174
timestamp 1621261055
transform 1 0 17856 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_182
timestamp 1621261055
transform 1 0 18624 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_190
timestamp 1621261055
transform 1 0 19392 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_198
timestamp 1621261055
transform 1 0 20160 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_206
timestamp 1621261055
transform 1 0 20928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_214
timestamp 1621261055
transform 1 0 21696 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_356
timestamp 1621261055
transform 1 0 22272 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_218
timestamp 1621261055
transform 1 0 22080 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_221
timestamp 1621261055
transform 1 0 22368 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_229
timestamp 1621261055
transform 1 0 23136 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_237
timestamp 1621261055
transform 1 0 23904 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_245
timestamp 1621261055
transform 1 0 24672 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_253
timestamp 1621261055
transform 1 0 25440 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_261
timestamp 1621261055
transform 1 0 26208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_269
timestamp 1621261055
transform 1 0 26976 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_357
timestamp 1621261055
transform 1 0 27552 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_273
timestamp 1621261055
transform 1 0 27360 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_276
timestamp 1621261055
transform 1 0 27648 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_284
timestamp 1621261055
transform 1 0 28416 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_292
timestamp 1621261055
transform 1 0 29184 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_300
timestamp 1621261055
transform 1 0 29952 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_308
timestamp 1621261055
transform 1 0 30720 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_316
timestamp 1621261055
transform 1 0 31488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_324
timestamp 1621261055
transform 1 0 32256 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_358
timestamp 1621261055
transform 1 0 32832 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_328
timestamp 1621261055
transform 1 0 32640 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_331
timestamp 1621261055
transform 1 0 32928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_339
timestamp 1621261055
transform 1 0 33696 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_347
timestamp 1621261055
transform 1 0 34464 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_355
timestamp 1621261055
transform 1 0 35232 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_363
timestamp 1621261055
transform 1 0 36000 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_371
timestamp 1621261055
transform 1 0 36768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_359
timestamp 1621261055
transform 1 0 38112 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_379
timestamp 1621261055
transform 1 0 37536 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_383
timestamp 1621261055
transform 1 0 37920 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_386
timestamp 1621261055
transform 1 0 38208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_394
timestamp 1621261055
transform 1 0 38976 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_402
timestamp 1621261055
transform 1 0 39744 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_410
timestamp 1621261055
transform 1 0 40512 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_418
timestamp 1621261055
transform 1 0 41280 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_426
timestamp 1621261055
transform 1 0 42048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_360
timestamp 1621261055
transform 1 0 43392 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_434
timestamp 1621261055
transform 1 0 42816 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_438
timestamp 1621261055
transform 1 0 43200 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_441
timestamp 1621261055
transform 1 0 43488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_449
timestamp 1621261055
transform 1 0 44256 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_457
timestamp 1621261055
transform 1 0 45024 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_465
timestamp 1621261055
transform 1 0 45792 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_473
timestamp 1621261055
transform 1 0 46560 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_481
timestamp 1621261055
transform 1 0 47328 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_361
timestamp 1621261055
transform 1 0 48672 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_489
timestamp 1621261055
transform 1 0 48096 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_493
timestamp 1621261055
transform 1 0 48480 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_496
timestamp 1621261055
transform 1 0 48768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_504
timestamp 1621261055
transform 1 0 49536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_512
timestamp 1621261055
transform 1 0 50304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_520
timestamp 1621261055
transform 1 0 51072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_528
timestamp 1621261055
transform 1 0 51840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_536
timestamp 1621261055
transform 1 0 52608 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_362
timestamp 1621261055
transform 1 0 53952 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_544
timestamp 1621261055
transform 1 0 53376 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_548
timestamp 1621261055
transform 1 0 53760 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_551
timestamp 1621261055
transform 1 0 54048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_559
timestamp 1621261055
transform 1 0 54816 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_567
timestamp 1621261055
transform 1 0 55584 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_575
timestamp 1621261055
transform 1 0 56352 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_583
timestamp 1621261055
transform 1 0 57120 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_591
timestamp 1621261055
transform 1 0 57888 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_35
timestamp 1621261055
transform -1 0 58848 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_595
timestamp 1621261055
transform 1 0 58272 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_36
timestamp 1621261055
transform 1 0 1152 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_4
timestamp 1621261055
transform 1 0 1536 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_12
timestamp 1621261055
transform 1 0 2304 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_20
timestamp 1621261055
transform 1 0 3072 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_363
timestamp 1621261055
transform 1 0 3840 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_29
timestamp 1621261055
transform 1 0 3936 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_37
timestamp 1621261055
transform 1 0 4704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_45
timestamp 1621261055
transform 1 0 5472 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_53
timestamp 1621261055
transform 1 0 6240 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_61
timestamp 1621261055
transform 1 0 7008 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_69
timestamp 1621261055
transform 1 0 7776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_77
timestamp 1621261055
transform 1 0 8544 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_81
timestamp 1621261055
transform 1 0 8928 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_364
timestamp 1621261055
transform 1 0 9120 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_84
timestamp 1621261055
transform 1 0 9216 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_92
timestamp 1621261055
transform 1 0 9984 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_100
timestamp 1621261055
transform 1 0 10752 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_108
timestamp 1621261055
transform 1 0 11520 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _022_
timestamp 1621261055
transform -1 0 12672 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_0
timestamp 1621261055
transform -1 0 12384 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_112
timestamp 1621261055
transform 1 0 11904 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_114
timestamp 1621261055
transform 1 0 12096 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_120
timestamp 1621261055
transform 1 0 12672 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_128
timestamp 1621261055
transform 1 0 13440 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_365
timestamp 1621261055
transform 1 0 14400 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_136
timestamp 1621261055
transform 1 0 14208 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_139
timestamp 1621261055
transform 1 0 14496 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_147
timestamp 1621261055
transform 1 0 15264 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_155
timestamp 1621261055
transform 1 0 16032 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_163
timestamp 1621261055
transform 1 0 16800 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_171
timestamp 1621261055
transform 1 0 17568 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_179
timestamp 1621261055
transform 1 0 18336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_187
timestamp 1621261055
transform 1 0 19104 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_366
timestamp 1621261055
transform 1 0 19680 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_191
timestamp 1621261055
transform 1 0 19488 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_194
timestamp 1621261055
transform 1 0 19776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_202
timestamp 1621261055
transform 1 0 20544 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_210
timestamp 1621261055
transform 1 0 21312 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _045_
timestamp 1621261055
transform -1 0 24480 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _198_
timestamp 1621261055
transform 1 0 23520 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_37
timestamp 1621261055
transform -1 0 24192 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_218
timestamp 1621261055
transform 1 0 22080 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_226
timestamp 1621261055
transform 1 0 22848 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_230
timestamp 1621261055
transform 1 0 23232 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_232
timestamp 1621261055
transform 1 0 23424 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_236
timestamp 1621261055
transform 1 0 23808 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_18_243
timestamp 1621261055
transform 1 0 24480 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_367
timestamp 1621261055
transform 1 0 24960 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_18_247
timestamp 1621261055
transform 1 0 24864 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_249
timestamp 1621261055
transform 1 0 25056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_257
timestamp 1621261055
transform 1 0 25824 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_265
timestamp 1621261055
transform 1 0 26592 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_273
timestamp 1621261055
transform 1 0 27360 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_281
timestamp 1621261055
transform 1 0 28128 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_289
timestamp 1621261055
transform 1 0 28896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_297
timestamp 1621261055
transform 1 0 29664 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_368
timestamp 1621261055
transform 1 0 30240 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_301
timestamp 1621261055
transform 1 0 30048 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_304
timestamp 1621261055
transform 1 0 30336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_312
timestamp 1621261055
transform 1 0 31104 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_320
timestamp 1621261055
transform 1 0 31872 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_328
timestamp 1621261055
transform 1 0 32640 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_336
timestamp 1621261055
transform 1 0 33408 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_344
timestamp 1621261055
transform 1 0 34176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_369
timestamp 1621261055
transform 1 0 35520 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_352
timestamp 1621261055
transform 1 0 34944 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_356
timestamp 1621261055
transform 1 0 35328 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_359
timestamp 1621261055
transform 1 0 35616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_367
timestamp 1621261055
transform 1 0 36384 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_375
timestamp 1621261055
transform 1 0 37152 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_383
timestamp 1621261055
transform 1 0 37920 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_391
timestamp 1621261055
transform 1 0 38688 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_399
timestamp 1621261055
transform 1 0 39456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_370
timestamp 1621261055
transform 1 0 40800 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_407
timestamp 1621261055
transform 1 0 40224 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_411
timestamp 1621261055
transform 1 0 40608 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_414
timestamp 1621261055
transform 1 0 40896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_422
timestamp 1621261055
transform 1 0 41664 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_430
timestamp 1621261055
transform 1 0 42432 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_438
timestamp 1621261055
transform 1 0 43200 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_446
timestamp 1621261055
transform 1 0 43968 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_454
timestamp 1621261055
transform 1 0 44736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_371
timestamp 1621261055
transform 1 0 46080 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_462
timestamp 1621261055
transform 1 0 45504 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_466
timestamp 1621261055
transform 1 0 45888 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_469
timestamp 1621261055
transform 1 0 46176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_477
timestamp 1621261055
transform 1 0 46944 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_485
timestamp 1621261055
transform 1 0 47712 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_493
timestamp 1621261055
transform 1 0 48480 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_501
timestamp 1621261055
transform 1 0 49248 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_509
timestamp 1621261055
transform 1 0 50016 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_372
timestamp 1621261055
transform 1 0 51360 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_517
timestamp 1621261055
transform 1 0 50784 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_521
timestamp 1621261055
transform 1 0 51168 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_524
timestamp 1621261055
transform 1 0 51456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_532
timestamp 1621261055
transform 1 0 52224 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_540
timestamp 1621261055
transform 1 0 52992 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_548
timestamp 1621261055
transform 1 0 53760 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_556
timestamp 1621261055
transform 1 0 54528 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_564
timestamp 1621261055
transform 1 0 55296 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _034_
timestamp 1621261055
transform 1 0 57792 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_373
timestamp 1621261055
transform 1 0 56640 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_27
timestamp 1621261055
transform 1 0 57600 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_18_572
timestamp 1621261055
transform 1 0 56064 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_576
timestamp 1621261055
transform 1 0 56448 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_579
timestamp 1621261055
transform 1 0 56736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_18_587
timestamp 1621261055
transform 1 0 57504 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_18_593
timestamp 1621261055
transform 1 0 58080 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_37
timestamp 1621261055
transform -1 0 58848 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_38
timestamp 1621261055
transform 1 0 1152 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_4
timestamp 1621261055
transform 1 0 1536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_12
timestamp 1621261055
transform 1 0 2304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_20
timestamp 1621261055
transform 1 0 3072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_28
timestamp 1621261055
transform 1 0 3840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_36
timestamp 1621261055
transform 1 0 4608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_44
timestamp 1621261055
transform 1 0 5376 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_52
timestamp 1621261055
transform 1 0 6144 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_54
timestamp 1621261055
transform 1 0 6336 0 1 15318
box -38 -49 134 715
use INVX1  INVX1
timestamp 1624893035
transform 1 0 7680 0 1 15318
box 0 -48 576 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_374
timestamp 1621261055
transform 1 0 6432 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_61
timestamp 1621261055
transform 1 0 7488 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_56
timestamp 1621261055
transform 1 0 6528 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_64
timestamp 1621261055
transform 1 0 7296 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_74
timestamp 1621261055
transform 1 0 8256 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_82
timestamp 1621261055
transform 1 0 9024 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_90
timestamp 1621261055
transform 1 0 9792 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_98
timestamp 1621261055
transform 1 0 10560 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_106
timestamp 1621261055
transform 1 0 11328 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_375
timestamp 1621261055
transform 1 0 11712 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_111
timestamp 1621261055
transform 1 0 11808 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_119
timestamp 1621261055
transform 1 0 12576 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_127
timestamp 1621261055
transform 1 0 13344 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_135
timestamp 1621261055
transform 1 0 14112 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_143
timestamp 1621261055
transform 1 0 14880 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_151
timestamp 1621261055
transform 1 0 15648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_159
timestamp 1621261055
transform 1 0 16416 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_376
timestamp 1621261055
transform 1 0 16992 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_163
timestamp 1621261055
transform 1 0 16800 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_166
timestamp 1621261055
transform 1 0 17088 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_174
timestamp 1621261055
transform 1 0 17856 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_182
timestamp 1621261055
transform 1 0 18624 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_190
timestamp 1621261055
transform 1 0 19392 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_198
timestamp 1621261055
transform 1 0 20160 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_206
timestamp 1621261055
transform 1 0 20928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_214
timestamp 1621261055
transform 1 0 21696 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_377
timestamp 1621261055
transform 1 0 22272 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_218
timestamp 1621261055
transform 1 0 22080 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_221
timestamp 1621261055
transform 1 0 22368 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_229
timestamp 1621261055
transform 1 0 23136 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_237
timestamp 1621261055
transform 1 0 23904 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_245
timestamp 1621261055
transform 1 0 24672 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_253
timestamp 1621261055
transform 1 0 25440 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_261
timestamp 1621261055
transform 1 0 26208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_269
timestamp 1621261055
transform 1 0 26976 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_378
timestamp 1621261055
transform 1 0 27552 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_273
timestamp 1621261055
transform 1 0 27360 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_276
timestamp 1621261055
transform 1 0 27648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_284
timestamp 1621261055
transform 1 0 28416 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_292
timestamp 1621261055
transform 1 0 29184 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_300
timestamp 1621261055
transform 1 0 29952 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_308
timestamp 1621261055
transform 1 0 30720 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_316
timestamp 1621261055
transform 1 0 31488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_324
timestamp 1621261055
transform 1 0 32256 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_379
timestamp 1621261055
transform 1 0 32832 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_328
timestamp 1621261055
transform 1 0 32640 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_331
timestamp 1621261055
transform 1 0 32928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_339
timestamp 1621261055
transform 1 0 33696 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_347
timestamp 1621261055
transform 1 0 34464 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_355
timestamp 1621261055
transform 1 0 35232 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_363
timestamp 1621261055
transform 1 0 36000 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_371
timestamp 1621261055
transform 1 0 36768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_380
timestamp 1621261055
transform 1 0 38112 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_379
timestamp 1621261055
transform 1 0 37536 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_383
timestamp 1621261055
transform 1 0 37920 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_386
timestamp 1621261055
transform 1 0 38208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_394
timestamp 1621261055
transform 1 0 38976 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_402
timestamp 1621261055
transform 1 0 39744 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_410
timestamp 1621261055
transform 1 0 40512 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_418
timestamp 1621261055
transform 1 0 41280 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_426
timestamp 1621261055
transform 1 0 42048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_381
timestamp 1621261055
transform 1 0 43392 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_434
timestamp 1621261055
transform 1 0 42816 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_438
timestamp 1621261055
transform 1 0 43200 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_441
timestamp 1621261055
transform 1 0 43488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_449
timestamp 1621261055
transform 1 0 44256 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_457
timestamp 1621261055
transform 1 0 45024 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _001_
timestamp 1621261055
transform 1 0 47040 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_2
timestamp 1621261055
transform 1 0 46848 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_465
timestamp 1621261055
transform 1 0 45792 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_473
timestamp 1621261055
transform 1 0 46560 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_475
timestamp 1621261055
transform 1 0 46752 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_481
timestamp 1621261055
transform 1 0 47328 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_382
timestamp 1621261055
transform 1 0 48672 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_489
timestamp 1621261055
transform 1 0 48096 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_493
timestamp 1621261055
transform 1 0 48480 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_496
timestamp 1621261055
transform 1 0 48768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_504
timestamp 1621261055
transform 1 0 49536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_512
timestamp 1621261055
transform 1 0 50304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_520
timestamp 1621261055
transform 1 0 51072 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_528
timestamp 1621261055
transform 1 0 51840 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_536
timestamp 1621261055
transform 1 0 52608 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_383
timestamp 1621261055
transform 1 0 53952 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_544
timestamp 1621261055
transform 1 0 53376 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_548
timestamp 1621261055
transform 1 0 53760 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_551
timestamp 1621261055
transform 1 0 54048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_559
timestamp 1621261055
transform 1 0 54816 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_567
timestamp 1621261055
transform 1 0 55584 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_575
timestamp 1621261055
transform 1 0 56352 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_583
timestamp 1621261055
transform 1 0 57120 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_591
timestamp 1621261055
transform 1 0 57888 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_39
timestamp 1621261055
transform -1 0 58848 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_595
timestamp 1621261055
transform 1 0 58272 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_40
timestamp 1621261055
transform 1 0 1152 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_20_4
timestamp 1621261055
transform 1 0 1536 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_12
timestamp 1621261055
transform 1 0 2304 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_20
timestamp 1621261055
transform 1 0 3072 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_384
timestamp 1621261055
transform 1 0 3840 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_29
timestamp 1621261055
transform 1 0 3936 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_37
timestamp 1621261055
transform 1 0 4704 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_45
timestamp 1621261055
transform 1 0 5472 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_53
timestamp 1621261055
transform 1 0 6240 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_61
timestamp 1621261055
transform 1 0 7008 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_69
timestamp 1621261055
transform 1 0 7776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_77
timestamp 1621261055
transform 1 0 8544 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_81
timestamp 1621261055
transform 1 0 8928 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_385
timestamp 1621261055
transform 1 0 9120 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_84
timestamp 1621261055
transform 1 0 9216 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_92
timestamp 1621261055
transform 1 0 9984 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_100
timestamp 1621261055
transform 1 0 10752 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_108
timestamp 1621261055
transform 1 0 11520 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_116
timestamp 1621261055
transform 1 0 12288 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_124
timestamp 1621261055
transform 1 0 13056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_132
timestamp 1621261055
transform 1 0 13824 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_386
timestamp 1621261055
transform 1 0 14400 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_136
timestamp 1621261055
transform 1 0 14208 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_139
timestamp 1621261055
transform 1 0 14496 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_147
timestamp 1621261055
transform 1 0 15264 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_155
timestamp 1621261055
transform 1 0 16032 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_163
timestamp 1621261055
transform 1 0 16800 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_171
timestamp 1621261055
transform 1 0 17568 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_179
timestamp 1621261055
transform 1 0 18336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_187
timestamp 1621261055
transform 1 0 19104 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_387
timestamp 1621261055
transform 1 0 19680 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_191
timestamp 1621261055
transform 1 0 19488 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_194
timestamp 1621261055
transform 1 0 19776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_202
timestamp 1621261055
transform 1 0 20544 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_210
timestamp 1621261055
transform 1 0 21312 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_218
timestamp 1621261055
transform 1 0 22080 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_226
timestamp 1621261055
transform 1 0 22848 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_234
timestamp 1621261055
transform 1 0 23616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_242
timestamp 1621261055
transform 1 0 24384 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _157_
timestamp 1621261055
transform 1 0 26880 0 -1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_388
timestamp 1621261055
transform 1 0 24960 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_246
timestamp 1621261055
transform 1 0 24768 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_249
timestamp 1621261055
transform 1 0 25056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_257
timestamp 1621261055
transform 1 0 25824 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_265
timestamp 1621261055
transform 1 0 26592 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_20_267
timestamp 1621261055
transform 1 0 26784 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_271
timestamp 1621261055
transform 1 0 27168 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_279
timestamp 1621261055
transform 1 0 27936 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_287
timestamp 1621261055
transform 1 0 28704 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_295
timestamp 1621261055
transform 1 0 29472 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_389
timestamp 1621261055
transform 1 0 30240 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_304
timestamp 1621261055
transform 1 0 30336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_312
timestamp 1621261055
transform 1 0 31104 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_320
timestamp 1621261055
transform 1 0 31872 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_328
timestamp 1621261055
transform 1 0 32640 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_336
timestamp 1621261055
transform 1 0 33408 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_344
timestamp 1621261055
transform 1 0 34176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_390
timestamp 1621261055
transform 1 0 35520 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_352
timestamp 1621261055
transform 1 0 34944 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_356
timestamp 1621261055
transform 1 0 35328 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_359
timestamp 1621261055
transform 1 0 35616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_367
timestamp 1621261055
transform 1 0 36384 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_375
timestamp 1621261055
transform 1 0 37152 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_383
timestamp 1621261055
transform 1 0 37920 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_391
timestamp 1621261055
transform 1 0 38688 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_399
timestamp 1621261055
transform 1 0 39456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_391
timestamp 1621261055
transform 1 0 40800 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_407
timestamp 1621261055
transform 1 0 40224 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_411
timestamp 1621261055
transform 1 0 40608 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_414
timestamp 1621261055
transform 1 0 40896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_422
timestamp 1621261055
transform 1 0 41664 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_430
timestamp 1621261055
transform 1 0 42432 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_438
timestamp 1621261055
transform 1 0 43200 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_446
timestamp 1621261055
transform 1 0 43968 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_454
timestamp 1621261055
transform 1 0 44736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_392
timestamp 1621261055
transform 1 0 46080 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_462
timestamp 1621261055
transform 1 0 45504 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_466
timestamp 1621261055
transform 1 0 45888 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_469
timestamp 1621261055
transform 1 0 46176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_477
timestamp 1621261055
transform 1 0 46944 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_485
timestamp 1621261055
transform 1 0 47712 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_493
timestamp 1621261055
transform 1 0 48480 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_501
timestamp 1621261055
transform 1 0 49248 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_509
timestamp 1621261055
transform 1 0 50016 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_393
timestamp 1621261055
transform 1 0 51360 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_517
timestamp 1621261055
transform 1 0 50784 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_521
timestamp 1621261055
transform 1 0 51168 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_524
timestamp 1621261055
transform 1 0 51456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_532
timestamp 1621261055
transform 1 0 52224 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_540
timestamp 1621261055
transform 1 0 52992 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_548
timestamp 1621261055
transform 1 0 53760 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_556
timestamp 1621261055
transform 1 0 54528 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_564
timestamp 1621261055
transform 1 0 55296 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_394
timestamp 1621261055
transform 1 0 56640 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_20_572
timestamp 1621261055
transform 1 0 56064 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_576
timestamp 1621261055
transform 1 0 56448 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_579
timestamp 1621261055
transform 1 0 56736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_587
timestamp 1621261055
transform 1 0 57504 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_41
timestamp 1621261055
transform -1 0 58848 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_595
timestamp 1621261055
transform 1 0 58272 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_42
timestamp 1621261055
transform 1 0 1152 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_4
timestamp 1621261055
transform 1 0 1536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_12
timestamp 1621261055
transform 1 0 2304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_20
timestamp 1621261055
transform 1 0 3072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _214_
timestamp 1621261055
transform 1 0 5760 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_21_28
timestamp 1621261055
transform 1 0 3840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_36
timestamp 1621261055
transform 1 0 4608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_44
timestamp 1621261055
transform 1 0 5376 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_21_51
timestamp 1621261055
transform 1 0 6048 0 1 16650
box -38 -49 422 715
use INVX2  INVX2
timestamp 1624893035
transform 1 0 7680 0 1 16650
box 0 -48 576 714
use sky130_fd_sc_ls__conb_1  _164_
timestamp 1621261055
transform 1 0 6912 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_395
timestamp 1621261055
transform 1 0 6432 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_66
timestamp 1621261055
transform 1 0 7488 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_21_56
timestamp 1621261055
transform 1 0 6528 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_63
timestamp 1621261055
transform 1 0 7200 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_65
timestamp 1621261055
transform 1 0 7392 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_74
timestamp 1621261055
transform 1 0 8256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_82
timestamp 1621261055
transform 1 0 9024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_90
timestamp 1621261055
transform 1 0 9792 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_98
timestamp 1621261055
transform 1 0 10560 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_106
timestamp 1621261055
transform 1 0 11328 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_396
timestamp 1621261055
transform 1 0 11712 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_111
timestamp 1621261055
transform 1 0 11808 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_119
timestamp 1621261055
transform 1 0 12576 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_127
timestamp 1621261055
transform 1 0 13344 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_135
timestamp 1621261055
transform 1 0 14112 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_143
timestamp 1621261055
transform 1 0 14880 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_151
timestamp 1621261055
transform 1 0 15648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_159
timestamp 1621261055
transform 1 0 16416 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_397
timestamp 1621261055
transform 1 0 16992 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_163
timestamp 1621261055
transform 1 0 16800 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_166
timestamp 1621261055
transform 1 0 17088 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_174
timestamp 1621261055
transform 1 0 17856 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_182
timestamp 1621261055
transform 1 0 18624 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_190
timestamp 1621261055
transform 1 0 19392 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_198
timestamp 1621261055
transform 1 0 20160 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_206
timestamp 1621261055
transform 1 0 20928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_214
timestamp 1621261055
transform 1 0 21696 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_398
timestamp 1621261055
transform 1 0 22272 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_218
timestamp 1621261055
transform 1 0 22080 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_221
timestamp 1621261055
transform 1 0 22368 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_229
timestamp 1621261055
transform 1 0 23136 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_237
timestamp 1621261055
transform 1 0 23904 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_245
timestamp 1621261055
transform 1 0 24672 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_253
timestamp 1621261055
transform 1 0 25440 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_261
timestamp 1621261055
transform 1 0 26208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_269
timestamp 1621261055
transform 1 0 26976 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_399
timestamp 1621261055
transform 1 0 27552 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_273
timestamp 1621261055
transform 1 0 27360 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_276
timestamp 1621261055
transform 1 0 27648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_284
timestamp 1621261055
transform 1 0 28416 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_292
timestamp 1621261055
transform 1 0 29184 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_300
timestamp 1621261055
transform 1 0 29952 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_308
timestamp 1621261055
transform 1 0 30720 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_316
timestamp 1621261055
transform 1 0 31488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_324
timestamp 1621261055
transform 1 0 32256 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_400
timestamp 1621261055
transform 1 0 32832 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_328
timestamp 1621261055
transform 1 0 32640 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_331
timestamp 1621261055
transform 1 0 32928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_339
timestamp 1621261055
transform 1 0 33696 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_347
timestamp 1621261055
transform 1 0 34464 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_355
timestamp 1621261055
transform 1 0 35232 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_363
timestamp 1621261055
transform 1 0 36000 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_371
timestamp 1621261055
transform 1 0 36768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_401
timestamp 1621261055
transform 1 0 38112 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_379
timestamp 1621261055
transform 1 0 37536 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_383
timestamp 1621261055
transform 1 0 37920 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_386
timestamp 1621261055
transform 1 0 38208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_394
timestamp 1621261055
transform 1 0 38976 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_402
timestamp 1621261055
transform 1 0 39744 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_410
timestamp 1621261055
transform 1 0 40512 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_418
timestamp 1621261055
transform 1 0 41280 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_426
timestamp 1621261055
transform 1 0 42048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_402
timestamp 1621261055
transform 1 0 43392 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_434
timestamp 1621261055
transform 1 0 42816 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_438
timestamp 1621261055
transform 1 0 43200 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_441
timestamp 1621261055
transform 1 0 43488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_449
timestamp 1621261055
transform 1 0 44256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_457
timestamp 1621261055
transform 1 0 45024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _091_
timestamp 1621261055
transform 1 0 46656 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_21_465
timestamp 1621261055
transform 1 0 45792 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_21_473
timestamp 1621261055
transform 1 0 46560 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_477
timestamp 1621261055
transform 1 0 46944 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_485
timestamp 1621261055
transform 1 0 47712 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_403
timestamp 1621261055
transform 1 0 48672 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_493
timestamp 1621261055
transform 1 0 48480 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_496
timestamp 1621261055
transform 1 0 48768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_504
timestamp 1621261055
transform 1 0 49536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_512
timestamp 1621261055
transform 1 0 50304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_520
timestamp 1621261055
transform 1 0 51072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_528
timestamp 1621261055
transform 1 0 51840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_536
timestamp 1621261055
transform 1 0 52608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_404
timestamp 1621261055
transform 1 0 53952 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_544
timestamp 1621261055
transform 1 0 53376 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_548
timestamp 1621261055
transform 1 0 53760 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_551
timestamp 1621261055
transform 1 0 54048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_559
timestamp 1621261055
transform 1 0 54816 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_567
timestamp 1621261055
transform 1 0 55584 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _178_
timestamp 1621261055
transform 1 0 55776 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _217_
timestamp 1621261055
transform 1 0 56544 0 1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_21_572
timestamp 1621261055
transform 1 0 56064 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_21_576
timestamp 1621261055
transform 1 0 56448 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_580
timestamp 1621261055
transform 1 0 56832 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_588
timestamp 1621261055
transform 1 0 57600 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_43
timestamp 1621261055
transform -1 0 58848 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_21_596
timestamp 1621261055
transform 1 0 58368 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _079_
timestamp 1621261055
transform 1 0 1728 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_44
timestamp 1621261055
transform 1 0 1152 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_4
timestamp 1621261055
transform 1 0 1536 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_9
timestamp 1621261055
transform 1 0 2016 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_17
timestamp 1621261055
transform 1 0 2784 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_25
timestamp 1621261055
transform 1 0 3552 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_22_27
timestamp 1621261055
transform 1 0 3744 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_405
timestamp 1621261055
transform 1 0 3840 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_29
timestamp 1621261055
transform 1 0 3936 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_37
timestamp 1621261055
transform 1 0 4704 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_45
timestamp 1621261055
transform 1 0 5472 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_53
timestamp 1621261055
transform 1 0 6240 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_61
timestamp 1621261055
transform 1 0 7008 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_69
timestamp 1621261055
transform 1 0 7776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_77
timestamp 1621261055
transform 1 0 8544 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_81
timestamp 1621261055
transform 1 0 8928 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_406
timestamp 1621261055
transform 1 0 9120 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_84
timestamp 1621261055
transform 1 0 9216 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_92
timestamp 1621261055
transform 1 0 9984 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_100
timestamp 1621261055
transform 1 0 10752 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_108
timestamp 1621261055
transform 1 0 11520 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_116
timestamp 1621261055
transform 1 0 12288 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_124
timestamp 1621261055
transform 1 0 13056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_132
timestamp 1621261055
transform 1 0 13824 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_407
timestamp 1621261055
transform 1 0 14400 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_136
timestamp 1621261055
transform 1 0 14208 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_139
timestamp 1621261055
transform 1 0 14496 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_147
timestamp 1621261055
transform 1 0 15264 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_155
timestamp 1621261055
transform 1 0 16032 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_163
timestamp 1621261055
transform 1 0 16800 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_171
timestamp 1621261055
transform 1 0 17568 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_179
timestamp 1621261055
transform 1 0 18336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_187
timestamp 1621261055
transform 1 0 19104 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_408
timestamp 1621261055
transform 1 0 19680 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_191
timestamp 1621261055
transform 1 0 19488 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_194
timestamp 1621261055
transform 1 0 19776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_202
timestamp 1621261055
transform 1 0 20544 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_210
timestamp 1621261055
transform 1 0 21312 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_218
timestamp 1621261055
transform 1 0 22080 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_226
timestamp 1621261055
transform 1 0 22848 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_234
timestamp 1621261055
transform 1 0 23616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_242
timestamp 1621261055
transform 1 0 24384 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_409
timestamp 1621261055
transform 1 0 24960 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_246
timestamp 1621261055
transform 1 0 24768 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_249
timestamp 1621261055
transform 1 0 25056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_257
timestamp 1621261055
transform 1 0 25824 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_265
timestamp 1621261055
transform 1 0 26592 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_273
timestamp 1621261055
transform 1 0 27360 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_281
timestamp 1621261055
transform 1 0 28128 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_289
timestamp 1621261055
transform 1 0 28896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_297
timestamp 1621261055
transform 1 0 29664 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _028_
timestamp 1621261055
transform 1 0 30720 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_410
timestamp 1621261055
transform 1 0 30240 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_8
timestamp 1621261055
transform 1 0 30528 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_301
timestamp 1621261055
transform 1 0 30048 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_304
timestamp 1621261055
transform 1 0 30336 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_311
timestamp 1621261055
transform 1 0 31008 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_319
timestamp 1621261055
transform 1 0 31776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_327
timestamp 1621261055
transform 1 0 32544 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_335
timestamp 1621261055
transform 1 0 33312 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_343
timestamp 1621261055
transform 1 0 34080 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_351
timestamp 1621261055
transform 1 0 34848 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_411
timestamp 1621261055
transform 1 0 35520 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_355
timestamp 1621261055
transform 1 0 35232 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_22_357
timestamp 1621261055
transform 1 0 35424 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_359
timestamp 1621261055
transform 1 0 35616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_367
timestamp 1621261055
transform 1 0 36384 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_375
timestamp 1621261055
transform 1 0 37152 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_383
timestamp 1621261055
transform 1 0 37920 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_391
timestamp 1621261055
transform 1 0 38688 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_399
timestamp 1621261055
transform 1 0 39456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_412
timestamp 1621261055
transform 1 0 40800 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_407
timestamp 1621261055
transform 1 0 40224 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_411
timestamp 1621261055
transform 1 0 40608 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_414
timestamp 1621261055
transform 1 0 40896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_422
timestamp 1621261055
transform 1 0 41664 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_430
timestamp 1621261055
transform 1 0 42432 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_438
timestamp 1621261055
transform 1 0 43200 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_446
timestamp 1621261055
transform 1 0 43968 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_454
timestamp 1621261055
transform 1 0 44736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_413
timestamp 1621261055
transform 1 0 46080 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_462
timestamp 1621261055
transform 1 0 45504 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_466
timestamp 1621261055
transform 1 0 45888 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_469
timestamp 1621261055
transform 1 0 46176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_477
timestamp 1621261055
transform 1 0 46944 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_485
timestamp 1621261055
transform 1 0 47712 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_493
timestamp 1621261055
transform 1 0 48480 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_501
timestamp 1621261055
transform 1 0 49248 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_509
timestamp 1621261055
transform 1 0 50016 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_414
timestamp 1621261055
transform 1 0 51360 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_517
timestamp 1621261055
transform 1 0 50784 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_521
timestamp 1621261055
transform 1 0 51168 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_524
timestamp 1621261055
transform 1 0 51456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_532
timestamp 1621261055
transform 1 0 52224 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_540
timestamp 1621261055
transform 1 0 52992 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_548
timestamp 1621261055
transform 1 0 53760 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_556
timestamp 1621261055
transform 1 0 54528 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_564
timestamp 1621261055
transform 1 0 55296 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_415
timestamp 1621261055
transform 1 0 56640 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_22_572
timestamp 1621261055
transform 1 0 56064 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_576
timestamp 1621261055
transform 1 0 56448 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_579
timestamp 1621261055
transform 1 0 56736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_587
timestamp 1621261055
transform 1 0 57504 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_45
timestamp 1621261055
transform -1 0 58848 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_595
timestamp 1621261055
transform 1 0 58272 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _201_
timestamp 1621261055
transform 1 0 1536 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_46
timestamp 1621261055
transform 1 0 1152 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_48
timestamp 1621261055
transform 1 0 1152 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_7
timestamp 1621261055
transform 1 0 1824 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_15
timestamp 1621261055
transform 1 0 2592 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_23
timestamp 1621261055
transform 1 0 3360 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_4
timestamp 1621261055
transform 1 0 1536 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_12
timestamp 1621261055
transform 1 0 2304 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_20
timestamp 1621261055
transform 1 0 3072 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_426
timestamp 1621261055
transform 1 0 3840 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_31
timestamp 1621261055
transform 1 0 4128 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_39
timestamp 1621261055
transform 1 0 4896 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_47
timestamp 1621261055
transform 1 0 5664 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_29
timestamp 1621261055
transform 1 0 3936 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_37
timestamp 1621261055
transform 1 0 4704 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_45
timestamp 1621261055
transform 1 0 5472 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_53
timestamp 1621261055
transform 1 0 6240 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_61
timestamp 1621261055
transform 1 0 7008 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_56
timestamp 1621261055
transform 1 0 6528 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_416
timestamp 1621261055
transform 1 0 6432 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_69
timestamp 1621261055
transform 1 0 7776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_64
timestamp 1621261055
transform 1 0 7296 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_70
timestamp 1621261055
transform 1 0 7488 0 1 17982
box -38 -49 230 715
use INVX4  INVX4
timestamp 1624893035
transform 1 0 7680 0 1 17982
box 0 -48 864 714
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_81
timestamp 1621261055
transform 1 0 8928 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_77
timestamp 1621261055
transform 1 0 8544 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_77
timestamp 1621261055
transform 1 0 8544 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_427
timestamp 1621261055
transform 1 0 9120 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_85
timestamp 1621261055
transform 1 0 9312 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_93
timestamp 1621261055
transform 1 0 10080 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_101
timestamp 1621261055
transform 1 0 10848 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_84
timestamp 1621261055
transform 1 0 9216 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_92
timestamp 1621261055
transform 1 0 9984 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_100
timestamp 1621261055
transform 1 0 10752 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_108
timestamp 1621261055
transform 1 0 11520 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_417
timestamp 1621261055
transform 1 0 11712 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_23_109
timestamp 1621261055
transform 1 0 11616 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_111
timestamp 1621261055
transform 1 0 11808 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_119
timestamp 1621261055
transform 1 0 12576 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_127
timestamp 1621261055
transform 1 0 13344 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_135
timestamp 1621261055
transform 1 0 14112 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_116
timestamp 1621261055
transform 1 0 12288 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_124
timestamp 1621261055
transform 1 0 13056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_132
timestamp 1621261055
transform 1 0 13824 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_428
timestamp 1621261055
transform 1 0 14400 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_143
timestamp 1621261055
transform 1 0 14880 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_151
timestamp 1621261055
transform 1 0 15648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_159
timestamp 1621261055
transform 1 0 16416 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_136
timestamp 1621261055
transform 1 0 14208 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_139
timestamp 1621261055
transform 1 0 14496 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_147
timestamp 1621261055
transform 1 0 15264 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_155
timestamp 1621261055
transform 1 0 16032 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_418
timestamp 1621261055
transform 1 0 16992 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_163
timestamp 1621261055
transform 1 0 16800 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_166
timestamp 1621261055
transform 1 0 17088 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_174
timestamp 1621261055
transform 1 0 17856 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_182
timestamp 1621261055
transform 1 0 18624 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_163
timestamp 1621261055
transform 1 0 16800 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_171
timestamp 1621261055
transform 1 0 17568 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_179
timestamp 1621261055
transform 1 0 18336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_187
timestamp 1621261055
transform 1 0 19104 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_194
timestamp 1621261055
transform 1 0 19776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_191
timestamp 1621261055
transform 1 0 19488 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_190
timestamp 1621261055
transform 1 0 19392 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_429
timestamp 1621261055
transform 1 0 19680 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_24_206
timestamp 1621261055
transform 1 0 20928 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_24_202
timestamp 1621261055
transform 1 0 20544 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_206
timestamp 1621261055
transform 1 0 20928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_198
timestamp 1621261055
transform 1 0 20160 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_210
timestamp 1621261055
transform 1 0 21312 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_214
timestamp 1621261055
transform 1 0 21696 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _084_
timestamp 1621261055
transform 1 0 21024 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_218
timestamp 1621261055
transform 1 0 22080 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_221
timestamp 1621261055
transform 1 0 22368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_218
timestamp 1621261055
transform 1 0 22080 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_419
timestamp 1621261055
transform 1 0 22272 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_226
timestamp 1621261055
transform 1 0 22848 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_229
timestamp 1621261055
transform 1 0 23136 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_242
timestamp 1621261055
transform 1 0 24384 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_234
timestamp 1621261055
transform 1 0 23616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_237
timestamp 1621261055
transform 1 0 23904 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _145_
timestamp 1621261055
transform 1 0 24288 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_249
timestamp 1621261055
transform 1 0 25056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_246
timestamp 1621261055
transform 1 0 24768 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_244
timestamp 1621261055
transform 1 0 24576 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_430
timestamp 1621261055
transform 1 0 24960 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_257
timestamp 1621261055
transform 1 0 25824 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_258
timestamp 1621261055
transform 1 0 25920 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_256
timestamp 1621261055
transform 1 0 25728 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_252
timestamp 1621261055
transform 1 0 25344 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_20
timestamp 1621261055
transform -1 0 26208 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_265
timestamp 1621261055
transform 1 0 26592 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_264
timestamp 1621261055
transform 1 0 26496 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _011_
timestamp 1621261055
transform -1 0 26496 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_273
timestamp 1621261055
transform 1 0 27360 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_276
timestamp 1621261055
transform 1 0 27648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_274
timestamp 1621261055
transform 1 0 27456 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_272
timestamp 1621261055
transform 1 0 27264 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_420
timestamp 1621261055
transform 1 0 27552 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_281
timestamp 1621261055
transform 1 0 28128 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_284
timestamp 1621261055
transform 1 0 28416 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_289
timestamp 1621261055
transform 1 0 28896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_292
timestamp 1621261055
transform 1 0 29184 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_297
timestamp 1621261055
transform 1 0 29664 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_431
timestamp 1621261055
transform 1 0 30240 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_300
timestamp 1621261055
transform 1 0 29952 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_308
timestamp 1621261055
transform 1 0 30720 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_316
timestamp 1621261055
transform 1 0 31488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_324
timestamp 1621261055
transform 1 0 32256 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_301
timestamp 1621261055
transform 1 0 30048 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_304
timestamp 1621261055
transform 1 0 30336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_312
timestamp 1621261055
transform 1 0 31104 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_320
timestamp 1621261055
transform 1 0 31872 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_421
timestamp 1621261055
transform 1 0 32832 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_328
timestamp 1621261055
transform 1 0 32640 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_331
timestamp 1621261055
transform 1 0 32928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_339
timestamp 1621261055
transform 1 0 33696 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_347
timestamp 1621261055
transform 1 0 34464 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_328
timestamp 1621261055
transform 1 0 32640 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_336
timestamp 1621261055
transform 1 0 33408 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_344
timestamp 1621261055
transform 1 0 34176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_432
timestamp 1621261055
transform 1 0 35520 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_355
timestamp 1621261055
transform 1 0 35232 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_363
timestamp 1621261055
transform 1 0 36000 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_371
timestamp 1621261055
transform 1 0 36768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_352
timestamp 1621261055
transform 1 0 34944 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_356
timestamp 1621261055
transform 1 0 35328 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_359
timestamp 1621261055
transform 1 0 35616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_367
timestamp 1621261055
transform 1 0 36384 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_375
timestamp 1621261055
transform 1 0 37152 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_422
timestamp 1621261055
transform 1 0 38112 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_23_379
timestamp 1621261055
transform 1 0 37536 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_383
timestamp 1621261055
transform 1 0 37920 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_386
timestamp 1621261055
transform 1 0 38208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_394
timestamp 1621261055
transform 1 0 38976 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_402
timestamp 1621261055
transform 1 0 39744 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_383
timestamp 1621261055
transform 1 0 37920 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_391
timestamp 1621261055
transform 1 0 38688 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_399
timestamp 1621261055
transform 1 0 39456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_411
timestamp 1621261055
transform 1 0 40608 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_407
timestamp 1621261055
transform 1 0 40224 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_413
timestamp 1621261055
transform 1 0 40800 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_433
timestamp 1621261055
transform 1 0 40800 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _154_
timestamp 1621261055
transform 1 0 40512 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_422
timestamp 1621261055
transform 1 0 41664 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_414
timestamp 1621261055
transform 1 0 40896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_421
timestamp 1621261055
transform 1 0 41568 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_430
timestamp 1621261055
transform 1 0 42432 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_429
timestamp 1621261055
transform 1 0 42336 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_423
timestamp 1621261055
transform 1 0 43392 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_437
timestamp 1621261055
transform 1 0 43104 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_23_439
timestamp 1621261055
transform 1 0 43296 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_441
timestamp 1621261055
transform 1 0 43488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_449
timestamp 1621261055
transform 1 0 44256 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_457
timestamp 1621261055
transform 1 0 45024 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_438
timestamp 1621261055
transform 1 0 43200 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_446
timestamp 1621261055
transform 1 0 43968 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_454
timestamp 1621261055
transform 1 0 44736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_434
timestamp 1621261055
transform 1 0 46080 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_465
timestamp 1621261055
transform 1 0 45792 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_473
timestamp 1621261055
transform 1 0 46560 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_481
timestamp 1621261055
transform 1 0 47328 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_462
timestamp 1621261055
transform 1 0 45504 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_466
timestamp 1621261055
transform 1 0 45888 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_24_469
timestamp 1621261055
transform 1 0 46176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_477
timestamp 1621261055
transform 1 0 46944 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_485
timestamp 1621261055
transform 1 0 47712 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_493
timestamp 1621261055
transform 1 0 48480 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_493
timestamp 1621261055
transform 1 0 48480 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_489
timestamp 1621261055
transform 1 0 48096 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_500
timestamp 1621261055
transform 1 0 49152 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_496
timestamp 1621261055
transform 1 0 48768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_14
timestamp 1621261055
transform 1 0 48672 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_424
timestamp 1621261055
transform 1 0 48672 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _007_
timestamp 1621261055
transform 1 0 48864 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_508
timestamp 1621261055
transform 1 0 49920 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_512
timestamp 1621261055
transform 1 0 50304 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_504
timestamp 1621261055
transform 1 0 49536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_520
timestamp 1621261055
transform 1 0 51072 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_516
timestamp 1621261055
transform 1 0 50688 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_23_518
timestamp 1621261055
transform 1 0 50880 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_516
timestamp 1621261055
transform 1 0 50688 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_91
timestamp 1621261055
transform -1 0 51168 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _038_
timestamp 1621261055
transform -1 0 51456 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_24_524
timestamp 1621261055
transform 1 0 51456 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_24_522
timestamp 1621261055
transform 1 0 51264 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_524
timestamp 1621261055
transform 1 0 51456 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_435
timestamp 1621261055
transform 1 0 51360 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _144_
timestamp 1621261055
transform 1 0 51840 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_539
timestamp 1621261055
transform 1 0 52896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_531
timestamp 1621261055
transform 1 0 52128 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_532
timestamp 1621261055
transform 1 0 52224 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_540
timestamp 1621261055
transform 1 0 52992 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_425
timestamp 1621261055
transform 1 0 53952 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_548
timestamp 1621261055
transform 1 0 53760 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_551
timestamp 1621261055
transform 1 0 54048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_559
timestamp 1621261055
transform 1 0 54816 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_567
timestamp 1621261055
transform 1 0 55584 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_547
timestamp 1621261055
transform 1 0 53664 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_555
timestamp 1621261055
transform 1 0 54432 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_563
timestamp 1621261055
transform 1 0 55200 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_436
timestamp 1621261055
transform 1 0 56640 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_575
timestamp 1621261055
transform 1 0 56352 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_583
timestamp 1621261055
transform 1 0 57120 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_591
timestamp 1621261055
transform 1 0 57888 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_24_571
timestamp 1621261055
transform 1 0 55968 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_575
timestamp 1621261055
transform 1 0 56352 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_24_577
timestamp 1621261055
transform 1 0 56544 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_579
timestamp 1621261055
transform 1 0 56736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_587
timestamp 1621261055
transform 1 0 57504 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_47
timestamp 1621261055
transform -1 0 58848 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_49
timestamp 1621261055
transform -1 0 58848 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_595
timestamp 1621261055
transform 1 0 58272 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_595
timestamp 1621261055
transform 1 0 58272 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_50
timestamp 1621261055
transform 1 0 1152 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_4
timestamp 1621261055
transform 1 0 1536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_12
timestamp 1621261055
transform 1 0 2304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_20
timestamp 1621261055
transform 1 0 3072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_28
timestamp 1621261055
transform 1 0 3840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_36
timestamp 1621261055
transform 1 0 4608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_44
timestamp 1621261055
transform 1 0 5376 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_52
timestamp 1621261055
transform 1 0 6144 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_54
timestamp 1621261055
transform 1 0 6336 0 1 19314
box -38 -49 134 715
use INVX8  INVX8
timestamp 1624893035
transform 1 0 7680 0 1 19314
box 0 -48 1440 714
use sky130_fd_sc_ls__conb_1  _160_
timestamp 1621261055
transform 1 0 6912 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_437
timestamp 1621261055
transform 1 0 6432 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_77
timestamp 1621261055
transform 1 0 7488 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_105
timestamp 1621261055
transform 1 0 6720 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_56
timestamp 1621261055
transform 1 0 6528 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_63
timestamp 1621261055
transform 1 0 7200 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_65
timestamp 1621261055
transform 1 0 7392 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_83
timestamp 1621261055
transform 1 0 9120 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_91
timestamp 1621261055
transform 1 0 9888 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_99
timestamp 1621261055
transform 1 0 10656 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_107
timestamp 1621261055
transform 1 0 11424 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_438
timestamp 1621261055
transform 1 0 11712 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_25_109
timestamp 1621261055
transform 1 0 11616 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_111
timestamp 1621261055
transform 1 0 11808 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_119
timestamp 1621261055
transform 1 0 12576 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_127
timestamp 1621261055
transform 1 0 13344 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_135
timestamp 1621261055
transform 1 0 14112 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_143
timestamp 1621261055
transform 1 0 14880 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_151
timestamp 1621261055
transform 1 0 15648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_159
timestamp 1621261055
transform 1 0 16416 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_439
timestamp 1621261055
transform 1 0 16992 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_163
timestamp 1621261055
transform 1 0 16800 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_166
timestamp 1621261055
transform 1 0 17088 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_174
timestamp 1621261055
transform 1 0 17856 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_182
timestamp 1621261055
transform 1 0 18624 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_190
timestamp 1621261055
transform 1 0 19392 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_198
timestamp 1621261055
transform 1 0 20160 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_206
timestamp 1621261055
transform 1 0 20928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_214
timestamp 1621261055
transform 1 0 21696 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_440
timestamp 1621261055
transform 1 0 22272 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_218
timestamp 1621261055
transform 1 0 22080 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_221
timestamp 1621261055
transform 1 0 22368 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_229
timestamp 1621261055
transform 1 0 23136 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_237
timestamp 1621261055
transform 1 0 23904 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_245
timestamp 1621261055
transform 1 0 24672 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_253
timestamp 1621261055
transform 1 0 25440 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_261
timestamp 1621261055
transform 1 0 26208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_269
timestamp 1621261055
transform 1 0 26976 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_441
timestamp 1621261055
transform 1 0 27552 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_273
timestamp 1621261055
transform 1 0 27360 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_276
timestamp 1621261055
transform 1 0 27648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_284
timestamp 1621261055
transform 1 0 28416 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_292
timestamp 1621261055
transform 1 0 29184 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_300
timestamp 1621261055
transform 1 0 29952 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_308
timestamp 1621261055
transform 1 0 30720 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_316
timestamp 1621261055
transform 1 0 31488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_324
timestamp 1621261055
transform 1 0 32256 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _184_
timestamp 1621261055
transform 1 0 34560 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_442
timestamp 1621261055
transform 1 0 32832 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_328
timestamp 1621261055
transform 1 0 32640 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_331
timestamp 1621261055
transform 1 0 32928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_339
timestamp 1621261055
transform 1 0 33696 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_25_347
timestamp 1621261055
transform 1 0 34464 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_351
timestamp 1621261055
transform 1 0 34848 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_359
timestamp 1621261055
transform 1 0 35616 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_367
timestamp 1621261055
transform 1 0 36384 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_375
timestamp 1621261055
transform 1 0 37152 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_443
timestamp 1621261055
transform 1 0 38112 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_383
timestamp 1621261055
transform 1 0 37920 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_386
timestamp 1621261055
transform 1 0 38208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_394
timestamp 1621261055
transform 1 0 38976 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_402
timestamp 1621261055
transform 1 0 39744 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_410
timestamp 1621261055
transform 1 0 40512 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_418
timestamp 1621261055
transform 1 0 41280 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_426
timestamp 1621261055
transform 1 0 42048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_444
timestamp 1621261055
transform 1 0 43392 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_434
timestamp 1621261055
transform 1 0 42816 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_438
timestamp 1621261055
transform 1 0 43200 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_441
timestamp 1621261055
transform 1 0 43488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_449
timestamp 1621261055
transform 1 0 44256 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_457
timestamp 1621261055
transform 1 0 45024 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_465
timestamp 1621261055
transform 1 0 45792 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_473
timestamp 1621261055
transform 1 0 46560 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_481
timestamp 1621261055
transform 1 0 47328 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_445
timestamp 1621261055
transform 1 0 48672 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_489
timestamp 1621261055
transform 1 0 48096 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_493
timestamp 1621261055
transform 1 0 48480 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_496
timestamp 1621261055
transform 1 0 48768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_504
timestamp 1621261055
transform 1 0 49536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_512
timestamp 1621261055
transform 1 0 50304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_520
timestamp 1621261055
transform 1 0 51072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_528
timestamp 1621261055
transform 1 0 51840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_536
timestamp 1621261055
transform 1 0 52608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_446
timestamp 1621261055
transform 1 0 53952 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_544
timestamp 1621261055
transform 1 0 53376 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_548
timestamp 1621261055
transform 1 0 53760 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_551
timestamp 1621261055
transform 1 0 54048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_559
timestamp 1621261055
transform 1 0 54816 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_567
timestamp 1621261055
transform 1 0 55584 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_575
timestamp 1621261055
transform 1 0 56352 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_583
timestamp 1621261055
transform 1 0 57120 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_591
timestamp 1621261055
transform 1 0 57888 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_51
timestamp 1621261055
transform -1 0 58848 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_595
timestamp 1621261055
transform 1 0 58272 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_52
timestamp 1621261055
transform 1 0 1152 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_26_4
timestamp 1621261055
transform 1 0 1536 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_12
timestamp 1621261055
transform 1 0 2304 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_20
timestamp 1621261055
transform 1 0 3072 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_447
timestamp 1621261055
transform 1 0 3840 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_29
timestamp 1621261055
transform 1 0 3936 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_37
timestamp 1621261055
transform 1 0 4704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_45
timestamp 1621261055
transform 1 0 5472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_53
timestamp 1621261055
transform 1 0 6240 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_61
timestamp 1621261055
transform 1 0 7008 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_69
timestamp 1621261055
transform 1 0 7776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_77
timestamp 1621261055
transform 1 0 8544 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_81
timestamp 1621261055
transform 1 0 8928 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_448
timestamp 1621261055
transform 1 0 9120 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_84
timestamp 1621261055
transform 1 0 9216 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_92
timestamp 1621261055
transform 1 0 9984 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_100
timestamp 1621261055
transform 1 0 10752 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_108
timestamp 1621261055
transform 1 0 11520 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_116
timestamp 1621261055
transform 1 0 12288 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_124
timestamp 1621261055
transform 1 0 13056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_132
timestamp 1621261055
transform 1 0 13824 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _126_
timestamp 1621261055
transform 1 0 15936 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_449
timestamp 1621261055
transform 1 0 14400 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_136
timestamp 1621261055
transform 1 0 14208 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_139
timestamp 1621261055
transform 1 0 14496 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_147
timestamp 1621261055
transform 1 0 15264 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_151
timestamp 1621261055
transform 1 0 15648 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_153
timestamp 1621261055
transform 1 0 15840 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_157
timestamp 1621261055
transform 1 0 16224 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_165
timestamp 1621261055
transform 1 0 16992 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_173
timestamp 1621261055
transform 1 0 17760 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_181
timestamp 1621261055
transform 1 0 18528 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_189
timestamp 1621261055
transform 1 0 19296 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_450
timestamp 1621261055
transform 1 0 19680 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_194
timestamp 1621261055
transform 1 0 19776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_202
timestamp 1621261055
transform 1 0 20544 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_210
timestamp 1621261055
transform 1 0 21312 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _052_
timestamp 1621261055
transform 1 0 24096 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_68
timestamp 1621261055
transform 1 0 23904 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_218
timestamp 1621261055
transform 1 0 22080 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_226
timestamp 1621261055
transform 1 0 22848 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_234
timestamp 1621261055
transform 1 0 23616 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_236
timestamp 1621261055
transform 1 0 23808 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_242
timestamp 1621261055
transform 1 0 24384 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_451
timestamp 1621261055
transform 1 0 24960 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_246
timestamp 1621261055
transform 1 0 24768 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_249
timestamp 1621261055
transform 1 0 25056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_257
timestamp 1621261055
transform 1 0 25824 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_265
timestamp 1621261055
transform 1 0 26592 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _108_
timestamp 1621261055
transform 1 0 27360 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_276
timestamp 1621261055
transform 1 0 27648 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_284
timestamp 1621261055
transform 1 0 28416 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_292
timestamp 1621261055
transform 1 0 29184 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_452
timestamp 1621261055
transform 1 0 30240 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_300
timestamp 1621261055
transform 1 0 29952 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_302
timestamp 1621261055
transform 1 0 30144 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_304
timestamp 1621261055
transform 1 0 30336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_312
timestamp 1621261055
transform 1 0 31104 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_320
timestamp 1621261055
transform 1 0 31872 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_328
timestamp 1621261055
transform 1 0 32640 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_336
timestamp 1621261055
transform 1 0 33408 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_344
timestamp 1621261055
transform 1 0 34176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_453
timestamp 1621261055
transform 1 0 35520 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_352
timestamp 1621261055
transform 1 0 34944 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_356
timestamp 1621261055
transform 1 0 35328 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_359
timestamp 1621261055
transform 1 0 35616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_367
timestamp 1621261055
transform 1 0 36384 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_375
timestamp 1621261055
transform 1 0 37152 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_383
timestamp 1621261055
transform 1 0 37920 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_391
timestamp 1621261055
transform 1 0 38688 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_399
timestamp 1621261055
transform 1 0 39456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_454
timestamp 1621261055
transform 1 0 40800 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_407
timestamp 1621261055
transform 1 0 40224 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_411
timestamp 1621261055
transform 1 0 40608 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_414
timestamp 1621261055
transform 1 0 40896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_422
timestamp 1621261055
transform 1 0 41664 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_430
timestamp 1621261055
transform 1 0 42432 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_438
timestamp 1621261055
transform 1 0 43200 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_446
timestamp 1621261055
transform 1 0 43968 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_454
timestamp 1621261055
transform 1 0 44736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_455
timestamp 1621261055
transform 1 0 46080 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_462
timestamp 1621261055
transform 1 0 45504 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_466
timestamp 1621261055
transform 1 0 45888 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_469
timestamp 1621261055
transform 1 0 46176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_477
timestamp 1621261055
transform 1 0 46944 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_485
timestamp 1621261055
transform 1 0 47712 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_493
timestamp 1621261055
transform 1 0 48480 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_501
timestamp 1621261055
transform 1 0 49248 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_509
timestamp 1621261055
transform 1 0 50016 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_456
timestamp 1621261055
transform 1 0 51360 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_517
timestamp 1621261055
transform 1 0 50784 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_521
timestamp 1621261055
transform 1 0 51168 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_524
timestamp 1621261055
transform 1 0 51456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_532
timestamp 1621261055
transform 1 0 52224 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_540
timestamp 1621261055
transform 1 0 52992 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_548
timestamp 1621261055
transform 1 0 53760 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_556
timestamp 1621261055
transform 1 0 54528 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_564
timestamp 1621261055
transform 1 0 55296 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_457
timestamp 1621261055
transform 1 0 56640 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_572
timestamp 1621261055
transform 1 0 56064 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_576
timestamp 1621261055
transform 1 0 56448 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_579
timestamp 1621261055
transform 1 0 56736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_587
timestamp 1621261055
transform 1 0 57504 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_53
timestamp 1621261055
transform -1 0 58848 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_595
timestamp 1621261055
transform 1 0 58272 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_54
timestamp 1621261055
transform 1 0 1152 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_4
timestamp 1621261055
transform 1 0 1536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_12
timestamp 1621261055
transform 1 0 2304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_20
timestamp 1621261055
transform 1 0 3072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_28
timestamp 1621261055
transform 1 0 3840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_36
timestamp 1621261055
transform 1 0 4608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_44
timestamp 1621261055
transform 1 0 5376 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_52
timestamp 1621261055
transform 1 0 6144 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_54
timestamp 1621261055
transform 1 0 6336 0 1 20646
box -38 -49 134 715
use MUX2X1  MUX2X1
timestamp 1624893035
transform 1 0 7680 0 1 20646
box 0 -48 1728 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_458
timestamp 1621261055
transform 1 0 6432 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_82
timestamp 1621261055
transform 1 0 7488 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_56
timestamp 1621261055
transform 1 0 6528 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_64
timestamp 1621261055
transform 1 0 7296 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_86
timestamp 1621261055
transform 1 0 9408 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_94
timestamp 1621261055
transform 1 0 10176 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_102
timestamp 1621261055
transform 1 0 10944 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_459
timestamp 1621261055
transform 1 0 11712 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_111
timestamp 1621261055
transform 1 0 11808 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_119
timestamp 1621261055
transform 1 0 12576 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_127
timestamp 1621261055
transform 1 0 13344 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_135
timestamp 1621261055
transform 1 0 14112 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_143
timestamp 1621261055
transform 1 0 14880 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_151
timestamp 1621261055
transform 1 0 15648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_159
timestamp 1621261055
transform 1 0 16416 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_460
timestamp 1621261055
transform 1 0 16992 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_163
timestamp 1621261055
transform 1 0 16800 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_166
timestamp 1621261055
transform 1 0 17088 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_174
timestamp 1621261055
transform 1 0 17856 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_182
timestamp 1621261055
transform 1 0 18624 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_190
timestamp 1621261055
transform 1 0 19392 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_198
timestamp 1621261055
transform 1 0 20160 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_206
timestamp 1621261055
transform 1 0 20928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_214
timestamp 1621261055
transform 1 0 21696 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_461
timestamp 1621261055
transform 1 0 22272 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_218
timestamp 1621261055
transform 1 0 22080 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_221
timestamp 1621261055
transform 1 0 22368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_229
timestamp 1621261055
transform 1 0 23136 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_237
timestamp 1621261055
transform 1 0 23904 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_245
timestamp 1621261055
transform 1 0 24672 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_253
timestamp 1621261055
transform 1 0 25440 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_261
timestamp 1621261055
transform 1 0 26208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_269
timestamp 1621261055
transform 1 0 26976 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_462
timestamp 1621261055
transform 1 0 27552 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_273
timestamp 1621261055
transform 1 0 27360 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_276
timestamp 1621261055
transform 1 0 27648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_284
timestamp 1621261055
transform 1 0 28416 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_292
timestamp 1621261055
transform 1 0 29184 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_300
timestamp 1621261055
transform 1 0 29952 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_308
timestamp 1621261055
transform 1 0 30720 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_316
timestamp 1621261055
transform 1 0 31488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_324
timestamp 1621261055
transform 1 0 32256 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_463
timestamp 1621261055
transform 1 0 32832 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_328
timestamp 1621261055
transform 1 0 32640 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_331
timestamp 1621261055
transform 1 0 32928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_339
timestamp 1621261055
transform 1 0 33696 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_347
timestamp 1621261055
transform 1 0 34464 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_355
timestamp 1621261055
transform 1 0 35232 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_363
timestamp 1621261055
transform 1 0 36000 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_371
timestamp 1621261055
transform 1 0 36768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_464
timestamp 1621261055
transform 1 0 38112 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_379
timestamp 1621261055
transform 1 0 37536 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_383
timestamp 1621261055
transform 1 0 37920 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_386
timestamp 1621261055
transform 1 0 38208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_394
timestamp 1621261055
transform 1 0 38976 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_402
timestamp 1621261055
transform 1 0 39744 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_410
timestamp 1621261055
transform 1 0 40512 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_418
timestamp 1621261055
transform 1 0 41280 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_426
timestamp 1621261055
transform 1 0 42048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_465
timestamp 1621261055
transform 1 0 43392 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_434
timestamp 1621261055
transform 1 0 42816 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_438
timestamp 1621261055
transform 1 0 43200 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_441
timestamp 1621261055
transform 1 0 43488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_449
timestamp 1621261055
transform 1 0 44256 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_457
timestamp 1621261055
transform 1 0 45024 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_465
timestamp 1621261055
transform 1 0 45792 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_473
timestamp 1621261055
transform 1 0 46560 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_481
timestamp 1621261055
transform 1 0 47328 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_466
timestamp 1621261055
transform 1 0 48672 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_489
timestamp 1621261055
transform 1 0 48096 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_493
timestamp 1621261055
transform 1 0 48480 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_496
timestamp 1621261055
transform 1 0 48768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_504
timestamp 1621261055
transform 1 0 49536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_512
timestamp 1621261055
transform 1 0 50304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_520
timestamp 1621261055
transform 1 0 51072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_528
timestamp 1621261055
transform 1 0 51840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_536
timestamp 1621261055
transform 1 0 52608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_467
timestamp 1621261055
transform 1 0 53952 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_544
timestamp 1621261055
transform 1 0 53376 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_548
timestamp 1621261055
transform 1 0 53760 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_551
timestamp 1621261055
transform 1 0 54048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_559
timestamp 1621261055
transform 1 0 54816 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_567
timestamp 1621261055
transform 1 0 55584 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_575
timestamp 1621261055
transform 1 0 56352 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_583
timestamp 1621261055
transform 1 0 57120 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_591
timestamp 1621261055
transform 1 0 57888 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_55
timestamp 1621261055
transform -1 0 58848 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_595
timestamp 1621261055
transform 1 0 58272 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_56
timestamp 1621261055
transform 1 0 1152 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_28_4
timestamp 1621261055
transform 1 0 1536 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_12
timestamp 1621261055
transform 1 0 2304 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_20
timestamp 1621261055
transform 1 0 3072 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_468
timestamp 1621261055
transform 1 0 3840 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_29
timestamp 1621261055
transform 1 0 3936 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_37
timestamp 1621261055
transform 1 0 4704 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_45
timestamp 1621261055
transform 1 0 5472 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_53
timestamp 1621261055
transform 1 0 6240 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _013_
timestamp 1621261055
transform -1 0 8352 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_24
timestamp 1621261055
transform -1 0 8064 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_61
timestamp 1621261055
transform 1 0 7008 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_28_69
timestamp 1621261055
transform 1 0 7776 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_75
timestamp 1621261055
transform 1 0 8352 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_469
timestamp 1621261055
transform 1 0 9120 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_84
timestamp 1621261055
transform 1 0 9216 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_92
timestamp 1621261055
transform 1 0 9984 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_100
timestamp 1621261055
transform 1 0 10752 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_108
timestamp 1621261055
transform 1 0 11520 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_116
timestamp 1621261055
transform 1 0 12288 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_124
timestamp 1621261055
transform 1 0 13056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_132
timestamp 1621261055
transform 1 0 13824 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_470
timestamp 1621261055
transform 1 0 14400 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_136
timestamp 1621261055
transform 1 0 14208 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_139
timestamp 1621261055
transform 1 0 14496 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_147
timestamp 1621261055
transform 1 0 15264 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_155
timestamp 1621261055
transform 1 0 16032 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_163
timestamp 1621261055
transform 1 0 16800 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_171
timestamp 1621261055
transform 1 0 17568 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_179
timestamp 1621261055
transform 1 0 18336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_187
timestamp 1621261055
transform 1 0 19104 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_471
timestamp 1621261055
transform 1 0 19680 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_191
timestamp 1621261055
transform 1 0 19488 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_194
timestamp 1621261055
transform 1 0 19776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_202
timestamp 1621261055
transform 1 0 20544 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_210
timestamp 1621261055
transform 1 0 21312 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_218
timestamp 1621261055
transform 1 0 22080 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_226
timestamp 1621261055
transform 1 0 22848 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_234
timestamp 1621261055
transform 1 0 23616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_242
timestamp 1621261055
transform 1 0 24384 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_472
timestamp 1621261055
transform 1 0 24960 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_246
timestamp 1621261055
transform 1 0 24768 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_249
timestamp 1621261055
transform 1 0 25056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_257
timestamp 1621261055
transform 1 0 25824 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_265
timestamp 1621261055
transform 1 0 26592 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_273
timestamp 1621261055
transform 1 0 27360 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_281
timestamp 1621261055
transform 1 0 28128 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_289
timestamp 1621261055
transform 1 0 28896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_297
timestamp 1621261055
transform 1 0 29664 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_473
timestamp 1621261055
transform 1 0 30240 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_301
timestamp 1621261055
transform 1 0 30048 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_304
timestamp 1621261055
transform 1 0 30336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_312
timestamp 1621261055
transform 1 0 31104 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_320
timestamp 1621261055
transform 1 0 31872 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _169_
timestamp 1621261055
transform 1 0 32640 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_28_331
timestamp 1621261055
transform 1 0 32928 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_339
timestamp 1621261055
transform 1 0 33696 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_347
timestamp 1621261055
transform 1 0 34464 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_474
timestamp 1621261055
transform 1 0 35520 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_355
timestamp 1621261055
transform 1 0 35232 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_28_357
timestamp 1621261055
transform 1 0 35424 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_359
timestamp 1621261055
transform 1 0 35616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_367
timestamp 1621261055
transform 1 0 36384 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_375
timestamp 1621261055
transform 1 0 37152 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_383
timestamp 1621261055
transform 1 0 37920 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_391
timestamp 1621261055
transform 1 0 38688 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_399
timestamp 1621261055
transform 1 0 39456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_475
timestamp 1621261055
transform 1 0 40800 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_407
timestamp 1621261055
transform 1 0 40224 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_411
timestamp 1621261055
transform 1 0 40608 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_414
timestamp 1621261055
transform 1 0 40896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_422
timestamp 1621261055
transform 1 0 41664 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_430
timestamp 1621261055
transform 1 0 42432 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_438
timestamp 1621261055
transform 1 0 43200 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_446
timestamp 1621261055
transform 1 0 43968 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_454
timestamp 1621261055
transform 1 0 44736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_476
timestamp 1621261055
transform 1 0 46080 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_462
timestamp 1621261055
transform 1 0 45504 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_466
timestamp 1621261055
transform 1 0 45888 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_469
timestamp 1621261055
transform 1 0 46176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_477
timestamp 1621261055
transform 1 0 46944 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_485
timestamp 1621261055
transform 1 0 47712 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_493
timestamp 1621261055
transform 1 0 48480 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_501
timestamp 1621261055
transform 1 0 49248 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_509
timestamp 1621261055
transform 1 0 50016 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_477
timestamp 1621261055
transform 1 0 51360 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_517
timestamp 1621261055
transform 1 0 50784 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_521
timestamp 1621261055
transform 1 0 51168 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_524
timestamp 1621261055
transform 1 0 51456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_532
timestamp 1621261055
transform 1 0 52224 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_540
timestamp 1621261055
transform 1 0 52992 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_548
timestamp 1621261055
transform 1 0 53760 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_556
timestamp 1621261055
transform 1 0 54528 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_564
timestamp 1621261055
transform 1 0 55296 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_478
timestamp 1621261055
transform 1 0 56640 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_572
timestamp 1621261055
transform 1 0 56064 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_576
timestamp 1621261055
transform 1 0 56448 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_579
timestamp 1621261055
transform 1 0 56736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_587
timestamp 1621261055
transform 1 0 57504 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_57
timestamp 1621261055
transform -1 0 58848 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_595
timestamp 1621261055
transform 1 0 58272 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_58
timestamp 1621261055
transform 1 0 1152 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_4
timestamp 1621261055
transform 1 0 1536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_12
timestamp 1621261055
transform 1 0 2304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_20
timestamp 1621261055
transform 1 0 3072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_28
timestamp 1621261055
transform 1 0 3840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_36
timestamp 1621261055
transform 1 0 4608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_44
timestamp 1621261055
transform 1 0 5376 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_52
timestamp 1621261055
transform 1 0 6144 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_54
timestamp 1621261055
transform 1 0 6336 0 1 21978
box -38 -49 134 715
use NAND2X1  NAND2X1
timestamp 1624893035
transform 1 0 7680 0 1 21978
box 0 -48 864 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_479
timestamp 1621261055
transform 1 0 6432 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_87
timestamp 1621261055
transform 1 0 7488 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_56
timestamp 1621261055
transform 1 0 6528 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_64
timestamp 1621261055
transform 1 0 7296 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_77
timestamp 1621261055
transform 1 0 8544 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_85
timestamp 1621261055
transform 1 0 9312 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_93
timestamp 1621261055
transform 1 0 10080 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_101
timestamp 1621261055
transform 1 0 10848 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_480
timestamp 1621261055
transform 1 0 11712 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_29_109
timestamp 1621261055
transform 1 0 11616 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_111
timestamp 1621261055
transform 1 0 11808 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_119
timestamp 1621261055
transform 1 0 12576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_127
timestamp 1621261055
transform 1 0 13344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_135
timestamp 1621261055
transform 1 0 14112 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_143
timestamp 1621261055
transform 1 0 14880 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_151
timestamp 1621261055
transform 1 0 15648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_159
timestamp 1621261055
transform 1 0 16416 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_481
timestamp 1621261055
transform 1 0 16992 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_163
timestamp 1621261055
transform 1 0 16800 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_166
timestamp 1621261055
transform 1 0 17088 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_174
timestamp 1621261055
transform 1 0 17856 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_182
timestamp 1621261055
transform 1 0 18624 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_190
timestamp 1621261055
transform 1 0 19392 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_198
timestamp 1621261055
transform 1 0 20160 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_206
timestamp 1621261055
transform 1 0 20928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_214
timestamp 1621261055
transform 1 0 21696 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_482
timestamp 1621261055
transform 1 0 22272 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_218
timestamp 1621261055
transform 1 0 22080 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_221
timestamp 1621261055
transform 1 0 22368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_229
timestamp 1621261055
transform 1 0 23136 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_237
timestamp 1621261055
transform 1 0 23904 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_245
timestamp 1621261055
transform 1 0 24672 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_253
timestamp 1621261055
transform 1 0 25440 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_261
timestamp 1621261055
transform 1 0 26208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_269
timestamp 1621261055
transform 1 0 26976 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_483
timestamp 1621261055
transform 1 0 27552 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_273
timestamp 1621261055
transform 1 0 27360 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_276
timestamp 1621261055
transform 1 0 27648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_284
timestamp 1621261055
transform 1 0 28416 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_292
timestamp 1621261055
transform 1 0 29184 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_300
timestamp 1621261055
transform 1 0 29952 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_308
timestamp 1621261055
transform 1 0 30720 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_316
timestamp 1621261055
transform 1 0 31488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_324
timestamp 1621261055
transform 1 0 32256 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_484
timestamp 1621261055
transform 1 0 32832 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_328
timestamp 1621261055
transform 1 0 32640 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_331
timestamp 1621261055
transform 1 0 32928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_339
timestamp 1621261055
transform 1 0 33696 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_347
timestamp 1621261055
transform 1 0 34464 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_355
timestamp 1621261055
transform 1 0 35232 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_363
timestamp 1621261055
transform 1 0 36000 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_371
timestamp 1621261055
transform 1 0 36768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_485
timestamp 1621261055
transform 1 0 38112 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_379
timestamp 1621261055
transform 1 0 37536 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_383
timestamp 1621261055
transform 1 0 37920 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_386
timestamp 1621261055
transform 1 0 38208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_394
timestamp 1621261055
transform 1 0 38976 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_402
timestamp 1621261055
transform 1 0 39744 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_410
timestamp 1621261055
transform 1 0 40512 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_418
timestamp 1621261055
transform 1 0 41280 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_426
timestamp 1621261055
transform 1 0 42048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_486
timestamp 1621261055
transform 1 0 43392 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_434
timestamp 1621261055
transform 1 0 42816 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_438
timestamp 1621261055
transform 1 0 43200 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_441
timestamp 1621261055
transform 1 0 43488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_449
timestamp 1621261055
transform 1 0 44256 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_457
timestamp 1621261055
transform 1 0 45024 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_465
timestamp 1621261055
transform 1 0 45792 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_473
timestamp 1621261055
transform 1 0 46560 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_481
timestamp 1621261055
transform 1 0 47328 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_487
timestamp 1621261055
transform 1 0 48672 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_489
timestamp 1621261055
transform 1 0 48096 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_493
timestamp 1621261055
transform 1 0 48480 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_496
timestamp 1621261055
transform 1 0 48768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_504
timestamp 1621261055
transform 1 0 49536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_512
timestamp 1621261055
transform 1 0 50304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_520
timestamp 1621261055
transform 1 0 51072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_528
timestamp 1621261055
transform 1 0 51840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_536
timestamp 1621261055
transform 1 0 52608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_488
timestamp 1621261055
transform 1 0 53952 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_544
timestamp 1621261055
transform 1 0 53376 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_548
timestamp 1621261055
transform 1 0 53760 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_551
timestamp 1621261055
transform 1 0 54048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_559
timestamp 1621261055
transform 1 0 54816 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_567
timestamp 1621261055
transform 1 0 55584 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_575
timestamp 1621261055
transform 1 0 56352 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_583
timestamp 1621261055
transform 1 0 57120 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_591
timestamp 1621261055
transform 1 0 57888 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_59
timestamp 1621261055
transform -1 0 58848 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_595
timestamp 1621261055
transform 1 0 58272 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_60
timestamp 1621261055
transform 1 0 1152 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_62
timestamp 1621261055
transform 1 0 1152 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_4
timestamp 1621261055
transform 1 0 1536 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_12
timestamp 1621261055
transform 1 0 2304 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_20
timestamp 1621261055
transform 1 0 3072 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_4
timestamp 1621261055
transform 1 0 1536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_12
timestamp 1621261055
transform 1 0 2304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_20
timestamp 1621261055
transform 1 0 3072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_28
timestamp 1621261055
transform 1 0 3840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_29
timestamp 1621261055
transform 1 0 3936 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_489
timestamp 1621261055
transform 1 0 3840 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_44
timestamp 1621261055
transform 1 0 5376 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_36
timestamp 1621261055
transform 1 0 4608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_37
timestamp 1621261055
transform 1 0 4704 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_52
timestamp 1621261055
transform 1 0 6144 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_53
timestamp 1621261055
transform 1 0 6240 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_45
timestamp 1621261055
transform 1 0 5472 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_54
timestamp 1621261055
transform 1 0 6336 0 1 23310
box -38 -49 134 715
use NAND3X1  NAND3X1
timestamp 1624893035
transform 1 0 7680 0 1 23310
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_500
timestamp 1621261055
transform 1 0 6432 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_61
timestamp 1621261055
transform 1 0 7008 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_69
timestamp 1621261055
transform 1 0 7776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_77
timestamp 1621261055
transform 1 0 8544 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_81
timestamp 1621261055
transform 1 0 8928 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_56
timestamp 1621261055
transform 1 0 6528 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_64
timestamp 1621261055
transform 1 0 7296 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_80
timestamp 1621261055
transform 1 0 8832 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _142_
timestamp 1621261055
transform 1 0 9984 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_490
timestamp 1621261055
transform 1 0 9120 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_84
timestamp 1621261055
transform 1 0 9216 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_95
timestamp 1621261055
transform 1 0 10272 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_103
timestamp 1621261055
transform 1 0 11040 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_88
timestamp 1621261055
transform 1 0 9600 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_96
timestamp 1621261055
transform 1 0 10368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_104
timestamp 1621261055
transform 1 0 11136 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_108
timestamp 1621261055
transform 1 0 11520 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_501
timestamp 1621261055
transform 1 0 11712 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_111
timestamp 1621261055
transform 1 0 11808 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_119
timestamp 1621261055
transform 1 0 12576 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_127
timestamp 1621261055
transform 1 0 13344 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_135
timestamp 1621261055
transform 1 0 14112 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_111
timestamp 1621261055
transform 1 0 11808 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_119
timestamp 1621261055
transform 1 0 12576 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_127
timestamp 1621261055
transform 1 0 13344 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_135
timestamp 1621261055
transform 1 0 14112 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_491
timestamp 1621261055
transform 1 0 14400 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_30_137
timestamp 1621261055
transform 1 0 14304 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_139
timestamp 1621261055
transform 1 0 14496 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_147
timestamp 1621261055
transform 1 0 15264 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_155
timestamp 1621261055
transform 1 0 16032 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_143
timestamp 1621261055
transform 1 0 14880 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_151
timestamp 1621261055
transform 1 0 15648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_159
timestamp 1621261055
transform 1 0 16416 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_502
timestamp 1621261055
transform 1 0 16992 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_163
timestamp 1621261055
transform 1 0 16800 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_171
timestamp 1621261055
transform 1 0 17568 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_179
timestamp 1621261055
transform 1 0 18336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_187
timestamp 1621261055
transform 1 0 19104 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_163
timestamp 1621261055
transform 1 0 16800 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_166
timestamp 1621261055
transform 1 0 17088 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_174
timestamp 1621261055
transform 1 0 17856 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_182
timestamp 1621261055
transform 1 0 18624 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_190
timestamp 1621261055
transform 1 0 19392 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_194
timestamp 1621261055
transform 1 0 19776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_191
timestamp 1621261055
transform 1 0 19488 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_55
timestamp 1621261055
transform 1 0 19776 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_492
timestamp 1621261055
transform 1 0 19680 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _049_
timestamp 1621261055
transform 1 0 19968 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_199
timestamp 1621261055
transform 1 0 20256 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_202
timestamp 1621261055
transform 1 0 20544 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_215
timestamp 1621261055
transform 1 0 21792 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_207
timestamp 1621261055
transform 1 0 21024 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_210
timestamp 1621261055
transform 1 0 21312 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_503
timestamp 1621261055
transform 1 0 22272 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_218
timestamp 1621261055
transform 1 0 22080 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_226
timestamp 1621261055
transform 1 0 22848 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_234
timestamp 1621261055
transform 1 0 23616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_242
timestamp 1621261055
transform 1 0 24384 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_31_219
timestamp 1621261055
transform 1 0 22176 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_221
timestamp 1621261055
transform 1 0 22368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_229
timestamp 1621261055
transform 1 0 23136 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_237
timestamp 1621261055
transform 1 0 23904 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_493
timestamp 1621261055
transform 1 0 24960 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_246
timestamp 1621261055
transform 1 0 24768 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_249
timestamp 1621261055
transform 1 0 25056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_257
timestamp 1621261055
transform 1 0 25824 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_265
timestamp 1621261055
transform 1 0 26592 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_245
timestamp 1621261055
transform 1 0 24672 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_253
timestamp 1621261055
transform 1 0 25440 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_261
timestamp 1621261055
transform 1 0 26208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_269
timestamp 1621261055
transform 1 0 26976 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_276
timestamp 1621261055
transform 1 0 27648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_273
timestamp 1621261055
transform 1 0 27360 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_273
timestamp 1621261055
transform 1 0 27360 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_504
timestamp 1621261055
transform 1 0 27552 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_284
timestamp 1621261055
transform 1 0 28416 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_281
timestamp 1621261055
transform 1 0 28128 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_296
timestamp 1621261055
transform 1 0 29568 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_292
timestamp 1621261055
transform 1 0 29184 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_289
timestamp 1621261055
transform 1 0 28896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_297
timestamp 1621261055
transform 1 0 29664 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _153_
timestamp 1621261055
transform 1 0 29760 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_494
timestamp 1621261055
transform 1 0 30240 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_301
timestamp 1621261055
transform 1 0 30048 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_304
timestamp 1621261055
transform 1 0 30336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_312
timestamp 1621261055
transform 1 0 31104 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_320
timestamp 1621261055
transform 1 0 31872 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_301
timestamp 1621261055
transform 1 0 30048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_309
timestamp 1621261055
transform 1 0 30816 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_317
timestamp 1621261055
transform 1 0 31584 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_505
timestamp 1621261055
transform 1 0 32832 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_328
timestamp 1621261055
transform 1 0 32640 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_336
timestamp 1621261055
transform 1 0 33408 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_344
timestamp 1621261055
transform 1 0 34176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_325
timestamp 1621261055
transform 1 0 32352 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_31_329
timestamp 1621261055
transform 1 0 32736 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_331
timestamp 1621261055
transform 1 0 32928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_339
timestamp 1621261055
transform 1 0 33696 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_347
timestamp 1621261055
transform 1 0 34464 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_355
timestamp 1621261055
transform 1 0 35232 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_359
timestamp 1621261055
transform 1 0 35616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_356
timestamp 1621261055
transform 1 0 35328 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_352
timestamp 1621261055
transform 1 0 34944 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_495
timestamp 1621261055
transform 1 0 35520 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_363
timestamp 1621261055
transform 1 0 36000 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_367
timestamp 1621261055
transform 1 0 36384 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_371
timestamp 1621261055
transform 1 0 36768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_375
timestamp 1621261055
transform 1 0 37152 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _085_
timestamp 1621261055
transform 1 0 37344 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_386
timestamp 1621261055
transform 1 0 38208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_383
timestamp 1621261055
transform 1 0 37920 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_379
timestamp 1621261055
transform 1 0 37536 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_380
timestamp 1621261055
transform 1 0 37632 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_506
timestamp 1621261055
transform 1 0 38112 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_394
timestamp 1621261055
transform 1 0 38976 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_388
timestamp 1621261055
transform 1 0 38400 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_402
timestamp 1621261055
transform 1 0 39744 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_404
timestamp 1621261055
transform 1 0 39936 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_396
timestamp 1621261055
transform 1 0 39168 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_410
timestamp 1621261055
transform 1 0 40512 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_412
timestamp 1621261055
transform 1 0 40704 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_496
timestamp 1621261055
transform 1 0 40800 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_31_420
timestamp 1621261055
transform 1 0 41472 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_418
timestamp 1621261055
transform 1 0 41280 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_422
timestamp 1621261055
transform 1 0 41664 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_414
timestamp 1621261055
transform 1 0 40896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _131_
timestamp 1621261055
transform 1 0 41568 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_424
timestamp 1621261055
transform 1 0 41856 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_430
timestamp 1621261055
transform 1 0 42432 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_432
timestamp 1621261055
transform 1 0 42624 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _098_
timestamp 1621261055
transform 1 0 44448 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_507
timestamp 1621261055
transform 1 0 43392 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_438
timestamp 1621261055
transform 1 0 43200 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_446
timestamp 1621261055
transform 1 0 43968 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_454
timestamp 1621261055
transform 1 0 44736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_441
timestamp 1621261055
transform 1 0 43488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_449
timestamp 1621261055
transform 1 0 44256 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_454
timestamp 1621261055
transform 1 0 44736 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_462
timestamp 1621261055
transform 1 0 45504 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_466
timestamp 1621261055
transform 1 0 45888 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_462
timestamp 1621261055
transform 1 0 45504 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_31_474
timestamp 1621261055
transform 1 0 46656 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_31_470
timestamp 1621261055
transform 1 0 46272 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_469
timestamp 1621261055
transform 1 0 46176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_497
timestamp 1621261055
transform 1 0 46080 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _168_
timestamp 1621261055
transform 1 0 46752 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_478
timestamp 1621261055
transform 1 0 47040 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_485
timestamp 1621261055
transform 1 0 47712 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_477
timestamp 1621261055
transform 1 0 46944 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_486
timestamp 1621261055
transform 1 0 47808 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_508
timestamp 1621261055
transform 1 0 48672 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_493
timestamp 1621261055
transform 1 0 48480 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_501
timestamp 1621261055
transform 1 0 49248 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_509
timestamp 1621261055
transform 1 0 50016 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_494
timestamp 1621261055
transform 1 0 48576 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_496
timestamp 1621261055
transform 1 0 48768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_504
timestamp 1621261055
transform 1 0 49536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_512
timestamp 1621261055
transform 1 0 50304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_498
timestamp 1621261055
transform 1 0 51360 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_517
timestamp 1621261055
transform 1 0 50784 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_521
timestamp 1621261055
transform 1 0 51168 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_524
timestamp 1621261055
transform 1 0 51456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_532
timestamp 1621261055
transform 1 0 52224 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_540
timestamp 1621261055
transform 1 0 52992 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_520
timestamp 1621261055
transform 1 0 51072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_528
timestamp 1621261055
transform 1 0 51840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_536
timestamp 1621261055
transform 1 0 52608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_509
timestamp 1621261055
transform 1 0 53952 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_548
timestamp 1621261055
transform 1 0 53760 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_556
timestamp 1621261055
transform 1 0 54528 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_564
timestamp 1621261055
transform 1 0 55296 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_544
timestamp 1621261055
transform 1 0 53376 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_548
timestamp 1621261055
transform 1 0 53760 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_551
timestamp 1621261055
transform 1 0 54048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_559
timestamp 1621261055
transform 1 0 54816 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_567
timestamp 1621261055
transform 1 0 55584 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_499
timestamp 1621261055
transform 1 0 56640 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_30_572
timestamp 1621261055
transform 1 0 56064 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_576
timestamp 1621261055
transform 1 0 56448 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_579
timestamp 1621261055
transform 1 0 56736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_587
timestamp 1621261055
transform 1 0 57504 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_575
timestamp 1621261055
transform 1 0 56352 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_583
timestamp 1621261055
transform 1 0 57120 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_591
timestamp 1621261055
transform 1 0 57888 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_61
timestamp 1621261055
transform -1 0 58848 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_63
timestamp 1621261055
transform -1 0 58848 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_595
timestamp 1621261055
transform 1 0 58272 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_595
timestamp 1621261055
transform 1 0 58272 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_64
timestamp 1621261055
transform 1 0 1152 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_4
timestamp 1621261055
transform 1 0 1536 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_12
timestamp 1621261055
transform 1 0 2304 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_20
timestamp 1621261055
transform 1 0 3072 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_510
timestamp 1621261055
transform 1 0 3840 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_29
timestamp 1621261055
transform 1 0 3936 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_37
timestamp 1621261055
transform 1 0 4704 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_45
timestamp 1621261055
transform 1 0 5472 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_53
timestamp 1621261055
transform 1 0 6240 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_61
timestamp 1621261055
transform 1 0 7008 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_69
timestamp 1621261055
transform 1 0 7776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_77
timestamp 1621261055
transform 1 0 8544 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_81
timestamp 1621261055
transform 1 0 8928 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _113_
timestamp 1621261055
transform 1 0 10272 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_511
timestamp 1621261055
transform 1 0 9120 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_84
timestamp 1621261055
transform 1 0 9216 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_92
timestamp 1621261055
transform 1 0 9984 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_32_94
timestamp 1621261055
transform 1 0 10176 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_98
timestamp 1621261055
transform 1 0 10560 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_106
timestamp 1621261055
transform 1 0 11328 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_114
timestamp 1621261055
transform 1 0 12096 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_122
timestamp 1621261055
transform 1 0 12864 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_130
timestamp 1621261055
transform 1 0 13632 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_512
timestamp 1621261055
transform 1 0 14400 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_139
timestamp 1621261055
transform 1 0 14496 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_147
timestamp 1621261055
transform 1 0 15264 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_155
timestamp 1621261055
transform 1 0 16032 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_163
timestamp 1621261055
transform 1 0 16800 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_171
timestamp 1621261055
transform 1 0 17568 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_179
timestamp 1621261055
transform 1 0 18336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_187
timestamp 1621261055
transform 1 0 19104 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_513
timestamp 1621261055
transform 1 0 19680 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_191
timestamp 1621261055
transform 1 0 19488 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_194
timestamp 1621261055
transform 1 0 19776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_202
timestamp 1621261055
transform 1 0 20544 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_210
timestamp 1621261055
transform 1 0 21312 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_218
timestamp 1621261055
transform 1 0 22080 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_226
timestamp 1621261055
transform 1 0 22848 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_234
timestamp 1621261055
transform 1 0 23616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_242
timestamp 1621261055
transform 1 0 24384 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_514
timestamp 1621261055
transform 1 0 24960 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_246
timestamp 1621261055
transform 1 0 24768 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_249
timestamp 1621261055
transform 1 0 25056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_257
timestamp 1621261055
transform 1 0 25824 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_265
timestamp 1621261055
transform 1 0 26592 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_273
timestamp 1621261055
transform 1 0 27360 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_281
timestamp 1621261055
transform 1 0 28128 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_289
timestamp 1621261055
transform 1 0 28896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_297
timestamp 1621261055
transform 1 0 29664 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_515
timestamp 1621261055
transform 1 0 30240 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_301
timestamp 1621261055
transform 1 0 30048 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_304
timestamp 1621261055
transform 1 0 30336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_312
timestamp 1621261055
transform 1 0 31104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_320
timestamp 1621261055
transform 1 0 31872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_328
timestamp 1621261055
transform 1 0 32640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_336
timestamp 1621261055
transform 1 0 33408 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_344
timestamp 1621261055
transform 1 0 34176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _086_
timestamp 1621261055
transform 1 0 36384 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_516
timestamp 1621261055
transform 1 0 35520 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_352
timestamp 1621261055
transform 1 0 34944 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_356
timestamp 1621261055
transform 1 0 35328 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_359
timestamp 1621261055
transform 1 0 35616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_370
timestamp 1621261055
transform 1 0 36672 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_378
timestamp 1621261055
transform 1 0 37440 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_386
timestamp 1621261055
transform 1 0 38208 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_394
timestamp 1621261055
transform 1 0 38976 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_402
timestamp 1621261055
transform 1 0 39744 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _136_
timestamp 1621261055
transform 1 0 41280 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_517
timestamp 1621261055
transform 1 0 40800 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_410
timestamp 1621261055
transform 1 0 40512 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_32_412
timestamp 1621261055
transform 1 0 40704 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_414
timestamp 1621261055
transform 1 0 40896 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_421
timestamp 1621261055
transform 1 0 41568 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_429
timestamp 1621261055
transform 1 0 42336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_437
timestamp 1621261055
transform 1 0 43104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_445
timestamp 1621261055
transform 1 0 43872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_453
timestamp 1621261055
transform 1 0 44640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_518
timestamp 1621261055
transform 1 0 46080 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_461
timestamp 1621261055
transform 1 0 45408 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_465
timestamp 1621261055
transform 1 0 45792 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_32_467
timestamp 1621261055
transform 1 0 45984 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_469
timestamp 1621261055
transform 1 0 46176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_477
timestamp 1621261055
transform 1 0 46944 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_485
timestamp 1621261055
transform 1 0 47712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_493
timestamp 1621261055
transform 1 0 48480 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_501
timestamp 1621261055
transform 1 0 49248 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_509
timestamp 1621261055
transform 1 0 50016 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_519
timestamp 1621261055
transform 1 0 51360 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_517
timestamp 1621261055
transform 1 0 50784 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_521
timestamp 1621261055
transform 1 0 51168 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_524
timestamp 1621261055
transform 1 0 51456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_532
timestamp 1621261055
transform 1 0 52224 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_540
timestamp 1621261055
transform 1 0 52992 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_548
timestamp 1621261055
transform 1 0 53760 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_556
timestamp 1621261055
transform 1 0 54528 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_564
timestamp 1621261055
transform 1 0 55296 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_520
timestamp 1621261055
transform 1 0 56640 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_32_572
timestamp 1621261055
transform 1 0 56064 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_576
timestamp 1621261055
transform 1 0 56448 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_579
timestamp 1621261055
transform 1 0 56736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_587
timestamp 1621261055
transform 1 0 57504 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_65
timestamp 1621261055
transform -1 0 58848 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_595
timestamp 1621261055
transform 1 0 58272 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_66
timestamp 1621261055
transform 1 0 1152 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_4
timestamp 1621261055
transform 1 0 1536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_12
timestamp 1621261055
transform 1 0 2304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_20
timestamp 1621261055
transform 1 0 3072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_28
timestamp 1621261055
transform 1 0 3840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_36
timestamp 1621261055
transform 1 0 4608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_44
timestamp 1621261055
transform 1 0 5376 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_52
timestamp 1621261055
transform 1 0 6144 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_54
timestamp 1621261055
transform 1 0 6336 0 1 24642
box -38 -49 134 715
use OR2X1  OR2X1
timestamp 1624893035
transform 1 0 7680 0 1 24642
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_521
timestamp 1621261055
transform 1 0 6432 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_56
timestamp 1621261055
transform 1 0 6528 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_64
timestamp 1621261055
transform 1 0 7296 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_80
timestamp 1621261055
transform 1 0 8832 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_88
timestamp 1621261055
transform 1 0 9600 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_96
timestamp 1621261055
transform 1 0 10368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_104
timestamp 1621261055
transform 1 0 11136 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_108
timestamp 1621261055
transform 1 0 11520 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_522
timestamp 1621261055
transform 1 0 11712 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_111
timestamp 1621261055
transform 1 0 11808 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_119
timestamp 1621261055
transform 1 0 12576 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_127
timestamp 1621261055
transform 1 0 13344 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_135
timestamp 1621261055
transform 1 0 14112 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_143
timestamp 1621261055
transform 1 0 14880 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_151
timestamp 1621261055
transform 1 0 15648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_159
timestamp 1621261055
transform 1 0 16416 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_523
timestamp 1621261055
transform 1 0 16992 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_163
timestamp 1621261055
transform 1 0 16800 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_166
timestamp 1621261055
transform 1 0 17088 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_174
timestamp 1621261055
transform 1 0 17856 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_182
timestamp 1621261055
transform 1 0 18624 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_190
timestamp 1621261055
transform 1 0 19392 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_198
timestamp 1621261055
transform 1 0 20160 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_206
timestamp 1621261055
transform 1 0 20928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_214
timestamp 1621261055
transform 1 0 21696 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_524
timestamp 1621261055
transform 1 0 22272 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_218
timestamp 1621261055
transform 1 0 22080 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_221
timestamp 1621261055
transform 1 0 22368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_229
timestamp 1621261055
transform 1 0 23136 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_237
timestamp 1621261055
transform 1 0 23904 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _165_
timestamp 1621261055
transform 1 0 26592 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_33_245
timestamp 1621261055
transform 1 0 24672 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_253
timestamp 1621261055
transform 1 0 25440 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_261
timestamp 1621261055
transform 1 0 26208 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_33_268
timestamp 1621261055
transform 1 0 26880 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_525
timestamp 1621261055
transform 1 0 27552 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_272
timestamp 1621261055
transform 1 0 27264 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_274
timestamp 1621261055
transform 1 0 27456 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_276
timestamp 1621261055
transform 1 0 27648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_284
timestamp 1621261055
transform 1 0 28416 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_292
timestamp 1621261055
transform 1 0 29184 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_300
timestamp 1621261055
transform 1 0 29952 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_308
timestamp 1621261055
transform 1 0 30720 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_316
timestamp 1621261055
transform 1 0 31488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_324
timestamp 1621261055
transform 1 0 32256 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _102_
timestamp 1621261055
transform 1 0 33312 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_526
timestamp 1621261055
transform 1 0 32832 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_328
timestamp 1621261055
transform 1 0 32640 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_33_331
timestamp 1621261055
transform 1 0 32928 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_338
timestamp 1621261055
transform 1 0 33600 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_346
timestamp 1621261055
transform 1 0 34368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_354
timestamp 1621261055
transform 1 0 35136 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_362
timestamp 1621261055
transform 1 0 35904 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_370
timestamp 1621261055
transform 1 0 36672 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_378
timestamp 1621261055
transform 1 0 37440 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_527
timestamp 1621261055
transform 1 0 38112 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_382
timestamp 1621261055
transform 1 0 37824 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_384
timestamp 1621261055
transform 1 0 38016 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_386
timestamp 1621261055
transform 1 0 38208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_394
timestamp 1621261055
transform 1 0 38976 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_402
timestamp 1621261055
transform 1 0 39744 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_410
timestamp 1621261055
transform 1 0 40512 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_418
timestamp 1621261055
transform 1 0 41280 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_426
timestamp 1621261055
transform 1 0 42048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_528
timestamp 1621261055
transform 1 0 43392 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_434
timestamp 1621261055
transform 1 0 42816 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_438
timestamp 1621261055
transform 1 0 43200 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_441
timestamp 1621261055
transform 1 0 43488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_449
timestamp 1621261055
transform 1 0 44256 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_457
timestamp 1621261055
transform 1 0 45024 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_465
timestamp 1621261055
transform 1 0 45792 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_473
timestamp 1621261055
transform 1 0 46560 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_481
timestamp 1621261055
transform 1 0 47328 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_529
timestamp 1621261055
transform 1 0 48672 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_489
timestamp 1621261055
transform 1 0 48096 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_493
timestamp 1621261055
transform 1 0 48480 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_496
timestamp 1621261055
transform 1 0 48768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_504
timestamp 1621261055
transform 1 0 49536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_512
timestamp 1621261055
transform 1 0 50304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _190_
timestamp 1621261055
transform 1 0 51072 0 1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_33_523
timestamp 1621261055
transform 1 0 51360 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_531
timestamp 1621261055
transform 1 0 52128 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_539
timestamp 1621261055
transform 1 0 52896 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_530
timestamp 1621261055
transform 1 0 53952 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_547
timestamp 1621261055
transform 1 0 53664 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_549
timestamp 1621261055
transform 1 0 53856 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_551
timestamp 1621261055
transform 1 0 54048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_559
timestamp 1621261055
transform 1 0 54816 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_567
timestamp 1621261055
transform 1 0 55584 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_575
timestamp 1621261055
transform 1 0 56352 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_583
timestamp 1621261055
transform 1 0 57120 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_591
timestamp 1621261055
transform 1 0 57888 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_67
timestamp 1621261055
transform -1 0 58848 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_595
timestamp 1621261055
transform 1 0 58272 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_68
timestamp 1621261055
transform 1 0 1152 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_4
timestamp 1621261055
transform 1 0 1536 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_12
timestamp 1621261055
transform 1 0 2304 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_20
timestamp 1621261055
transform 1 0 3072 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_531
timestamp 1621261055
transform 1 0 3840 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_29
timestamp 1621261055
transform 1 0 3936 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_37
timestamp 1621261055
transform 1 0 4704 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_45
timestamp 1621261055
transform 1 0 5472 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_53
timestamp 1621261055
transform 1 0 6240 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_61
timestamp 1621261055
transform 1 0 7008 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_69
timestamp 1621261055
transform 1 0 7776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_77
timestamp 1621261055
transform 1 0 8544 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_81
timestamp 1621261055
transform 1 0 8928 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_532
timestamp 1621261055
transform 1 0 9120 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_84
timestamp 1621261055
transform 1 0 9216 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_92
timestamp 1621261055
transform 1 0 9984 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_100
timestamp 1621261055
transform 1 0 10752 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_108
timestamp 1621261055
transform 1 0 11520 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_116
timestamp 1621261055
transform 1 0 12288 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_124
timestamp 1621261055
transform 1 0 13056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_132
timestamp 1621261055
transform 1 0 13824 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_533
timestamp 1621261055
transform 1 0 14400 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_136
timestamp 1621261055
transform 1 0 14208 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_139
timestamp 1621261055
transform 1 0 14496 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_147
timestamp 1621261055
transform 1 0 15264 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_155
timestamp 1621261055
transform 1 0 16032 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_163
timestamp 1621261055
transform 1 0 16800 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_171
timestamp 1621261055
transform 1 0 17568 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_179
timestamp 1621261055
transform 1 0 18336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_187
timestamp 1621261055
transform 1 0 19104 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_534
timestamp 1621261055
transform 1 0 19680 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_191
timestamp 1621261055
transform 1 0 19488 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_194
timestamp 1621261055
transform 1 0 19776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_202
timestamp 1621261055
transform 1 0 20544 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_210
timestamp 1621261055
transform 1 0 21312 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_218
timestamp 1621261055
transform 1 0 22080 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_226
timestamp 1621261055
transform 1 0 22848 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_234
timestamp 1621261055
transform 1 0 23616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_242
timestamp 1621261055
transform 1 0 24384 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _006_
timestamp 1621261055
transform -1 0 25728 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_535
timestamp 1621261055
transform 1 0 24960 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_10
timestamp 1621261055
transform -1 0 25440 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_246
timestamp 1621261055
transform 1 0 24768 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_249
timestamp 1621261055
transform 1 0 25056 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_256
timestamp 1621261055
transform 1 0 25728 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_264
timestamp 1621261055
transform 1 0 26496 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_272
timestamp 1621261055
transform 1 0 27264 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_280
timestamp 1621261055
transform 1 0 28032 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_288
timestamp 1621261055
transform 1 0 28800 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_296
timestamp 1621261055
transform 1 0 29568 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_536
timestamp 1621261055
transform 1 0 30240 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_300
timestamp 1621261055
transform 1 0 29952 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_34_302
timestamp 1621261055
transform 1 0 30144 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_304
timestamp 1621261055
transform 1 0 30336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_312
timestamp 1621261055
transform 1 0 31104 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_320
timestamp 1621261055
transform 1 0 31872 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _204_
timestamp 1621261055
transform 1 0 33312 0 -1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_34_328
timestamp 1621261055
transform 1 0 32640 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_332
timestamp 1621261055
transform 1 0 33024 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_34_334
timestamp 1621261055
transform 1 0 33216 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_338
timestamp 1621261055
transform 1 0 33600 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_346
timestamp 1621261055
transform 1 0 34368 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_537
timestamp 1621261055
transform 1 0 35520 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_354
timestamp 1621261055
transform 1 0 35136 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_34_359
timestamp 1621261055
transform 1 0 35616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_367
timestamp 1621261055
transform 1 0 36384 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_375
timestamp 1621261055
transform 1 0 37152 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_383
timestamp 1621261055
transform 1 0 37920 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_391
timestamp 1621261055
transform 1 0 38688 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_399
timestamp 1621261055
transform 1 0 39456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_538
timestamp 1621261055
transform 1 0 40800 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_407
timestamp 1621261055
transform 1 0 40224 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_411
timestamp 1621261055
transform 1 0 40608 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_414
timestamp 1621261055
transform 1 0 40896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_422
timestamp 1621261055
transform 1 0 41664 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_430
timestamp 1621261055
transform 1 0 42432 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_438
timestamp 1621261055
transform 1 0 43200 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_446
timestamp 1621261055
transform 1 0 43968 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_454
timestamp 1621261055
transform 1 0 44736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_539
timestamp 1621261055
transform 1 0 46080 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_462
timestamp 1621261055
transform 1 0 45504 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_466
timestamp 1621261055
transform 1 0 45888 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_469
timestamp 1621261055
transform 1 0 46176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_477
timestamp 1621261055
transform 1 0 46944 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_485
timestamp 1621261055
transform 1 0 47712 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_493
timestamp 1621261055
transform 1 0 48480 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_501
timestamp 1621261055
transform 1 0 49248 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_509
timestamp 1621261055
transform 1 0 50016 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_540
timestamp 1621261055
transform 1 0 51360 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_517
timestamp 1621261055
transform 1 0 50784 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_521
timestamp 1621261055
transform 1 0 51168 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_524
timestamp 1621261055
transform 1 0 51456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_532
timestamp 1621261055
transform 1 0 52224 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_540
timestamp 1621261055
transform 1 0 52992 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_548
timestamp 1621261055
transform 1 0 53760 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_556
timestamp 1621261055
transform 1 0 54528 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_564
timestamp 1621261055
transform 1 0 55296 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_541
timestamp 1621261055
transform 1 0 56640 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_34_572
timestamp 1621261055
transform 1 0 56064 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_576
timestamp 1621261055
transform 1 0 56448 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_579
timestamp 1621261055
transform 1 0 56736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_587
timestamp 1621261055
transform 1 0 57504 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_69
timestamp 1621261055
transform -1 0 58848 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_595
timestamp 1621261055
transform 1 0 58272 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _109_
timestamp 1621261055
transform 1 0 1728 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_70
timestamp 1621261055
transform 1 0 1152 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_4
timestamp 1621261055
transform 1 0 1536 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_9
timestamp 1621261055
transform 1 0 2016 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_17
timestamp 1621261055
transform 1 0 2784 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_25
timestamp 1621261055
transform 1 0 3552 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_33
timestamp 1621261055
transform 1 0 4320 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_41
timestamp 1621261055
transform 1 0 5088 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_49
timestamp 1621261055
transform 1 0 5856 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_53
timestamp 1621261055
transform 1 0 6240 0 1 25974
box -38 -49 230 715
use OR2X2  OR2X2
timestamp 1624893035
transform 1 0 7680 0 1 25974
box 0 -48 1152 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_542
timestamp 1621261055
transform 1 0 6432 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_56
timestamp 1621261055
transform 1 0 6528 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_64
timestamp 1621261055
transform 1 0 7296 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_80
timestamp 1621261055
transform 1 0 8832 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_88
timestamp 1621261055
transform 1 0 9600 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_96
timestamp 1621261055
transform 1 0 10368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_104
timestamp 1621261055
transform 1 0 11136 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_108
timestamp 1621261055
transform 1 0 11520 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_543
timestamp 1621261055
transform 1 0 11712 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_111
timestamp 1621261055
transform 1 0 11808 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_119
timestamp 1621261055
transform 1 0 12576 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_127
timestamp 1621261055
transform 1 0 13344 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_135
timestamp 1621261055
transform 1 0 14112 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_143
timestamp 1621261055
transform 1 0 14880 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_151
timestamp 1621261055
transform 1 0 15648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_159
timestamp 1621261055
transform 1 0 16416 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_544
timestamp 1621261055
transform 1 0 16992 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_163
timestamp 1621261055
transform 1 0 16800 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_166
timestamp 1621261055
transform 1 0 17088 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_174
timestamp 1621261055
transform 1 0 17856 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_182
timestamp 1621261055
transform 1 0 18624 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_190
timestamp 1621261055
transform 1 0 19392 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_198
timestamp 1621261055
transform 1 0 20160 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_206
timestamp 1621261055
transform 1 0 20928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_214
timestamp 1621261055
transform 1 0 21696 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_545
timestamp 1621261055
transform 1 0 22272 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_218
timestamp 1621261055
transform 1 0 22080 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_221
timestamp 1621261055
transform 1 0 22368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_229
timestamp 1621261055
transform 1 0 23136 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_237
timestamp 1621261055
transform 1 0 23904 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_245
timestamp 1621261055
transform 1 0 24672 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_253
timestamp 1621261055
transform 1 0 25440 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_261
timestamp 1621261055
transform 1 0 26208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_269
timestamp 1621261055
transform 1 0 26976 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_546
timestamp 1621261055
transform 1 0 27552 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_273
timestamp 1621261055
transform 1 0 27360 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_276
timestamp 1621261055
transform 1 0 27648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_284
timestamp 1621261055
transform 1 0 28416 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_292
timestamp 1621261055
transform 1 0 29184 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_300
timestamp 1621261055
transform 1 0 29952 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_308
timestamp 1621261055
transform 1 0 30720 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_316
timestamp 1621261055
transform 1 0 31488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_324
timestamp 1621261055
transform 1 0 32256 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_547
timestamp 1621261055
transform 1 0 32832 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_328
timestamp 1621261055
transform 1 0 32640 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_331
timestamp 1621261055
transform 1 0 32928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_339
timestamp 1621261055
transform 1 0 33696 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_347
timestamp 1621261055
transform 1 0 34464 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_355
timestamp 1621261055
transform 1 0 35232 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_363
timestamp 1621261055
transform 1 0 36000 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_371
timestamp 1621261055
transform 1 0 36768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_548
timestamp 1621261055
transform 1 0 38112 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_379
timestamp 1621261055
transform 1 0 37536 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_383
timestamp 1621261055
transform 1 0 37920 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_386
timestamp 1621261055
transform 1 0 38208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_394
timestamp 1621261055
transform 1 0 38976 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_402
timestamp 1621261055
transform 1 0 39744 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_410
timestamp 1621261055
transform 1 0 40512 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_418
timestamp 1621261055
transform 1 0 41280 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_426
timestamp 1621261055
transform 1 0 42048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_549
timestamp 1621261055
transform 1 0 43392 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_434
timestamp 1621261055
transform 1 0 42816 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_438
timestamp 1621261055
transform 1 0 43200 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_441
timestamp 1621261055
transform 1 0 43488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_449
timestamp 1621261055
transform 1 0 44256 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_457
timestamp 1621261055
transform 1 0 45024 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_465
timestamp 1621261055
transform 1 0 45792 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_473
timestamp 1621261055
transform 1 0 46560 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_481
timestamp 1621261055
transform 1 0 47328 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_550
timestamp 1621261055
transform 1 0 48672 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_489
timestamp 1621261055
transform 1 0 48096 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_493
timestamp 1621261055
transform 1 0 48480 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_496
timestamp 1621261055
transform 1 0 48768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_504
timestamp 1621261055
transform 1 0 49536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_512
timestamp 1621261055
transform 1 0 50304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_520
timestamp 1621261055
transform 1 0 51072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_528
timestamp 1621261055
transform 1 0 51840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_536
timestamp 1621261055
transform 1 0 52608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_551
timestamp 1621261055
transform 1 0 53952 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_544
timestamp 1621261055
transform 1 0 53376 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_548
timestamp 1621261055
transform 1 0 53760 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_551
timestamp 1621261055
transform 1 0 54048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_559
timestamp 1621261055
transform 1 0 54816 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_567
timestamp 1621261055
transform 1 0 55584 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _050_
timestamp 1621261055
transform -1 0 58080 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_59
timestamp 1621261055
transform -1 0 57792 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_575
timestamp 1621261055
transform 1 0 56352 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_583
timestamp 1621261055
transform 1 0 57120 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_35_587
timestamp 1621261055
transform 1 0 57504 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_593
timestamp 1621261055
transform 1 0 58080 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_71
timestamp 1621261055
transform -1 0 58848 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_72
timestamp 1621261055
transform 1 0 1152 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_4
timestamp 1621261055
transform 1 0 1536 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_12
timestamp 1621261055
transform 1 0 2304 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_20
timestamp 1621261055
transform 1 0 3072 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_552
timestamp 1621261055
transform 1 0 3840 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_29
timestamp 1621261055
transform 1 0 3936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_37
timestamp 1621261055
transform 1 0 4704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_45
timestamp 1621261055
transform 1 0 5472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_53
timestamp 1621261055
transform 1 0 6240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_61
timestamp 1621261055
transform 1 0 7008 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_69
timestamp 1621261055
transform 1 0 7776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_77
timestamp 1621261055
transform 1 0 8544 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_81
timestamp 1621261055
transform 1 0 8928 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_553
timestamp 1621261055
transform 1 0 9120 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_84
timestamp 1621261055
transform 1 0 9216 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_92
timestamp 1621261055
transform 1 0 9984 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_100
timestamp 1621261055
transform 1 0 10752 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_108
timestamp 1621261055
transform 1 0 11520 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_116
timestamp 1621261055
transform 1 0 12288 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_124
timestamp 1621261055
transform 1 0 13056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_132
timestamp 1621261055
transform 1 0 13824 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _087_
timestamp 1621261055
transform 1 0 14880 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_554
timestamp 1621261055
transform 1 0 14400 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_136
timestamp 1621261055
transform 1 0 14208 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_36_139
timestamp 1621261055
transform 1 0 14496 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_146
timestamp 1621261055
transform 1 0 15168 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_154
timestamp 1621261055
transform 1 0 15936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_162
timestamp 1621261055
transform 1 0 16704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_170
timestamp 1621261055
transform 1 0 17472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_178
timestamp 1621261055
transform 1 0 18240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_186
timestamp 1621261055
transform 1 0 19008 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_555
timestamp 1621261055
transform 1 0 19680 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_190
timestamp 1621261055
transform 1 0 19392 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_36_192
timestamp 1621261055
transform 1 0 19584 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_194
timestamp 1621261055
transform 1 0 19776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_202
timestamp 1621261055
transform 1 0 20544 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_210
timestamp 1621261055
transform 1 0 21312 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_218
timestamp 1621261055
transform 1 0 22080 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_226
timestamp 1621261055
transform 1 0 22848 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_234
timestamp 1621261055
transform 1 0 23616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_242
timestamp 1621261055
transform 1 0 24384 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_556
timestamp 1621261055
transform 1 0 24960 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_246
timestamp 1621261055
transform 1 0 24768 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_249
timestamp 1621261055
transform 1 0 25056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_257
timestamp 1621261055
transform 1 0 25824 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_265
timestamp 1621261055
transform 1 0 26592 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_273
timestamp 1621261055
transform 1 0 27360 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_281
timestamp 1621261055
transform 1 0 28128 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_289
timestamp 1621261055
transform 1 0 28896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_297
timestamp 1621261055
transform 1 0 29664 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_557
timestamp 1621261055
transform 1 0 30240 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_301
timestamp 1621261055
transform 1 0 30048 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_304
timestamp 1621261055
transform 1 0 30336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_312
timestamp 1621261055
transform 1 0 31104 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_320
timestamp 1621261055
transform 1 0 31872 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_328
timestamp 1621261055
transform 1 0 32640 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_336
timestamp 1621261055
transform 1 0 33408 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_344
timestamp 1621261055
transform 1 0 34176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _094_
timestamp 1621261055
transform 1 0 36000 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_558
timestamp 1621261055
transform 1 0 35520 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_352
timestamp 1621261055
transform 1 0 34944 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_356
timestamp 1621261055
transform 1 0 35328 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_36_359
timestamp 1621261055
transform 1 0 35616 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_366
timestamp 1621261055
transform 1 0 36288 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_374
timestamp 1621261055
transform 1 0 37056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _048_
timestamp 1621261055
transform -1 0 39072 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_49
timestamp 1621261055
transform -1 0 38784 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_382
timestamp 1621261055
transform 1 0 37824 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_395
timestamp 1621261055
transform 1 0 39072 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_403
timestamp 1621261055
transform 1 0 39840 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _065_
timestamp 1621261055
transform 1 0 42048 0 -1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_559
timestamp 1621261055
transform 1 0 40800 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_411
timestamp 1621261055
transform 1 0 40608 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_414
timestamp 1621261055
transform 1 0 40896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_422
timestamp 1621261055
transform 1 0 41664 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_36_429
timestamp 1621261055
transform 1 0 42336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_437
timestamp 1621261055
transform 1 0 43104 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_445
timestamp 1621261055
transform 1 0 43872 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_453
timestamp 1621261055
transform 1 0 44640 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_560
timestamp 1621261055
transform 1 0 46080 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_461
timestamp 1621261055
transform 1 0 45408 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_465
timestamp 1621261055
transform 1 0 45792 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_36_467
timestamp 1621261055
transform 1 0 45984 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_469
timestamp 1621261055
transform 1 0 46176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_477
timestamp 1621261055
transform 1 0 46944 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_485
timestamp 1621261055
transform 1 0 47712 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_493
timestamp 1621261055
transform 1 0 48480 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_501
timestamp 1621261055
transform 1 0 49248 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_509
timestamp 1621261055
transform 1 0 50016 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_561
timestamp 1621261055
transform 1 0 51360 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_517
timestamp 1621261055
transform 1 0 50784 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_521
timestamp 1621261055
transform 1 0 51168 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_524
timestamp 1621261055
transform 1 0 51456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_532
timestamp 1621261055
transform 1 0 52224 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_540
timestamp 1621261055
transform 1 0 52992 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_548
timestamp 1621261055
transform 1 0 53760 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_556
timestamp 1621261055
transform 1 0 54528 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_564
timestamp 1621261055
transform 1 0 55296 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_562
timestamp 1621261055
transform 1 0 56640 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_36_572
timestamp 1621261055
transform 1 0 56064 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_576
timestamp 1621261055
transform 1 0 56448 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_579
timestamp 1621261055
transform 1 0 56736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_587
timestamp 1621261055
transform 1 0 57504 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_73
timestamp 1621261055
transform -1 0 58848 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_595
timestamp 1621261055
transform 1 0 58272 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_74
timestamp 1621261055
transform 1 0 1152 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_4
timestamp 1621261055
transform 1 0 1536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_12
timestamp 1621261055
transform 1 0 2304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_20
timestamp 1621261055
transform 1 0 3072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _210_
timestamp 1621261055
transform 1 0 5088 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_37_28
timestamp 1621261055
transform 1 0 3840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_36
timestamp 1621261055
transform 1 0 4608 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_37_40
timestamp 1621261055
transform 1 0 4992 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_44
timestamp 1621261055
transform 1 0 5376 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_52
timestamp 1621261055
transform 1 0 6144 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_54
timestamp 1621261055
transform 1 0 6336 0 1 27306
box -38 -49 134 715
use XNOR2X1  XNOR2X1
timestamp 1624893035
transform 1 0 7680 0 1 27306
box 0 -48 2016 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_563
timestamp 1621261055
transform 1 0 6432 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_56
timestamp 1621261055
transform 1 0 6528 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_64
timestamp 1621261055
transform 1 0 7296 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_89
timestamp 1621261055
transform 1 0 9696 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_97
timestamp 1621261055
transform 1 0 10464 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_105
timestamp 1621261055
transform 1 0 11232 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_564
timestamp 1621261055
transform 1 0 11712 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_37_109
timestamp 1621261055
transform 1 0 11616 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_111
timestamp 1621261055
transform 1 0 11808 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_119
timestamp 1621261055
transform 1 0 12576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_127
timestamp 1621261055
transform 1 0 13344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_135
timestamp 1621261055
transform 1 0 14112 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _037_
timestamp 1621261055
transform -1 0 14880 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_89
timestamp 1621261055
transform -1 0 14592 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_137
timestamp 1621261055
transform 1 0 14304 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_143
timestamp 1621261055
transform 1 0 14880 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_151
timestamp 1621261055
transform 1 0 15648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_159
timestamp 1621261055
transform 1 0 16416 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_565
timestamp 1621261055
transform 1 0 16992 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_163
timestamp 1621261055
transform 1 0 16800 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_166
timestamp 1621261055
transform 1 0 17088 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_174
timestamp 1621261055
transform 1 0 17856 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_182
timestamp 1621261055
transform 1 0 18624 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_190
timestamp 1621261055
transform 1 0 19392 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_198
timestamp 1621261055
transform 1 0 20160 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_206
timestamp 1621261055
transform 1 0 20928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_214
timestamp 1621261055
transform 1 0 21696 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_566
timestamp 1621261055
transform 1 0 22272 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_218
timestamp 1621261055
transform 1 0 22080 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_221
timestamp 1621261055
transform 1 0 22368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_229
timestamp 1621261055
transform 1 0 23136 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_237
timestamp 1621261055
transform 1 0 23904 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_245
timestamp 1621261055
transform 1 0 24672 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_253
timestamp 1621261055
transform 1 0 25440 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_261
timestamp 1621261055
transform 1 0 26208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_269
timestamp 1621261055
transform 1 0 26976 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_567
timestamp 1621261055
transform 1 0 27552 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_273
timestamp 1621261055
transform 1 0 27360 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_276
timestamp 1621261055
transform 1 0 27648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_284
timestamp 1621261055
transform 1 0 28416 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_292
timestamp 1621261055
transform 1 0 29184 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_300
timestamp 1621261055
transform 1 0 29952 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_308
timestamp 1621261055
transform 1 0 30720 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_316
timestamp 1621261055
transform 1 0 31488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_324
timestamp 1621261055
transform 1 0 32256 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_568
timestamp 1621261055
transform 1 0 32832 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_328
timestamp 1621261055
transform 1 0 32640 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_331
timestamp 1621261055
transform 1 0 32928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_339
timestamp 1621261055
transform 1 0 33696 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_347
timestamp 1621261055
transform 1 0 34464 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_355
timestamp 1621261055
transform 1 0 35232 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_363
timestamp 1621261055
transform 1 0 36000 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_371
timestamp 1621261055
transform 1 0 36768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_569
timestamp 1621261055
transform 1 0 38112 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_379
timestamp 1621261055
transform 1 0 37536 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_383
timestamp 1621261055
transform 1 0 37920 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_386
timestamp 1621261055
transform 1 0 38208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_394
timestamp 1621261055
transform 1 0 38976 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_402
timestamp 1621261055
transform 1 0 39744 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_410
timestamp 1621261055
transform 1 0 40512 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_418
timestamp 1621261055
transform 1 0 41280 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_426
timestamp 1621261055
transform 1 0 42048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_570
timestamp 1621261055
transform 1 0 43392 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_434
timestamp 1621261055
transform 1 0 42816 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_438
timestamp 1621261055
transform 1 0 43200 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_441
timestamp 1621261055
transform 1 0 43488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_449
timestamp 1621261055
transform 1 0 44256 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_457
timestamp 1621261055
transform 1 0 45024 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_465
timestamp 1621261055
transform 1 0 45792 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_473
timestamp 1621261055
transform 1 0 46560 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_481
timestamp 1621261055
transform 1 0 47328 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_571
timestamp 1621261055
transform 1 0 48672 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_489
timestamp 1621261055
transform 1 0 48096 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_493
timestamp 1621261055
transform 1 0 48480 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_496
timestamp 1621261055
transform 1 0 48768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_504
timestamp 1621261055
transform 1 0 49536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_512
timestamp 1621261055
transform 1 0 50304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_520
timestamp 1621261055
transform 1 0 51072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_528
timestamp 1621261055
transform 1 0 51840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_536
timestamp 1621261055
transform 1 0 52608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_572
timestamp 1621261055
transform 1 0 53952 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_544
timestamp 1621261055
transform 1 0 53376 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_548
timestamp 1621261055
transform 1 0 53760 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_551
timestamp 1621261055
transform 1 0 54048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_559
timestamp 1621261055
transform 1 0 54816 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_567
timestamp 1621261055
transform 1 0 55584 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _088_
timestamp 1621261055
transform 1 0 57504 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_37_575
timestamp 1621261055
transform 1 0 56352 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_583
timestamp 1621261055
transform 1 0 57120 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_37_590
timestamp 1621261055
transform 1 0 57792 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_594
timestamp 1621261055
transform 1 0 58176 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_75
timestamp 1621261055
transform -1 0 58848 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_37_596
timestamp 1621261055
transform 1 0 58368 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_76
timestamp 1621261055
transform 1 0 1152 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_78
timestamp 1621261055
transform 1 0 1152 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_4
timestamp 1621261055
transform 1 0 1536 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_12
timestamp 1621261055
transform 1 0 2304 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_20
timestamp 1621261055
transform 1 0 3072 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_4
timestamp 1621261055
transform 1 0 1536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_12
timestamp 1621261055
transform 1 0 2304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_20
timestamp 1621261055
transform 1 0 3072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_28
timestamp 1621261055
transform 1 0 3840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_29
timestamp 1621261055
transform 1 0 3936 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_573
timestamp 1621261055
transform 1 0 3840 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_44
timestamp 1621261055
transform 1 0 5376 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_36
timestamp 1621261055
transform 1 0 4608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_37
timestamp 1621261055
transform 1 0 4704 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_52
timestamp 1621261055
transform 1 0 6144 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_53
timestamp 1621261055
transform 1 0 6240 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_45
timestamp 1621261055
transform 1 0 5472 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_54
timestamp 1621261055
transform 1 0 6336 0 1 28638
box -38 -49 134 715
use XOR2X1  XOR2X1
timestamp 1624893035
transform 1 0 7680 0 1 28638
box 0 -48 2016 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_584
timestamp 1621261055
transform 1 0 6432 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_61
timestamp 1621261055
transform 1 0 7008 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_69
timestamp 1621261055
transform 1 0 7776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_77
timestamp 1621261055
transform 1 0 8544 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_81
timestamp 1621261055
transform 1 0 8928 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_56
timestamp 1621261055
transform 1 0 6528 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_64
timestamp 1621261055
transform 1 0 7296 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_89
timestamp 1621261055
transform 1 0 9696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_38_88
timestamp 1621261055
transform 1 0 9600 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_84
timestamp 1621261055
transform 1 0 9216 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_574
timestamp 1621261055
transform 1 0 9120 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _186_
timestamp 1621261055
transform 1 0 9696 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_97
timestamp 1621261055
transform 1 0 10464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_92
timestamp 1621261055
transform 1 0 9984 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_105
timestamp 1621261055
transform 1 0 11232 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_100
timestamp 1621261055
transform 1 0 10752 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_108
timestamp 1621261055
transform 1 0 11520 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_585
timestamp 1621261055
transform 1 0 11712 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_116
timestamp 1621261055
transform 1 0 12288 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_124
timestamp 1621261055
transform 1 0 13056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_132
timestamp 1621261055
transform 1 0 13824 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_39_109
timestamp 1621261055
transform 1 0 11616 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_111
timestamp 1621261055
transform 1 0 11808 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_119
timestamp 1621261055
transform 1 0 12576 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_127
timestamp 1621261055
transform 1 0 13344 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_135
timestamp 1621261055
transform 1 0 14112 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_575
timestamp 1621261055
transform 1 0 14400 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_136
timestamp 1621261055
transform 1 0 14208 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_139
timestamp 1621261055
transform 1 0 14496 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_147
timestamp 1621261055
transform 1 0 15264 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_155
timestamp 1621261055
transform 1 0 16032 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_143
timestamp 1621261055
transform 1 0 14880 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_151
timestamp 1621261055
transform 1 0 15648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_159
timestamp 1621261055
transform 1 0 16416 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_586
timestamp 1621261055
transform 1 0 16992 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_163
timestamp 1621261055
transform 1 0 16800 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_171
timestamp 1621261055
transform 1 0 17568 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_179
timestamp 1621261055
transform 1 0 18336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_187
timestamp 1621261055
transform 1 0 19104 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_163
timestamp 1621261055
transform 1 0 16800 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_166
timestamp 1621261055
transform 1 0 17088 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_174
timestamp 1621261055
transform 1 0 17856 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_182
timestamp 1621261055
transform 1 0 18624 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_190
timestamp 1621261055
transform 1 0 19392 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_194
timestamp 1621261055
transform 1 0 19776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_191
timestamp 1621261055
transform 1 0 19488 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_576
timestamp 1621261055
transform 1 0 19680 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_206
timestamp 1621261055
transform 1 0 20928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_198
timestamp 1621261055
transform 1 0 20160 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_206
timestamp 1621261055
transform 1 0 20928 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_202
timestamp 1621261055
transform 1 0 20544 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_39_214
timestamp 1621261055
transform 1 0 21696 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_211
timestamp 1621261055
transform 1 0 21408 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _149_
timestamp 1621261055
transform 1 0 21120 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_587
timestamp 1621261055
transform 1 0 22272 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_219
timestamp 1621261055
transform 1 0 22176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_227
timestamp 1621261055
transform 1 0 22944 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_235
timestamp 1621261055
transform 1 0 23712 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_243
timestamp 1621261055
transform 1 0 24480 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_218
timestamp 1621261055
transform 1 0 22080 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_221
timestamp 1621261055
transform 1 0 22368 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_229
timestamp 1621261055
transform 1 0 23136 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_237
timestamp 1621261055
transform 1 0 23904 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_577
timestamp 1621261055
transform 1 0 24960 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_38_247
timestamp 1621261055
transform 1 0 24864 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_249
timestamp 1621261055
transform 1 0 25056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_257
timestamp 1621261055
transform 1 0 25824 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_265
timestamp 1621261055
transform 1 0 26592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_245
timestamp 1621261055
transform 1 0 24672 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_253
timestamp 1621261055
transform 1 0 25440 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_261
timestamp 1621261055
transform 1 0 26208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_269
timestamp 1621261055
transform 1 0 26976 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_588
timestamp 1621261055
transform 1 0 27552 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_273
timestamp 1621261055
transform 1 0 27360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_281
timestamp 1621261055
transform 1 0 28128 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_289
timestamp 1621261055
transform 1 0 28896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_297
timestamp 1621261055
transform 1 0 29664 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_273
timestamp 1621261055
transform 1 0 27360 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_276
timestamp 1621261055
transform 1 0 27648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_284
timestamp 1621261055
transform 1 0 28416 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_292
timestamp 1621261055
transform 1 0 29184 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_300
timestamp 1621261055
transform 1 0 29952 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_304
timestamp 1621261055
transform 1 0 30336 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_301
timestamp 1621261055
transform 1 0 30048 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_578
timestamp 1621261055
transform 1 0 30240 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_308
timestamp 1621261055
transform 1 0 30720 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_38_310
timestamp 1621261055
transform 1 0 30912 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_308
timestamp 1621261055
transform 1 0 30720 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_51
timestamp 1621261055
transform -1 0 31200 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _036_
timestamp 1621261055
transform -1 0 31488 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_316
timestamp 1621261055
transform 1 0 31488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_316
timestamp 1621261055
transform 1 0 31488 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_324
timestamp 1621261055
transform 1 0 32256 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_324
timestamp 1621261055
transform 1 0 32256 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_589
timestamp 1621261055
transform 1 0 32832 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_332
timestamp 1621261055
transform 1 0 33024 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_340
timestamp 1621261055
transform 1 0 33792 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_348
timestamp 1621261055
transform 1 0 34560 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_328
timestamp 1621261055
transform 1 0 32640 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_331
timestamp 1621261055
transform 1 0 32928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_339
timestamp 1621261055
transform 1 0 33696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_347
timestamp 1621261055
transform 1 0 34464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_579
timestamp 1621261055
transform 1 0 35520 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_356
timestamp 1621261055
transform 1 0 35328 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_359
timestamp 1621261055
transform 1 0 35616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_367
timestamp 1621261055
transform 1 0 36384 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_375
timestamp 1621261055
transform 1 0 37152 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_355
timestamp 1621261055
transform 1 0 35232 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_363
timestamp 1621261055
transform 1 0 36000 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_371
timestamp 1621261055
transform 1 0 36768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_590
timestamp 1621261055
transform 1 0 38112 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_383
timestamp 1621261055
transform 1 0 37920 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_391
timestamp 1621261055
transform 1 0 38688 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_399
timestamp 1621261055
transform 1 0 39456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_379
timestamp 1621261055
transform 1 0 37536 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_383
timestamp 1621261055
transform 1 0 37920 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_386
timestamp 1621261055
transform 1 0 38208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_394
timestamp 1621261055
transform 1 0 38976 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_402
timestamp 1621261055
transform 1 0 39744 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_580
timestamp 1621261055
transform 1 0 40800 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_407
timestamp 1621261055
transform 1 0 40224 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_411
timestamp 1621261055
transform 1 0 40608 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_414
timestamp 1621261055
transform 1 0 40896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_422
timestamp 1621261055
transform 1 0 41664 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_430
timestamp 1621261055
transform 1 0 42432 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_410
timestamp 1621261055
transform 1 0 40512 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_418
timestamp 1621261055
transform 1 0 41280 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_426
timestamp 1621261055
transform 1 0 42048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_591
timestamp 1621261055
transform 1 0 43392 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_438
timestamp 1621261055
transform 1 0 43200 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_446
timestamp 1621261055
transform 1 0 43968 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_454
timestamp 1621261055
transform 1 0 44736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_434
timestamp 1621261055
transform 1 0 42816 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_438
timestamp 1621261055
transform 1 0 43200 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_441
timestamp 1621261055
transform 1 0 43488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_449
timestamp 1621261055
transform 1 0 44256 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_457
timestamp 1621261055
transform 1 0 45024 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_465
timestamp 1621261055
transform 1 0 45792 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_466
timestamp 1621261055
transform 1 0 45888 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_462
timestamp 1621261055
transform 1 0 45504 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_473
timestamp 1621261055
transform 1 0 46560 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_469
timestamp 1621261055
transform 1 0 46176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_581
timestamp 1621261055
transform 1 0 46080 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_485
timestamp 1621261055
transform 1 0 47712 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_477
timestamp 1621261055
transform 1 0 46944 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_31
timestamp 1621261055
transform 1 0 47328 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _019_
timestamp 1621261055
transform 1 0 47520 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_486
timestamp 1621261055
transform 1 0 47808 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_592
timestamp 1621261055
transform 1 0 48672 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_493
timestamp 1621261055
transform 1 0 48480 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_501
timestamp 1621261055
transform 1 0 49248 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_509
timestamp 1621261055
transform 1 0 50016 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_494
timestamp 1621261055
transform 1 0 48576 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_496
timestamp 1621261055
transform 1 0 48768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_504
timestamp 1621261055
transform 1 0 49536 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_512
timestamp 1621261055
transform 1 0 50304 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_582
timestamp 1621261055
transform 1 0 51360 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_38_517
timestamp 1621261055
transform 1 0 50784 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_521
timestamp 1621261055
transform 1 0 51168 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_524
timestamp 1621261055
transform 1 0 51456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_532
timestamp 1621261055
transform 1 0 52224 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_540
timestamp 1621261055
transform 1 0 52992 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_520
timestamp 1621261055
transform 1 0 51072 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_528
timestamp 1621261055
transform 1 0 51840 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_536
timestamp 1621261055
transform 1 0 52608 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_593
timestamp 1621261055
transform 1 0 53952 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_548
timestamp 1621261055
transform 1 0 53760 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_556
timestamp 1621261055
transform 1 0 54528 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_564
timestamp 1621261055
transform 1 0 55296 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_544
timestamp 1621261055
transform 1 0 53376 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_548
timestamp 1621261055
transform 1 0 53760 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_39_551
timestamp 1621261055
transform 1 0 54048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_559
timestamp 1621261055
transform 1 0 54816 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_567
timestamp 1621261055
transform 1 0 55584 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_575
timestamp 1621261055
transform 1 0 56352 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_576
timestamp 1621261055
transform 1 0 56448 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_572
timestamp 1621261055
transform 1 0 56064 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_583
timestamp 1621261055
transform 1 0 57120 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_579
timestamp 1621261055
transform 1 0 56736 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_583
timestamp 1621261055
transform 1 0 56640 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _093_
timestamp 1621261055
transform 1 0 57120 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_39_591
timestamp 1621261055
transform 1 0 57888 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_586
timestamp 1621261055
transform 1 0 57408 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_594
timestamp 1621261055
transform 1 0 58176 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_77
timestamp 1621261055
transform -1 0 58848 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_79
timestamp 1621261055
transform -1 0 58848 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_38_596
timestamp 1621261055
transform 1 0 58368 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_595
timestamp 1621261055
transform 1 0 58272 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_80
timestamp 1621261055
transform 1 0 1152 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_40_4
timestamp 1621261055
transform 1 0 1536 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_12
timestamp 1621261055
transform 1 0 2304 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_20
timestamp 1621261055
transform 1 0 3072 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _021_
timestamp 1621261055
transform -1 0 6144 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_594
timestamp 1621261055
transform 1 0 3840 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_33
timestamp 1621261055
transform -1 0 5856 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_29
timestamp 1621261055
transform 1 0 3936 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_37
timestamp 1621261055
transform 1 0 4704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_45
timestamp 1621261055
transform 1 0 5472 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_52
timestamp 1621261055
transform 1 0 6144 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_60
timestamp 1621261055
transform 1 0 6912 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_68
timestamp 1621261055
transform 1 0 7680 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_76
timestamp 1621261055
transform 1 0 8448 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_80
timestamp 1621261055
transform 1 0 8832 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_595
timestamp 1621261055
transform 1 0 9120 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_40_82
timestamp 1621261055
transform 1 0 9024 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_84
timestamp 1621261055
transform 1 0 9216 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_92
timestamp 1621261055
transform 1 0 9984 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_100
timestamp 1621261055
transform 1 0 10752 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_108
timestamp 1621261055
transform 1 0 11520 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_116
timestamp 1621261055
transform 1 0 12288 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_124
timestamp 1621261055
transform 1 0 13056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_132
timestamp 1621261055
transform 1 0 13824 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_596
timestamp 1621261055
transform 1 0 14400 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_136
timestamp 1621261055
transform 1 0 14208 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_139
timestamp 1621261055
transform 1 0 14496 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_147
timestamp 1621261055
transform 1 0 15264 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_155
timestamp 1621261055
transform 1 0 16032 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _073_
timestamp 1621261055
transform 1 0 18144 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_40_163
timestamp 1621261055
transform 1 0 16800 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_171
timestamp 1621261055
transform 1 0 17568 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_175
timestamp 1621261055
transform 1 0 17952 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_180
timestamp 1621261055
transform 1 0 18432 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_188
timestamp 1621261055
transform 1 0 19200 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_597
timestamp 1621261055
transform 1 0 19680 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_40_192
timestamp 1621261055
transform 1 0 19584 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_194
timestamp 1621261055
transform 1 0 19776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_202
timestamp 1621261055
transform 1 0 20544 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_210
timestamp 1621261055
transform 1 0 21312 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_218
timestamp 1621261055
transform 1 0 22080 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_226
timestamp 1621261055
transform 1 0 22848 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_234
timestamp 1621261055
transform 1 0 23616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_242
timestamp 1621261055
transform 1 0 24384 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_598
timestamp 1621261055
transform 1 0 24960 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_246
timestamp 1621261055
transform 1 0 24768 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_249
timestamp 1621261055
transform 1 0 25056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_257
timestamp 1621261055
transform 1 0 25824 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_265
timestamp 1621261055
transform 1 0 26592 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_273
timestamp 1621261055
transform 1 0 27360 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_281
timestamp 1621261055
transform 1 0 28128 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_289
timestamp 1621261055
transform 1 0 28896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_297
timestamp 1621261055
transform 1 0 29664 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_599
timestamp 1621261055
transform 1 0 30240 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_301
timestamp 1621261055
transform 1 0 30048 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_304
timestamp 1621261055
transform 1 0 30336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_312
timestamp 1621261055
transform 1 0 31104 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_320
timestamp 1621261055
transform 1 0 31872 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_328
timestamp 1621261055
transform 1 0 32640 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_336
timestamp 1621261055
transform 1 0 33408 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_344
timestamp 1621261055
transform 1 0 34176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_600
timestamp 1621261055
transform 1 0 35520 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_352
timestamp 1621261055
transform 1 0 34944 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_356
timestamp 1621261055
transform 1 0 35328 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_359
timestamp 1621261055
transform 1 0 35616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_367
timestamp 1621261055
transform 1 0 36384 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_375
timestamp 1621261055
transform 1 0 37152 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_383
timestamp 1621261055
transform 1 0 37920 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_391
timestamp 1621261055
transform 1 0 38688 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_399
timestamp 1621261055
transform 1 0 39456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_601
timestamp 1621261055
transform 1 0 40800 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_407
timestamp 1621261055
transform 1 0 40224 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_411
timestamp 1621261055
transform 1 0 40608 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_414
timestamp 1621261055
transform 1 0 40896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_422
timestamp 1621261055
transform 1 0 41664 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_430
timestamp 1621261055
transform 1 0 42432 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_438
timestamp 1621261055
transform 1 0 43200 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_446
timestamp 1621261055
transform 1 0 43968 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_454
timestamp 1621261055
transform 1 0 44736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_602
timestamp 1621261055
transform 1 0 46080 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_462
timestamp 1621261055
transform 1 0 45504 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_466
timestamp 1621261055
transform 1 0 45888 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_469
timestamp 1621261055
transform 1 0 46176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_477
timestamp 1621261055
transform 1 0 46944 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_485
timestamp 1621261055
transform 1 0 47712 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_493
timestamp 1621261055
transform 1 0 48480 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_501
timestamp 1621261055
transform 1 0 49248 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_509
timestamp 1621261055
transform 1 0 50016 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_603
timestamp 1621261055
transform 1 0 51360 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_517
timestamp 1621261055
transform 1 0 50784 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_521
timestamp 1621261055
transform 1 0 51168 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_524
timestamp 1621261055
transform 1 0 51456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_532
timestamp 1621261055
transform 1 0 52224 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_540
timestamp 1621261055
transform 1 0 52992 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_548
timestamp 1621261055
transform 1 0 53760 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_556
timestamp 1621261055
transform 1 0 54528 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_564
timestamp 1621261055
transform 1 0 55296 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_604
timestamp 1621261055
transform 1 0 56640 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_40_572
timestamp 1621261055
transform 1 0 56064 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_576
timestamp 1621261055
transform 1 0 56448 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_579
timestamp 1621261055
transform 1 0 56736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_587
timestamp 1621261055
transform 1 0 57504 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_81
timestamp 1621261055
transform -1 0 58848 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_595
timestamp 1621261055
transform 1 0 58272 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_82
timestamp 1621261055
transform 1 0 1152 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_4
timestamp 1621261055
transform 1 0 1536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_12
timestamp 1621261055
transform 1 0 2304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_20
timestamp 1621261055
transform 1 0 3072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_28
timestamp 1621261055
transform 1 0 3840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_36
timestamp 1621261055
transform 1 0 4608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_44
timestamp 1621261055
transform 1 0 5376 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_52
timestamp 1621261055
transform 1 0 6144 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_41_54
timestamp 1621261055
transform 1 0 6336 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_605
timestamp 1621261055
transform 1 0 6432 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_56
timestamp 1621261055
transform 1 0 6528 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_64
timestamp 1621261055
transform 1 0 7296 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_72
timestamp 1621261055
transform 1 0 8064 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_80
timestamp 1621261055
transform 1 0 8832 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_88
timestamp 1621261055
transform 1 0 9600 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_96
timestamp 1621261055
transform 1 0 10368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_104
timestamp 1621261055
transform 1 0 11136 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_108
timestamp 1621261055
transform 1 0 11520 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_606
timestamp 1621261055
transform 1 0 11712 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_111
timestamp 1621261055
transform 1 0 11808 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_119
timestamp 1621261055
transform 1 0 12576 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_127
timestamp 1621261055
transform 1 0 13344 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_135
timestamp 1621261055
transform 1 0 14112 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _170_
timestamp 1621261055
transform 1 0 15936 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_41_143
timestamp 1621261055
transform 1 0 14880 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_151
timestamp 1621261055
transform 1 0 15648 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_41_153
timestamp 1621261055
transform 1 0 15840 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_157
timestamp 1621261055
transform 1 0 16224 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_607
timestamp 1621261055
transform 1 0 16992 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_166
timestamp 1621261055
transform 1 0 17088 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_174
timestamp 1621261055
transform 1 0 17856 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_182
timestamp 1621261055
transform 1 0 18624 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_190
timestamp 1621261055
transform 1 0 19392 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_198
timestamp 1621261055
transform 1 0 20160 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_206
timestamp 1621261055
transform 1 0 20928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_214
timestamp 1621261055
transform 1 0 21696 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_608
timestamp 1621261055
transform 1 0 22272 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_218
timestamp 1621261055
transform 1 0 22080 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_221
timestamp 1621261055
transform 1 0 22368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_229
timestamp 1621261055
transform 1 0 23136 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_237
timestamp 1621261055
transform 1 0 23904 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_245
timestamp 1621261055
transform 1 0 24672 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_253
timestamp 1621261055
transform 1 0 25440 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_261
timestamp 1621261055
transform 1 0 26208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_269
timestamp 1621261055
transform 1 0 26976 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_609
timestamp 1621261055
transform 1 0 27552 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_273
timestamp 1621261055
transform 1 0 27360 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_276
timestamp 1621261055
transform 1 0 27648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_284
timestamp 1621261055
transform 1 0 28416 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_292
timestamp 1621261055
transform 1 0 29184 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_300
timestamp 1621261055
transform 1 0 29952 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_308
timestamp 1621261055
transform 1 0 30720 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_316
timestamp 1621261055
transform 1 0 31488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_324
timestamp 1621261055
transform 1 0 32256 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_610
timestamp 1621261055
transform 1 0 32832 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_328
timestamp 1621261055
transform 1 0 32640 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_331
timestamp 1621261055
transform 1 0 32928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_339
timestamp 1621261055
transform 1 0 33696 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_347
timestamp 1621261055
transform 1 0 34464 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_355
timestamp 1621261055
transform 1 0 35232 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_363
timestamp 1621261055
transform 1 0 36000 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_371
timestamp 1621261055
transform 1 0 36768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_611
timestamp 1621261055
transform 1 0 38112 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_379
timestamp 1621261055
transform 1 0 37536 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_383
timestamp 1621261055
transform 1 0 37920 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_386
timestamp 1621261055
transform 1 0 38208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_394
timestamp 1621261055
transform 1 0 38976 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_402
timestamp 1621261055
transform 1 0 39744 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_410
timestamp 1621261055
transform 1 0 40512 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_418
timestamp 1621261055
transform 1 0 41280 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_426
timestamp 1621261055
transform 1 0 42048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_612
timestamp 1621261055
transform 1 0 43392 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_434
timestamp 1621261055
transform 1 0 42816 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_438
timestamp 1621261055
transform 1 0 43200 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_441
timestamp 1621261055
transform 1 0 43488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_449
timestamp 1621261055
transform 1 0 44256 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_457
timestamp 1621261055
transform 1 0 45024 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_465
timestamp 1621261055
transform 1 0 45792 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_473
timestamp 1621261055
transform 1 0 46560 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_481
timestamp 1621261055
transform 1 0 47328 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_613
timestamp 1621261055
transform 1 0 48672 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_489
timestamp 1621261055
transform 1 0 48096 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_493
timestamp 1621261055
transform 1 0 48480 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_496
timestamp 1621261055
transform 1 0 48768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_504
timestamp 1621261055
transform 1 0 49536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_512
timestamp 1621261055
transform 1 0 50304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_520
timestamp 1621261055
transform 1 0 51072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_528
timestamp 1621261055
transform 1 0 51840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_536
timestamp 1621261055
transform 1 0 52608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_614
timestamp 1621261055
transform 1 0 53952 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_544
timestamp 1621261055
transform 1 0 53376 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_548
timestamp 1621261055
transform 1 0 53760 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_551
timestamp 1621261055
transform 1 0 54048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_559
timestamp 1621261055
transform 1 0 54816 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_567
timestamp 1621261055
transform 1 0 55584 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_575
timestamp 1621261055
transform 1 0 56352 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_583
timestamp 1621261055
transform 1 0 57120 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_591
timestamp 1621261055
transform 1 0 57888 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_83
timestamp 1621261055
transform -1 0 58848 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_595
timestamp 1621261055
transform 1 0 58272 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_84
timestamp 1621261055
transform 1 0 1152 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_42_4
timestamp 1621261055
transform 1 0 1536 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_12
timestamp 1621261055
transform 1 0 2304 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_20
timestamp 1621261055
transform 1 0 3072 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_615
timestamp 1621261055
transform 1 0 3840 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_29
timestamp 1621261055
transform 1 0 3936 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_37
timestamp 1621261055
transform 1 0 4704 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_45
timestamp 1621261055
transform 1 0 5472 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_53
timestamp 1621261055
transform 1 0 6240 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _130_
timestamp 1621261055
transform 1 0 8064 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_190
timestamp 1621261055
transform 1 0 7872 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_61
timestamp 1621261055
transform 1 0 7008 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_42_69
timestamp 1621261055
transform 1 0 7776 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_75
timestamp 1621261055
transform 1 0 8352 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_616
timestamp 1621261055
transform 1 0 9120 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_84
timestamp 1621261055
transform 1 0 9216 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_92
timestamp 1621261055
transform 1 0 9984 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_100
timestamp 1621261055
transform 1 0 10752 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_108
timestamp 1621261055
transform 1 0 11520 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_116
timestamp 1621261055
transform 1 0 12288 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_124
timestamp 1621261055
transform 1 0 13056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_132
timestamp 1621261055
transform 1 0 13824 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_617
timestamp 1621261055
transform 1 0 14400 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_136
timestamp 1621261055
transform 1 0 14208 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_139
timestamp 1621261055
transform 1 0 14496 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_147
timestamp 1621261055
transform 1 0 15264 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_155
timestamp 1621261055
transform 1 0 16032 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_163
timestamp 1621261055
transform 1 0 16800 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_171
timestamp 1621261055
transform 1 0 17568 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_179
timestamp 1621261055
transform 1 0 18336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_187
timestamp 1621261055
transform 1 0 19104 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_618
timestamp 1621261055
transform 1 0 19680 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_191
timestamp 1621261055
transform 1 0 19488 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_194
timestamp 1621261055
transform 1 0 19776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_202
timestamp 1621261055
transform 1 0 20544 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_210
timestamp 1621261055
transform 1 0 21312 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_218
timestamp 1621261055
transform 1 0 22080 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_226
timestamp 1621261055
transform 1 0 22848 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_234
timestamp 1621261055
transform 1 0 23616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_242
timestamp 1621261055
transform 1 0 24384 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_619
timestamp 1621261055
transform 1 0 24960 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_246
timestamp 1621261055
transform 1 0 24768 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_249
timestamp 1621261055
transform 1 0 25056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_257
timestamp 1621261055
transform 1 0 25824 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_265
timestamp 1621261055
transform 1 0 26592 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_273
timestamp 1621261055
transform 1 0 27360 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_281
timestamp 1621261055
transform 1 0 28128 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_289
timestamp 1621261055
transform 1 0 28896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_297
timestamp 1621261055
transform 1 0 29664 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_620
timestamp 1621261055
transform 1 0 30240 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_301
timestamp 1621261055
transform 1 0 30048 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_304
timestamp 1621261055
transform 1 0 30336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_312
timestamp 1621261055
transform 1 0 31104 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_320
timestamp 1621261055
transform 1 0 31872 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_328
timestamp 1621261055
transform 1 0 32640 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_336
timestamp 1621261055
transform 1 0 33408 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_344
timestamp 1621261055
transform 1 0 34176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_621
timestamp 1621261055
transform 1 0 35520 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_352
timestamp 1621261055
transform 1 0 34944 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_356
timestamp 1621261055
transform 1 0 35328 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_359
timestamp 1621261055
transform 1 0 35616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_367
timestamp 1621261055
transform 1 0 36384 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_375
timestamp 1621261055
transform 1 0 37152 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_383
timestamp 1621261055
transform 1 0 37920 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_391
timestamp 1621261055
transform 1 0 38688 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_399
timestamp 1621261055
transform 1 0 39456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_622
timestamp 1621261055
transform 1 0 40800 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_407
timestamp 1621261055
transform 1 0 40224 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_411
timestamp 1621261055
transform 1 0 40608 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_414
timestamp 1621261055
transform 1 0 40896 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_422
timestamp 1621261055
transform 1 0 41664 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_430
timestamp 1621261055
transform 1 0 42432 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_438
timestamp 1621261055
transform 1 0 43200 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_446
timestamp 1621261055
transform 1 0 43968 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_454
timestamp 1621261055
transform 1 0 44736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_623
timestamp 1621261055
transform 1 0 46080 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_462
timestamp 1621261055
transform 1 0 45504 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_466
timestamp 1621261055
transform 1 0 45888 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_469
timestamp 1621261055
transform 1 0 46176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_477
timestamp 1621261055
transform 1 0 46944 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_485
timestamp 1621261055
transform 1 0 47712 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_493
timestamp 1621261055
transform 1 0 48480 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_501
timestamp 1621261055
transform 1 0 49248 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_509
timestamp 1621261055
transform 1 0 50016 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_624
timestamp 1621261055
transform 1 0 51360 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_517
timestamp 1621261055
transform 1 0 50784 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_521
timestamp 1621261055
transform 1 0 51168 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_524
timestamp 1621261055
transform 1 0 51456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_532
timestamp 1621261055
transform 1 0 52224 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_540
timestamp 1621261055
transform 1 0 52992 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _033_
timestamp 1621261055
transform 1 0 54528 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_548
timestamp 1621261055
transform 1 0 53760 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_559
timestamp 1621261055
transform 1 0 54816 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_567
timestamp 1621261055
transform 1 0 55584 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_625
timestamp 1621261055
transform 1 0 56640 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_575
timestamp 1621261055
transform 1 0 56352 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_42_577
timestamp 1621261055
transform 1 0 56544 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_579
timestamp 1621261055
transform 1 0 56736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_587
timestamp 1621261055
transform 1 0 57504 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_85
timestamp 1621261055
transform -1 0 58848 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_595
timestamp 1621261055
transform 1 0 58272 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_86
timestamp 1621261055
transform 1 0 1152 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_43_4
timestamp 1621261055
transform 1 0 1536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_12
timestamp 1621261055
transform 1 0 2304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_20
timestamp 1621261055
transform 1 0 3072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_28
timestamp 1621261055
transform 1 0 3840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_36
timestamp 1621261055
transform 1 0 4608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_44
timestamp 1621261055
transform 1 0 5376 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_52
timestamp 1621261055
transform 1 0 6144 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_54
timestamp 1621261055
transform 1 0 6336 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_626
timestamp 1621261055
transform 1 0 6432 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_56
timestamp 1621261055
transform 1 0 6528 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_64
timestamp 1621261055
transform 1 0 7296 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_72
timestamp 1621261055
transform 1 0 8064 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_80
timestamp 1621261055
transform 1 0 8832 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_88
timestamp 1621261055
transform 1 0 9600 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_96
timestamp 1621261055
transform 1 0 10368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_104
timestamp 1621261055
transform 1 0 11136 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_108
timestamp 1621261055
transform 1 0 11520 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_627
timestamp 1621261055
transform 1 0 11712 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_111
timestamp 1621261055
transform 1 0 11808 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_119
timestamp 1621261055
transform 1 0 12576 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_127
timestamp 1621261055
transform 1 0 13344 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_135
timestamp 1621261055
transform 1 0 14112 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_143
timestamp 1621261055
transform 1 0 14880 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_151
timestamp 1621261055
transform 1 0 15648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_159
timestamp 1621261055
transform 1 0 16416 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_628
timestamp 1621261055
transform 1 0 16992 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_163
timestamp 1621261055
transform 1 0 16800 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_166
timestamp 1621261055
transform 1 0 17088 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_174
timestamp 1621261055
transform 1 0 17856 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_182
timestamp 1621261055
transform 1 0 18624 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _173_
timestamp 1621261055
transform 1 0 21120 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_43_190
timestamp 1621261055
transform 1 0 19392 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_198
timestamp 1621261055
transform 1 0 20160 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_206
timestamp 1621261055
transform 1 0 20928 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_211
timestamp 1621261055
transform 1 0 21408 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_629
timestamp 1621261055
transform 1 0 22272 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_43_219
timestamp 1621261055
transform 1 0 22176 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_221
timestamp 1621261055
transform 1 0 22368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_229
timestamp 1621261055
transform 1 0 23136 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_237
timestamp 1621261055
transform 1 0 23904 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_245
timestamp 1621261055
transform 1 0 24672 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_253
timestamp 1621261055
transform 1 0 25440 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_261
timestamp 1621261055
transform 1 0 26208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_269
timestamp 1621261055
transform 1 0 26976 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _000_
timestamp 1621261055
transform 1 0 28992 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_630
timestamp 1621261055
transform 1 0 27552 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_273
timestamp 1621261055
transform 1 0 27360 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_276
timestamp 1621261055
transform 1 0 27648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_284
timestamp 1621261055
transform 1 0 28416 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_288
timestamp 1621261055
transform 1 0 28800 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_293
timestamp 1621261055
transform 1 0 29280 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_301
timestamp 1621261055
transform 1 0 30048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_309
timestamp 1621261055
transform 1 0 30816 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_317
timestamp 1621261055
transform 1 0 31584 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _116_
timestamp 1621261055
transform 1 0 34464 0 1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_631
timestamp 1621261055
transform 1 0 32832 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_325
timestamp 1621261055
transform 1 0 32352 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_43_329
timestamp 1621261055
transform 1 0 32736 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_331
timestamp 1621261055
transform 1 0 32928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_339
timestamp 1621261055
transform 1 0 33696 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_350
timestamp 1621261055
transform 1 0 34752 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_358
timestamp 1621261055
transform 1 0 35520 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_366
timestamp 1621261055
transform 1 0 36288 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_374
timestamp 1621261055
transform 1 0 37056 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_632
timestamp 1621261055
transform 1 0 38112 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_382
timestamp 1621261055
transform 1 0 37824 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_384
timestamp 1621261055
transform 1 0 38016 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_386
timestamp 1621261055
transform 1 0 38208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_394
timestamp 1621261055
transform 1 0 38976 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_402
timestamp 1621261055
transform 1 0 39744 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_410
timestamp 1621261055
transform 1 0 40512 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_418
timestamp 1621261055
transform 1 0 41280 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_426
timestamp 1621261055
transform 1 0 42048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_633
timestamp 1621261055
transform 1 0 43392 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_434
timestamp 1621261055
transform 1 0 42816 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_438
timestamp 1621261055
transform 1 0 43200 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_441
timestamp 1621261055
transform 1 0 43488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_449
timestamp 1621261055
transform 1 0 44256 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_457
timestamp 1621261055
transform 1 0 45024 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_465
timestamp 1621261055
transform 1 0 45792 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_473
timestamp 1621261055
transform 1 0 46560 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_481
timestamp 1621261055
transform 1 0 47328 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_634
timestamp 1621261055
transform 1 0 48672 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_489
timestamp 1621261055
transform 1 0 48096 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_493
timestamp 1621261055
transform 1 0 48480 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_496
timestamp 1621261055
transform 1 0 48768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_504
timestamp 1621261055
transform 1 0 49536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_512
timestamp 1621261055
transform 1 0 50304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_520
timestamp 1621261055
transform 1 0 51072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_528
timestamp 1621261055
transform 1 0 51840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_536
timestamp 1621261055
transform 1 0 52608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_635
timestamp 1621261055
transform 1 0 53952 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_544
timestamp 1621261055
transform 1 0 53376 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_548
timestamp 1621261055
transform 1 0 53760 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_551
timestamp 1621261055
transform 1 0 54048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_559
timestamp 1621261055
transform 1 0 54816 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_567
timestamp 1621261055
transform 1 0 55584 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_575
timestamp 1621261055
transform 1 0 56352 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_583
timestamp 1621261055
transform 1 0 57120 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_591
timestamp 1621261055
transform 1 0 57888 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_87
timestamp 1621261055
transform -1 0 58848 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_595
timestamp 1621261055
transform 1 0 58272 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_88
timestamp 1621261055
transform 1 0 1152 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_4
timestamp 1621261055
transform 1 0 1536 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_12
timestamp 1621261055
transform 1 0 2304 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_20
timestamp 1621261055
transform 1 0 3072 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_636
timestamp 1621261055
transform 1 0 3840 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_29
timestamp 1621261055
transform 1 0 3936 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_37
timestamp 1621261055
transform 1 0 4704 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_45
timestamp 1621261055
transform 1 0 5472 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_53
timestamp 1621261055
transform 1 0 6240 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _056_
timestamp 1621261055
transform 1 0 8256 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_44_61
timestamp 1621261055
transform 1 0 7008 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_69
timestamp 1621261055
transform 1 0 7776 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_44_73
timestamp 1621261055
transform 1 0 8160 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_77
timestamp 1621261055
transform 1 0 8544 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_81
timestamp 1621261055
transform 1 0 8928 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_637
timestamp 1621261055
transform 1 0 9120 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_84
timestamp 1621261055
transform 1 0 9216 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_92
timestamp 1621261055
transform 1 0 9984 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_100
timestamp 1621261055
transform 1 0 10752 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_108
timestamp 1621261055
transform 1 0 11520 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_116
timestamp 1621261055
transform 1 0 12288 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_124
timestamp 1621261055
transform 1 0 13056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_132
timestamp 1621261055
transform 1 0 13824 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_638
timestamp 1621261055
transform 1 0 14400 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_136
timestamp 1621261055
transform 1 0 14208 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_139
timestamp 1621261055
transform 1 0 14496 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_147
timestamp 1621261055
transform 1 0 15264 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_155
timestamp 1621261055
transform 1 0 16032 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_163
timestamp 1621261055
transform 1 0 16800 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_171
timestamp 1621261055
transform 1 0 17568 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_179
timestamp 1621261055
transform 1 0 18336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_187
timestamp 1621261055
transform 1 0 19104 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_639
timestamp 1621261055
transform 1 0 19680 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_191
timestamp 1621261055
transform 1 0 19488 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_194
timestamp 1621261055
transform 1 0 19776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_202
timestamp 1621261055
transform 1 0 20544 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_210
timestamp 1621261055
transform 1 0 21312 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_218
timestamp 1621261055
transform 1 0 22080 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_226
timestamp 1621261055
transform 1 0 22848 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_234
timestamp 1621261055
transform 1 0 23616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_242
timestamp 1621261055
transform 1 0 24384 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_640
timestamp 1621261055
transform 1 0 24960 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_246
timestamp 1621261055
transform 1 0 24768 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_249
timestamp 1621261055
transform 1 0 25056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_257
timestamp 1621261055
transform 1 0 25824 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_265
timestamp 1621261055
transform 1 0 26592 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_273
timestamp 1621261055
transform 1 0 27360 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_281
timestamp 1621261055
transform 1 0 28128 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_289
timestamp 1621261055
transform 1 0 28896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_297
timestamp 1621261055
transform 1 0 29664 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _158_
timestamp 1621261055
transform 1 0 31968 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_641
timestamp 1621261055
transform 1 0 30240 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_301
timestamp 1621261055
transform 1 0 30048 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_304
timestamp 1621261055
transform 1 0 30336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_312
timestamp 1621261055
transform 1 0 31104 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_44_320
timestamp 1621261055
transform 1 0 31872 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_324
timestamp 1621261055
transform 1 0 32256 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_332
timestamp 1621261055
transform 1 0 33024 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_340
timestamp 1621261055
transform 1 0 33792 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_348
timestamp 1621261055
transform 1 0 34560 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_642
timestamp 1621261055
transform 1 0 35520 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_356
timestamp 1621261055
transform 1 0 35328 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_359
timestamp 1621261055
transform 1 0 35616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_367
timestamp 1621261055
transform 1 0 36384 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_375
timestamp 1621261055
transform 1 0 37152 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_383
timestamp 1621261055
transform 1 0 37920 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_391
timestamp 1621261055
transform 1 0 38688 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_399
timestamp 1621261055
transform 1 0 39456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_643
timestamp 1621261055
transform 1 0 40800 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_407
timestamp 1621261055
transform 1 0 40224 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_411
timestamp 1621261055
transform 1 0 40608 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_414
timestamp 1621261055
transform 1 0 40896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_422
timestamp 1621261055
transform 1 0 41664 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_430
timestamp 1621261055
transform 1 0 42432 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _121_
timestamp 1621261055
transform 1 0 42816 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_44_437
timestamp 1621261055
transform 1 0 43104 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_445
timestamp 1621261055
transform 1 0 43872 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_453
timestamp 1621261055
transform 1 0 44640 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_644
timestamp 1621261055
transform 1 0 46080 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_461
timestamp 1621261055
transform 1 0 45408 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_465
timestamp 1621261055
transform 1 0 45792 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_44_467
timestamp 1621261055
transform 1 0 45984 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_469
timestamp 1621261055
transform 1 0 46176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_477
timestamp 1621261055
transform 1 0 46944 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_485
timestamp 1621261055
transform 1 0 47712 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_493
timestamp 1621261055
transform 1 0 48480 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_501
timestamp 1621261055
transform 1 0 49248 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_509
timestamp 1621261055
transform 1 0 50016 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_645
timestamp 1621261055
transform 1 0 51360 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_517
timestamp 1621261055
transform 1 0 50784 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_521
timestamp 1621261055
transform 1 0 51168 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_524
timestamp 1621261055
transform 1 0 51456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_532
timestamp 1621261055
transform 1 0 52224 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_540
timestamp 1621261055
transform 1 0 52992 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_548
timestamp 1621261055
transform 1 0 53760 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_556
timestamp 1621261055
transform 1 0 54528 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_564
timestamp 1621261055
transform 1 0 55296 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_646
timestamp 1621261055
transform 1 0 56640 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_44_572
timestamp 1621261055
transform 1 0 56064 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_576
timestamp 1621261055
transform 1 0 56448 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_579
timestamp 1621261055
transform 1 0 56736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_587
timestamp 1621261055
transform 1 0 57504 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_89
timestamp 1621261055
transform -1 0 58848 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_595
timestamp 1621261055
transform 1 0 58272 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _015_
timestamp 1621261055
transform 1 0 2496 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_90
timestamp 1621261055
transform 1 0 1152 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_4
timestamp 1621261055
transform 1 0 1536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_12
timestamp 1621261055
transform 1 0 2304 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_17
timestamp 1621261055
transform 1 0 2784 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_25
timestamp 1621261055
transform 1 0 3552 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_33
timestamp 1621261055
transform 1 0 4320 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_41
timestamp 1621261055
transform 1 0 5088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_49
timestamp 1621261055
transform 1 0 5856 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_53
timestamp 1621261055
transform 1 0 6240 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_647
timestamp 1621261055
transform 1 0 6432 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_56
timestamp 1621261055
transform 1 0 6528 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_64
timestamp 1621261055
transform 1 0 7296 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_72
timestamp 1621261055
transform 1 0 8064 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_80
timestamp 1621261055
transform 1 0 8832 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_88
timestamp 1621261055
transform 1 0 9600 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_96
timestamp 1621261055
transform 1 0 10368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_104
timestamp 1621261055
transform 1 0 11136 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_108
timestamp 1621261055
transform 1 0 11520 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_648
timestamp 1621261055
transform 1 0 11712 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_111
timestamp 1621261055
transform 1 0 11808 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_119
timestamp 1621261055
transform 1 0 12576 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_127
timestamp 1621261055
transform 1 0 13344 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_135
timestamp 1621261055
transform 1 0 14112 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_143
timestamp 1621261055
transform 1 0 14880 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_151
timestamp 1621261055
transform 1 0 15648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_159
timestamp 1621261055
transform 1 0 16416 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_649
timestamp 1621261055
transform 1 0 16992 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_163
timestamp 1621261055
transform 1 0 16800 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_166
timestamp 1621261055
transform 1 0 17088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_174
timestamp 1621261055
transform 1 0 17856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_182
timestamp 1621261055
transform 1 0 18624 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_190
timestamp 1621261055
transform 1 0 19392 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_198
timestamp 1621261055
transform 1 0 20160 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_206
timestamp 1621261055
transform 1 0 20928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_214
timestamp 1621261055
transform 1 0 21696 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_650
timestamp 1621261055
transform 1 0 22272 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_218
timestamp 1621261055
transform 1 0 22080 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_221
timestamp 1621261055
transform 1 0 22368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_229
timestamp 1621261055
transform 1 0 23136 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_237
timestamp 1621261055
transform 1 0 23904 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_245
timestamp 1621261055
transform 1 0 24672 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_253
timestamp 1621261055
transform 1 0 25440 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_261
timestamp 1621261055
transform 1 0 26208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_269
timestamp 1621261055
transform 1 0 26976 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_651
timestamp 1621261055
transform 1 0 27552 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_273
timestamp 1621261055
transform 1 0 27360 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_276
timestamp 1621261055
transform 1 0 27648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_284
timestamp 1621261055
transform 1 0 28416 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_292
timestamp 1621261055
transform 1 0 29184 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_300
timestamp 1621261055
transform 1 0 29952 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_308
timestamp 1621261055
transform 1 0 30720 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_316
timestamp 1621261055
transform 1 0 31488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_324
timestamp 1621261055
transform 1 0 32256 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_652
timestamp 1621261055
transform 1 0 32832 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_328
timestamp 1621261055
transform 1 0 32640 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_331
timestamp 1621261055
transform 1 0 32928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_339
timestamp 1621261055
transform 1 0 33696 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_347
timestamp 1621261055
transform 1 0 34464 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_355
timestamp 1621261055
transform 1 0 35232 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_363
timestamp 1621261055
transform 1 0 36000 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_371
timestamp 1621261055
transform 1 0 36768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _106_
timestamp 1621261055
transform -1 0 40320 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_653
timestamp 1621261055
transform 1 0 38112 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_167
timestamp 1621261055
transform -1 0 40032 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_45_379
timestamp 1621261055
transform 1 0 37536 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_383
timestamp 1621261055
transform 1 0 37920 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_386
timestamp 1621261055
transform 1 0 38208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_394
timestamp 1621261055
transform 1 0 38976 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_45_402
timestamp 1621261055
transform 1 0 39744 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_408
timestamp 1621261055
transform 1 0 40320 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_416
timestamp 1621261055
transform 1 0 41088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_424
timestamp 1621261055
transform 1 0 41856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_432
timestamp 1621261055
transform 1 0 42624 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _054_
timestamp 1621261055
transform 1 0 44544 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_654
timestamp 1621261055
transform 1 0 43392 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_441
timestamp 1621261055
transform 1 0 43488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_449
timestamp 1621261055
transform 1 0 44256 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_451
timestamp 1621261055
transform 1 0 44448 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_455
timestamp 1621261055
transform 1 0 44832 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _092_
timestamp 1621261055
transform -1 0 47232 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_153
timestamp 1621261055
transform -1 0 46944 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_463
timestamp 1621261055
transform 1 0 45600 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_471
timestamp 1621261055
transform 1 0 46368 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_480
timestamp 1621261055
transform 1 0 47232 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_655
timestamp 1621261055
transform 1 0 48672 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_488
timestamp 1621261055
transform 1 0 48000 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_492
timestamp 1621261055
transform 1 0 48384 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_494
timestamp 1621261055
transform 1 0 48576 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_496
timestamp 1621261055
transform 1 0 48768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_504
timestamp 1621261055
transform 1 0 49536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_512
timestamp 1621261055
transform 1 0 50304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_520
timestamp 1621261055
transform 1 0 51072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_528
timestamp 1621261055
transform 1 0 51840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_536
timestamp 1621261055
transform 1 0 52608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_656
timestamp 1621261055
transform 1 0 53952 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_544
timestamp 1621261055
transform 1 0 53376 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_548
timestamp 1621261055
transform 1 0 53760 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_551
timestamp 1621261055
transform 1 0 54048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_559
timestamp 1621261055
transform 1 0 54816 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_567
timestamp 1621261055
transform 1 0 55584 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_575
timestamp 1621261055
transform 1 0 56352 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_583
timestamp 1621261055
transform 1 0 57120 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_591
timestamp 1621261055
transform 1 0 57888 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_91
timestamp 1621261055
transform -1 0 58848 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_595
timestamp 1621261055
transform 1 0 58272 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_92
timestamp 1621261055
transform 1 0 1152 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_94
timestamp 1621261055
transform 1 0 1152 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_4
timestamp 1621261055
transform 1 0 1536 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_12
timestamp 1621261055
transform 1 0 2304 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_20
timestamp 1621261055
transform 1 0 3072 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_4
timestamp 1621261055
transform 1 0 1536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_12
timestamp 1621261055
transform 1 0 2304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_20
timestamp 1621261055
transform 1 0 3072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_28
timestamp 1621261055
transform 1 0 3840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_29
timestamp 1621261055
transform 1 0 3936 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_657
timestamp 1621261055
transform 1 0 3840 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_44
timestamp 1621261055
transform 1 0 5376 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_36
timestamp 1621261055
transform 1 0 4608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_37
timestamp 1621261055
transform 1 0 4704 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_52
timestamp 1621261055
transform 1 0 6144 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_53
timestamp 1621261055
transform 1 0 6240 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_45
timestamp 1621261055
transform 1 0 5472 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_54
timestamp 1621261055
transform 1 0 6336 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_668
timestamp 1621261055
transform 1 0 6432 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_61
timestamp 1621261055
transform 1 0 7008 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_69
timestamp 1621261055
transform 1 0 7776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_77
timestamp 1621261055
transform 1 0 8544 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_81
timestamp 1621261055
transform 1 0 8928 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_56
timestamp 1621261055
transform 1 0 6528 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_64
timestamp 1621261055
transform 1 0 7296 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_72
timestamp 1621261055
transform 1 0 8064 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_80
timestamp 1621261055
transform 1 0 8832 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_658
timestamp 1621261055
transform 1 0 9120 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_84
timestamp 1621261055
transform 1 0 9216 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_92
timestamp 1621261055
transform 1 0 9984 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_100
timestamp 1621261055
transform 1 0 10752 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_108
timestamp 1621261055
transform 1 0 11520 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_88
timestamp 1621261055
transform 1 0 9600 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_96
timestamp 1621261055
transform 1 0 10368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_104
timestamp 1621261055
transform 1 0 11136 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_108
timestamp 1621261055
transform 1 0 11520 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_669
timestamp 1621261055
transform 1 0 11712 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_116
timestamp 1621261055
transform 1 0 12288 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_124
timestamp 1621261055
transform 1 0 13056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_132
timestamp 1621261055
transform 1 0 13824 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_111
timestamp 1621261055
transform 1 0 11808 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_119
timestamp 1621261055
transform 1 0 12576 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_127
timestamp 1621261055
transform 1 0 13344 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_135
timestamp 1621261055
transform 1 0 14112 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_659
timestamp 1621261055
transform 1 0 14400 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_136
timestamp 1621261055
transform 1 0 14208 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_139
timestamp 1621261055
transform 1 0 14496 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_147
timestamp 1621261055
transform 1 0 15264 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_155
timestamp 1621261055
transform 1 0 16032 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_143
timestamp 1621261055
transform 1 0 14880 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_151
timestamp 1621261055
transform 1 0 15648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_159
timestamp 1621261055
transform 1 0 16416 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_166
timestamp 1621261055
transform 1 0 17088 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_163
timestamp 1621261055
transform 1 0 16800 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_46_165
timestamp 1621261055
transform 1 0 16992 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_163
timestamp 1621261055
transform 1 0 16800 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_172
timestamp 1621261055
transform -1 0 17280 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_670
timestamp 1621261055
transform 1 0 16992 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _063_
timestamp 1621261055
transform -1 0 17568 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_174
timestamp 1621261055
transform 1 0 17856 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_179
timestamp 1621261055
transform 1 0 18336 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_171
timestamp 1621261055
transform 1 0 17568 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_182
timestamp 1621261055
transform 1 0 18624 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_184
timestamp 1621261055
transform 1 0 18816 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _032_
timestamp 1621261055
transform 1 0 18528 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_660
timestamp 1621261055
transform 1 0 19680 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_46_192
timestamp 1621261055
transform 1 0 19584 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_194
timestamp 1621261055
transform 1 0 19776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_202
timestamp 1621261055
transform 1 0 20544 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_210
timestamp 1621261055
transform 1 0 21312 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_190
timestamp 1621261055
transform 1 0 19392 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_198
timestamp 1621261055
transform 1 0 20160 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_206
timestamp 1621261055
transform 1 0 20928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_214
timestamp 1621261055
transform 1 0 21696 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_47_221
timestamp 1621261055
transform 1 0 22368 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_218
timestamp 1621261055
transform 1 0 22080 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_218
timestamp 1621261055
transform 1 0 22080 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_671
timestamp 1621261055
transform 1 0 22272 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_228
timestamp 1621261055
transform 1 0 23040 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_226
timestamp 1621261055
transform 1 0 22848 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _211_
timestamp 1621261055
transform 1 0 22752 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_236
timestamp 1621261055
transform 1 0 23808 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_242
timestamp 1621261055
transform 1 0 24384 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_234
timestamp 1621261055
transform 1 0 23616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_661
timestamp 1621261055
transform 1 0 24960 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_246
timestamp 1621261055
transform 1 0 24768 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_249
timestamp 1621261055
transform 1 0 25056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_257
timestamp 1621261055
transform 1 0 25824 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_265
timestamp 1621261055
transform 1 0 26592 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_244
timestamp 1621261055
transform 1 0 24576 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_252
timestamp 1621261055
transform 1 0 25344 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_260
timestamp 1621261055
transform 1 0 26112 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_268
timestamp 1621261055
transform 1 0 26880 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_276
timestamp 1621261055
transform 1 0 27648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_274
timestamp 1621261055
transform 1 0 27456 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_272
timestamp 1621261055
transform 1 0 27264 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_273
timestamp 1621261055
transform 1 0 27360 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_672
timestamp 1621261055
transform 1 0 27552 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_284
timestamp 1621261055
transform 1 0 28416 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_286
timestamp 1621261055
transform 1 0 28608 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_235
timestamp 1621261055
transform -1 0 28320 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _203_
timestamp 1621261055
transform -1 0 28608 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_292
timestamp 1621261055
transform 1 0 29184 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_294
timestamp 1621261055
transform 1 0 29376 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_662
timestamp 1621261055
transform 1 0 30240 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_46_302
timestamp 1621261055
transform 1 0 30144 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_304
timestamp 1621261055
transform 1 0 30336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_312
timestamp 1621261055
transform 1 0 31104 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_320
timestamp 1621261055
transform 1 0 31872 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_300
timestamp 1621261055
transform 1 0 29952 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_308
timestamp 1621261055
transform 1 0 30720 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_316
timestamp 1621261055
transform 1 0 31488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_324
timestamp 1621261055
transform 1 0 32256 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_673
timestamp 1621261055
transform 1 0 32832 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_328
timestamp 1621261055
transform 1 0 32640 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_336
timestamp 1621261055
transform 1 0 33408 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_344
timestamp 1621261055
transform 1 0 34176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_328
timestamp 1621261055
transform 1 0 32640 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_331
timestamp 1621261055
transform 1 0 32928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_339
timestamp 1621261055
transform 1 0 33696 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_347
timestamp 1621261055
transform 1 0 34464 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_663
timestamp 1621261055
transform 1 0 35520 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_352
timestamp 1621261055
transform 1 0 34944 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_356
timestamp 1621261055
transform 1 0 35328 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_359
timestamp 1621261055
transform 1 0 35616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_367
timestamp 1621261055
transform 1 0 36384 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_375
timestamp 1621261055
transform 1 0 37152 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_355
timestamp 1621261055
transform 1 0 35232 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_363
timestamp 1621261055
transform 1 0 36000 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_371
timestamp 1621261055
transform 1 0 36768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_674
timestamp 1621261055
transform 1 0 38112 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_383
timestamp 1621261055
transform 1 0 37920 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_391
timestamp 1621261055
transform 1 0 38688 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_399
timestamp 1621261055
transform 1 0 39456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_379
timestamp 1621261055
transform 1 0 37536 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_383
timestamp 1621261055
transform 1 0 37920 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_386
timestamp 1621261055
transform 1 0 38208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_394
timestamp 1621261055
transform 1 0 38976 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_402
timestamp 1621261055
transform 1 0 39744 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_664
timestamp 1621261055
transform 1 0 40800 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_407
timestamp 1621261055
transform 1 0 40224 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_411
timestamp 1621261055
transform 1 0 40608 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_414
timestamp 1621261055
transform 1 0 40896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_422
timestamp 1621261055
transform 1 0 41664 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_430
timestamp 1621261055
transform 1 0 42432 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_410
timestamp 1621261055
transform 1 0 40512 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_418
timestamp 1621261055
transform 1 0 41280 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_426
timestamp 1621261055
transform 1 0 42048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_438
timestamp 1621261055
transform 1 0 43200 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_434
timestamp 1621261055
transform 1 0 42816 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_438
timestamp 1621261055
transform 1 0 43200 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_434
timestamp 1621261055
transform 1 0 42816 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_675
timestamp 1621261055
transform 1 0 43392 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _212_
timestamp 1621261055
transform 1 0 42912 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_449
timestamp 1621261055
transform 1 0 44256 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_441
timestamp 1621261055
transform 1 0 43488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_446
timestamp 1621261055
transform 1 0 43968 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_457
timestamp 1621261055
transform 1 0 45024 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_454
timestamp 1621261055
transform 1 0 44736 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_665
timestamp 1621261055
transform 1 0 46080 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_462
timestamp 1621261055
transform 1 0 45504 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_466
timestamp 1621261055
transform 1 0 45888 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_469
timestamp 1621261055
transform 1 0 46176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_477
timestamp 1621261055
transform 1 0 46944 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_485
timestamp 1621261055
transform 1 0 47712 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_465
timestamp 1621261055
transform 1 0 45792 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_473
timestamp 1621261055
transform 1 0 46560 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_481
timestamp 1621261055
transform 1 0 47328 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_676
timestamp 1621261055
transform 1 0 48672 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_493
timestamp 1621261055
transform 1 0 48480 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_501
timestamp 1621261055
transform 1 0 49248 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_509
timestamp 1621261055
transform 1 0 50016 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_489
timestamp 1621261055
transform 1 0 48096 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_493
timestamp 1621261055
transform 1 0 48480 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_496
timestamp 1621261055
transform 1 0 48768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_504
timestamp 1621261055
transform 1 0 49536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_512
timestamp 1621261055
transform 1 0 50304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_666
timestamp 1621261055
transform 1 0 51360 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_517
timestamp 1621261055
transform 1 0 50784 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_521
timestamp 1621261055
transform 1 0 51168 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_524
timestamp 1621261055
transform 1 0 51456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_532
timestamp 1621261055
transform 1 0 52224 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_540
timestamp 1621261055
transform 1 0 52992 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_520
timestamp 1621261055
transform 1 0 51072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_528
timestamp 1621261055
transform 1 0 51840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_536
timestamp 1621261055
transform 1 0 52608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _175_
timestamp 1621261055
transform 1 0 55584 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_677
timestamp 1621261055
transform 1 0 53952 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_548
timestamp 1621261055
transform 1 0 53760 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_556
timestamp 1621261055
transform 1 0 54528 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_564
timestamp 1621261055
transform 1 0 55296 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_544
timestamp 1621261055
transform 1 0 53376 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_548
timestamp 1621261055
transform 1 0 53760 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_551
timestamp 1621261055
transform 1 0 54048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_559
timestamp 1621261055
transform 1 0 54816 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_570
timestamp 1621261055
transform 1 0 55872 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_576
timestamp 1621261055
transform 1 0 56448 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_572
timestamp 1621261055
transform 1 0 56064 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_578
timestamp 1621261055
transform 1 0 56640 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_583
timestamp 1621261055
transform 1 0 57120 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_579
timestamp 1621261055
transform 1 0 56736 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_667
timestamp 1621261055
transform 1 0 56640 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_586
timestamp 1621261055
transform 1 0 57408 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_589
timestamp 1621261055
transform 1 0 57696 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_585
timestamp 1621261055
transform 1 0 57312 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _112_
timestamp 1621261055
transform 1 0 57408 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_594
timestamp 1621261055
transform 1 0 58176 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_93
timestamp 1621261055
transform -1 0 58848 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_95
timestamp 1621261055
transform -1 0 58848 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_47_596
timestamp 1621261055
transform 1 0 58368 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_96
timestamp 1621261055
transform 1 0 1152 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_4
timestamp 1621261055
transform 1 0 1536 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_12
timestamp 1621261055
transform 1 0 2304 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_20
timestamp 1621261055
transform 1 0 3072 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _040_
timestamp 1621261055
transform 1 0 5856 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_678
timestamp 1621261055
transform 1 0 3840 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_29
timestamp 1621261055
transform 1 0 3936 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_37
timestamp 1621261055
transform 1 0 4704 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_45
timestamp 1621261055
transform 1 0 5472 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_52
timestamp 1621261055
transform 1 0 6144 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_60
timestamp 1621261055
transform 1 0 6912 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_68
timestamp 1621261055
transform 1 0 7680 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_76
timestamp 1621261055
transform 1 0 8448 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_80
timestamp 1621261055
transform 1 0 8832 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_679
timestamp 1621261055
transform 1 0 9120 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_48_82
timestamp 1621261055
transform 1 0 9024 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_84
timestamp 1621261055
transform 1 0 9216 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_92
timestamp 1621261055
transform 1 0 9984 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_100
timestamp 1621261055
transform 1 0 10752 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_108
timestamp 1621261055
transform 1 0 11520 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_116
timestamp 1621261055
transform 1 0 12288 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_124
timestamp 1621261055
transform 1 0 13056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_132
timestamp 1621261055
transform 1 0 13824 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_680
timestamp 1621261055
transform 1 0 14400 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_136
timestamp 1621261055
transform 1 0 14208 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_139
timestamp 1621261055
transform 1 0 14496 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_147
timestamp 1621261055
transform 1 0 15264 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_155
timestamp 1621261055
transform 1 0 16032 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_163
timestamp 1621261055
transform 1 0 16800 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_171
timestamp 1621261055
transform 1 0 17568 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_179
timestamp 1621261055
transform 1 0 18336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_187
timestamp 1621261055
transform 1 0 19104 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _117_
timestamp 1621261055
transform 1 0 21120 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_681
timestamp 1621261055
transform 1 0 19680 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_176
timestamp 1621261055
transform 1 0 20928 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_191
timestamp 1621261055
transform 1 0 19488 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_194
timestamp 1621261055
transform 1 0 19776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_202
timestamp 1621261055
transform 1 0 20544 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_211
timestamp 1621261055
transform 1 0 21408 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _205_
timestamp 1621261055
transform -1 0 23232 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_237
timestamp 1621261055
transform -1 0 22944 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_219
timestamp 1621261055
transform 1 0 22176 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_223
timestamp 1621261055
transform 1 0 22560 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_230
timestamp 1621261055
transform 1 0 23232 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_238
timestamp 1621261055
transform 1 0 24000 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_682
timestamp 1621261055
transform 1 0 24960 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_246
timestamp 1621261055
transform 1 0 24768 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_249
timestamp 1621261055
transform 1 0 25056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_257
timestamp 1621261055
transform 1 0 25824 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_265
timestamp 1621261055
transform 1 0 26592 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _068_
timestamp 1621261055
transform -1 0 28992 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_131
timestamp 1621261055
transform -1 0 28704 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_273
timestamp 1621261055
transform 1 0 27360 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_281
timestamp 1621261055
transform 1 0 28128 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_48_290
timestamp 1621261055
transform 1 0 28992 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_683
timestamp 1621261055
transform 1 0 30240 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_298
timestamp 1621261055
transform 1 0 29760 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_48_302
timestamp 1621261055
transform 1 0 30144 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_304
timestamp 1621261055
transform 1 0 30336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_312
timestamp 1621261055
transform 1 0 31104 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_320
timestamp 1621261055
transform 1 0 31872 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _027_
timestamp 1621261055
transform 1 0 32928 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_328
timestamp 1621261055
transform 1 0 32640 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_330
timestamp 1621261055
transform 1 0 32832 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_334
timestamp 1621261055
transform 1 0 33216 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_342
timestamp 1621261055
transform 1 0 33984 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_350
timestamp 1621261055
transform 1 0 34752 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_684
timestamp 1621261055
transform 1 0 35520 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_359
timestamp 1621261055
transform 1 0 35616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_367
timestamp 1621261055
transform 1 0 36384 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_375
timestamp 1621261055
transform 1 0 37152 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_383
timestamp 1621261055
transform 1 0 37920 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_391
timestamp 1621261055
transform 1 0 38688 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_399
timestamp 1621261055
transform 1 0 39456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_685
timestamp 1621261055
transform 1 0 40800 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_407
timestamp 1621261055
transform 1 0 40224 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_411
timestamp 1621261055
transform 1 0 40608 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_414
timestamp 1621261055
transform 1 0 40896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_422
timestamp 1621261055
transform 1 0 41664 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_430
timestamp 1621261055
transform 1 0 42432 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_438
timestamp 1621261055
transform 1 0 43200 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_446
timestamp 1621261055
transform 1 0 43968 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_454
timestamp 1621261055
transform 1 0 44736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_686
timestamp 1621261055
transform 1 0 46080 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_48_462
timestamp 1621261055
transform 1 0 45504 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_466
timestamp 1621261055
transform 1 0 45888 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_469
timestamp 1621261055
transform 1 0 46176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_477
timestamp 1621261055
transform 1 0 46944 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_485
timestamp 1621261055
transform 1 0 47712 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_493
timestamp 1621261055
transform 1 0 48480 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_501
timestamp 1621261055
transform 1 0 49248 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_509
timestamp 1621261055
transform 1 0 50016 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_521
timestamp 1621261055
transform 1 0 51168 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_517
timestamp 1621261055
transform 1 0 50784 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_524
timestamp 1621261055
transform 1 0 51456 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_141
timestamp 1621261055
transform -1 0 51840 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_687
timestamp 1621261055
transform 1 0 51360 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _075_
timestamp 1621261055
transform -1 0 52128 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_48_538
timestamp 1621261055
transform 1 0 52800 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_531
timestamp 1621261055
transform 1 0 52128 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_195
timestamp 1621261055
transform -1 0 52512 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _135_
timestamp 1621261055
transform -1 0 52800 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_48_546
timestamp 1621261055
transform 1 0 53568 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_554
timestamp 1621261055
transform 1 0 54336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_562
timestamp 1621261055
transform 1 0 55104 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_688
timestamp 1621261055
transform 1 0 56640 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_570
timestamp 1621261055
transform 1 0 55872 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_579
timestamp 1621261055
transform 1 0 56736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_587
timestamp 1621261055
transform 1 0 57504 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_97
timestamp 1621261055
transform -1 0 58848 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_595
timestamp 1621261055
transform 1 0 58272 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_98
timestamp 1621261055
transform 1 0 1152 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_49_4
timestamp 1621261055
transform 1 0 1536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_12
timestamp 1621261055
transform 1 0 2304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_20
timestamp 1621261055
transform 1 0 3072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_28
timestamp 1621261055
transform 1 0 3840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_36
timestamp 1621261055
transform 1 0 4608 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_44
timestamp 1621261055
transform 1 0 5376 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_52
timestamp 1621261055
transform 1 0 6144 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_54
timestamp 1621261055
transform 1 0 6336 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_689
timestamp 1621261055
transform 1 0 6432 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_56
timestamp 1621261055
transform 1 0 6528 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_64
timestamp 1621261055
transform 1 0 7296 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_72
timestamp 1621261055
transform 1 0 8064 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_80
timestamp 1621261055
transform 1 0 8832 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_88
timestamp 1621261055
transform 1 0 9600 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_96
timestamp 1621261055
transform 1 0 10368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_104
timestamp 1621261055
transform 1 0 11136 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_108
timestamp 1621261055
transform 1 0 11520 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _191_
timestamp 1621261055
transform -1 0 13536 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_690
timestamp 1621261055
transform 1 0 11712 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_251
timestamp 1621261055
transform -1 0 13248 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_111
timestamp 1621261055
transform 1 0 11808 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_119
timestamp 1621261055
transform 1 0 12576 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_49_123
timestamp 1621261055
transform 1 0 12960 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_129
timestamp 1621261055
transform 1 0 13536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_137
timestamp 1621261055
transform 1 0 14304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_145
timestamp 1621261055
transform 1 0 15072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_153
timestamp 1621261055
transform 1 0 15840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_161
timestamp 1621261055
transform 1 0 16608 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_691
timestamp 1621261055
transform 1 0 16992 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_166
timestamp 1621261055
transform 1 0 17088 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_174
timestamp 1621261055
transform 1 0 17856 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_182
timestamp 1621261055
transform 1 0 18624 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_190
timestamp 1621261055
transform 1 0 19392 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_198
timestamp 1621261055
transform 1 0 20160 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_206
timestamp 1621261055
transform 1 0 20928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_214
timestamp 1621261055
transform 1 0 21696 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_692
timestamp 1621261055
transform 1 0 22272 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_218
timestamp 1621261055
transform 1 0 22080 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_221
timestamp 1621261055
transform 1 0 22368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_229
timestamp 1621261055
transform 1 0 23136 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_237
timestamp 1621261055
transform 1 0 23904 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_245
timestamp 1621261055
transform 1 0 24672 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_253
timestamp 1621261055
transform 1 0 25440 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_261
timestamp 1621261055
transform 1 0 26208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_269
timestamp 1621261055
transform 1 0 26976 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_693
timestamp 1621261055
transform 1 0 27552 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_273
timestamp 1621261055
transform 1 0 27360 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_276
timestamp 1621261055
transform 1 0 27648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_284
timestamp 1621261055
transform 1 0 28416 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_292
timestamp 1621261055
transform 1 0 29184 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_300
timestamp 1621261055
transform 1 0 29952 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_308
timestamp 1621261055
transform 1 0 30720 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_316
timestamp 1621261055
transform 1 0 31488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_324
timestamp 1621261055
transform 1 0 32256 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_694
timestamp 1621261055
transform 1 0 32832 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_328
timestamp 1621261055
transform 1 0 32640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_331
timestamp 1621261055
transform 1 0 32928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_339
timestamp 1621261055
transform 1 0 33696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_347
timestamp 1621261055
transform 1 0 34464 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_355
timestamp 1621261055
transform 1 0 35232 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_363
timestamp 1621261055
transform 1 0 36000 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_371
timestamp 1621261055
transform 1 0 36768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _024_
timestamp 1621261055
transform 1 0 38880 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_695
timestamp 1621261055
transform 1 0 38112 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_379
timestamp 1621261055
transform 1 0 37536 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_383
timestamp 1621261055
transform 1 0 37920 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_49_386
timestamp 1621261055
transform 1 0 38208 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_390
timestamp 1621261055
transform 1 0 38592 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_392
timestamp 1621261055
transform 1 0 38784 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_396
timestamp 1621261055
transform 1 0 39168 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_404
timestamp 1621261055
transform 1 0 39936 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_412
timestamp 1621261055
transform 1 0 40704 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_420
timestamp 1621261055
transform 1 0 41472 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_428
timestamp 1621261055
transform 1 0 42240 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _194_
timestamp 1621261055
transform -1 0 44160 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_696
timestamp 1621261055
transform 1 0 43392 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_224
timestamp 1621261055
transform -1 0 43872 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_49_436
timestamp 1621261055
transform 1 0 43008 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_441
timestamp 1621261055
transform 1 0 43488 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_448
timestamp 1621261055
transform 1 0 44160 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_456
timestamp 1621261055
transform 1 0 44928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_464
timestamp 1621261055
transform 1 0 45696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_472
timestamp 1621261055
transform 1 0 46464 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_480
timestamp 1621261055
transform 1 0 47232 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_697
timestamp 1621261055
transform 1 0 48672 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_488
timestamp 1621261055
transform 1 0 48000 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_492
timestamp 1621261055
transform 1 0 48384 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_494
timestamp 1621261055
transform 1 0 48576 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_496
timestamp 1621261055
transform 1 0 48768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_504
timestamp 1621261055
transform 1 0 49536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_512
timestamp 1621261055
transform 1 0 50304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_520
timestamp 1621261055
transform 1 0 51072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_528
timestamp 1621261055
transform 1 0 51840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_536
timestamp 1621261055
transform 1 0 52608 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_698
timestamp 1621261055
transform 1 0 53952 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_544
timestamp 1621261055
transform 1 0 53376 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_548
timestamp 1621261055
transform 1 0 53760 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_551
timestamp 1621261055
transform 1 0 54048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_559
timestamp 1621261055
transform 1 0 54816 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_567
timestamp 1621261055
transform 1 0 55584 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_575
timestamp 1621261055
transform 1 0 56352 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_583
timestamp 1621261055
transform 1 0 57120 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_591
timestamp 1621261055
transform 1 0 57888 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_99
timestamp 1621261055
transform -1 0 58848 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_595
timestamp 1621261055
transform 1 0 58272 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _002_
timestamp 1621261055
transform 1 0 2400 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_100
timestamp 1621261055
transform 1 0 1152 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_4
timestamp 1621261055
transform 1 0 1536 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_50_12
timestamp 1621261055
transform 1 0 2304 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_16
timestamp 1621261055
transform 1 0 2688 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_24
timestamp 1621261055
transform 1 0 3456 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_699
timestamp 1621261055
transform 1 0 3840 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_29
timestamp 1621261055
transform 1 0 3936 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_37
timestamp 1621261055
transform 1 0 4704 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_45
timestamp 1621261055
transform 1 0 5472 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_53
timestamp 1621261055
transform 1 0 6240 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _057_
timestamp 1621261055
transform 1 0 7104 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_50_61
timestamp 1621261055
transform 1 0 7008 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_65
timestamp 1621261055
transform 1 0 7392 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_73
timestamp 1621261055
transform 1 0 8160 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_81
timestamp 1621261055
transform 1 0 8928 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_700
timestamp 1621261055
transform 1 0 9120 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_84
timestamp 1621261055
transform 1 0 9216 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_92
timestamp 1621261055
transform 1 0 9984 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_100
timestamp 1621261055
transform 1 0 10752 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_108
timestamp 1621261055
transform 1 0 11520 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_116
timestamp 1621261055
transform 1 0 12288 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_124
timestamp 1621261055
transform 1 0 13056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_132
timestamp 1621261055
transform 1 0 13824 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _089_
timestamp 1621261055
transform 1 0 16608 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_701
timestamp 1621261055
transform 1 0 14400 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_151
timestamp 1621261055
transform 1 0 16416 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_136
timestamp 1621261055
transform 1 0 14208 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_139
timestamp 1621261055
transform 1 0 14496 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_147
timestamp 1621261055
transform 1 0 15264 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_155
timestamp 1621261055
transform 1 0 16032 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_164
timestamp 1621261055
transform 1 0 16896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_172
timestamp 1621261055
transform 1 0 17664 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_180
timestamp 1621261055
transform 1 0 18432 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_188
timestamp 1621261055
transform 1 0 19200 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_702
timestamp 1621261055
transform 1 0 19680 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_50_192
timestamp 1621261055
transform 1 0 19584 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_194
timestamp 1621261055
transform 1 0 19776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_202
timestamp 1621261055
transform 1 0 20544 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_210
timestamp 1621261055
transform 1 0 21312 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_218
timestamp 1621261055
transform 1 0 22080 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_226
timestamp 1621261055
transform 1 0 22848 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_234
timestamp 1621261055
transform 1 0 23616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_242
timestamp 1621261055
transform 1 0 24384 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_703
timestamp 1621261055
transform 1 0 24960 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_246
timestamp 1621261055
transform 1 0 24768 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_249
timestamp 1621261055
transform 1 0 25056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_257
timestamp 1621261055
transform 1 0 25824 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_265
timestamp 1621261055
transform 1 0 26592 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_273
timestamp 1621261055
transform 1 0 27360 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_281
timestamp 1621261055
transform 1 0 28128 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_289
timestamp 1621261055
transform 1 0 28896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_297
timestamp 1621261055
transform 1 0 29664 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_704
timestamp 1621261055
transform 1 0 30240 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_301
timestamp 1621261055
transform 1 0 30048 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_304
timestamp 1621261055
transform 1 0 30336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_312
timestamp 1621261055
transform 1 0 31104 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_320
timestamp 1621261055
transform 1 0 31872 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_328
timestamp 1621261055
transform 1 0 32640 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_336
timestamp 1621261055
transform 1 0 33408 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_344
timestamp 1621261055
transform 1 0 34176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_705
timestamp 1621261055
transform 1 0 35520 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_352
timestamp 1621261055
transform 1 0 34944 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_356
timestamp 1621261055
transform 1 0 35328 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_359
timestamp 1621261055
transform 1 0 35616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_367
timestamp 1621261055
transform 1 0 36384 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_375
timestamp 1621261055
transform 1 0 37152 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_383
timestamp 1621261055
transform 1 0 37920 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_391
timestamp 1621261055
transform 1 0 38688 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_399
timestamp 1621261055
transform 1 0 39456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_706
timestamp 1621261055
transform 1 0 40800 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_407
timestamp 1621261055
transform 1 0 40224 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_411
timestamp 1621261055
transform 1 0 40608 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_414
timestamp 1621261055
transform 1 0 40896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_422
timestamp 1621261055
transform 1 0 41664 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_430
timestamp 1621261055
transform 1 0 42432 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_438
timestamp 1621261055
transform 1 0 43200 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_446
timestamp 1621261055
transform 1 0 43968 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_454
timestamp 1621261055
transform 1 0 44736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_707
timestamp 1621261055
transform 1 0 46080 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_462
timestamp 1621261055
transform 1 0 45504 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_466
timestamp 1621261055
transform 1 0 45888 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_469
timestamp 1621261055
transform 1 0 46176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_477
timestamp 1621261055
transform 1 0 46944 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_485
timestamp 1621261055
transform 1 0 47712 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_493
timestamp 1621261055
transform 1 0 48480 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_501
timestamp 1621261055
transform 1 0 49248 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_509
timestamp 1621261055
transform 1 0 50016 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_708
timestamp 1621261055
transform 1 0 51360 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_517
timestamp 1621261055
transform 1 0 50784 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_521
timestamp 1621261055
transform 1 0 51168 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_524
timestamp 1621261055
transform 1 0 51456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_532
timestamp 1621261055
transform 1 0 52224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_540
timestamp 1621261055
transform 1 0 52992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_548
timestamp 1621261055
transform 1 0 53760 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_556
timestamp 1621261055
transform 1 0 54528 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_564
timestamp 1621261055
transform 1 0 55296 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_709
timestamp 1621261055
transform 1 0 56640 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_572
timestamp 1621261055
transform 1 0 56064 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_576
timestamp 1621261055
transform 1 0 56448 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_579
timestamp 1621261055
transform 1 0 56736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_587
timestamp 1621261055
transform 1 0 57504 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_101
timestamp 1621261055
transform -1 0 58848 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_595
timestamp 1621261055
transform 1 0 58272 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_102
timestamp 1621261055
transform 1 0 1152 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_4
timestamp 1621261055
transform 1 0 1536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_12
timestamp 1621261055
transform 1 0 2304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_20
timestamp 1621261055
transform 1 0 3072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _041_
timestamp 1621261055
transform 1 0 4800 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_51_28
timestamp 1621261055
transform 1 0 3840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_36
timestamp 1621261055
transform 1 0 4608 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_41
timestamp 1621261055
transform 1 0 5088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_49
timestamp 1621261055
transform 1 0 5856 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_53
timestamp 1621261055
transform 1 0 6240 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_710
timestamp 1621261055
transform 1 0 6432 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_56
timestamp 1621261055
transform 1 0 6528 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_64
timestamp 1621261055
transform 1 0 7296 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_72
timestamp 1621261055
transform 1 0 8064 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_80
timestamp 1621261055
transform 1 0 8832 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_88
timestamp 1621261055
transform 1 0 9600 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_96
timestamp 1621261055
transform 1 0 10368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_104
timestamp 1621261055
transform 1 0 11136 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_108
timestamp 1621261055
transform 1 0 11520 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_711
timestamp 1621261055
transform 1 0 11712 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_111
timestamp 1621261055
transform 1 0 11808 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_119
timestamp 1621261055
transform 1 0 12576 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_127
timestamp 1621261055
transform 1 0 13344 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_135
timestamp 1621261055
transform 1 0 14112 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_143
timestamp 1621261055
transform 1 0 14880 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_151
timestamp 1621261055
transform 1 0 15648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_159
timestamp 1621261055
transform 1 0 16416 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_712
timestamp 1621261055
transform 1 0 16992 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_163
timestamp 1621261055
transform 1 0 16800 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_166
timestamp 1621261055
transform 1 0 17088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_174
timestamp 1621261055
transform 1 0 17856 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_182
timestamp 1621261055
transform 1 0 18624 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_190
timestamp 1621261055
transform 1 0 19392 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_198
timestamp 1621261055
transform 1 0 20160 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_206
timestamp 1621261055
transform 1 0 20928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_214
timestamp 1621261055
transform 1 0 21696 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_713
timestamp 1621261055
transform 1 0 22272 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_218
timestamp 1621261055
transform 1 0 22080 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_221
timestamp 1621261055
transform 1 0 22368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_229
timestamp 1621261055
transform 1 0 23136 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_237
timestamp 1621261055
transform 1 0 23904 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_245
timestamp 1621261055
transform 1 0 24672 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_253
timestamp 1621261055
transform 1 0 25440 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_261
timestamp 1621261055
transform 1 0 26208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_269
timestamp 1621261055
transform 1 0 26976 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_714
timestamp 1621261055
transform 1 0 27552 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_273
timestamp 1621261055
transform 1 0 27360 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_276
timestamp 1621261055
transform 1 0 27648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_284
timestamp 1621261055
transform 1 0 28416 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_292
timestamp 1621261055
transform 1 0 29184 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_300
timestamp 1621261055
transform 1 0 29952 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_308
timestamp 1621261055
transform 1 0 30720 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_316
timestamp 1621261055
transform 1 0 31488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_324
timestamp 1621261055
transform 1 0 32256 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _159_
timestamp 1621261055
transform 1 0 33888 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_715
timestamp 1621261055
transform 1 0 32832 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_103
timestamp 1621261055
transform 1 0 33696 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_328
timestamp 1621261055
transform 1 0 32640 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_331
timestamp 1621261055
transform 1 0 32928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_344
timestamp 1621261055
transform 1 0 34176 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_352
timestamp 1621261055
transform 1 0 34944 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_360
timestamp 1621261055
transform 1 0 35712 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_368
timestamp 1621261055
transform 1 0 36480 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_376
timestamp 1621261055
transform 1 0 37248 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_716
timestamp 1621261055
transform 1 0 38112 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_51_384
timestamp 1621261055
transform 1 0 38016 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_386
timestamp 1621261055
transform 1 0 38208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_394
timestamp 1621261055
transform 1 0 38976 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_402
timestamp 1621261055
transform 1 0 39744 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_410
timestamp 1621261055
transform 1 0 40512 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_418
timestamp 1621261055
transform 1 0 41280 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_426
timestamp 1621261055
transform 1 0 42048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_717
timestamp 1621261055
transform 1 0 43392 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_434
timestamp 1621261055
transform 1 0 42816 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_438
timestamp 1621261055
transform 1 0 43200 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_441
timestamp 1621261055
transform 1 0 43488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_449
timestamp 1621261055
transform 1 0 44256 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_457
timestamp 1621261055
transform 1 0 45024 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_465
timestamp 1621261055
transform 1 0 45792 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_473
timestamp 1621261055
transform 1 0 46560 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_481
timestamp 1621261055
transform 1 0 47328 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_718
timestamp 1621261055
transform 1 0 48672 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_489
timestamp 1621261055
transform 1 0 48096 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_493
timestamp 1621261055
transform 1 0 48480 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_496
timestamp 1621261055
transform 1 0 48768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_504
timestamp 1621261055
transform 1 0 49536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_512
timestamp 1621261055
transform 1 0 50304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_520
timestamp 1621261055
transform 1 0 51072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_528
timestamp 1621261055
transform 1 0 51840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_536
timestamp 1621261055
transform 1 0 52608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_719
timestamp 1621261055
transform 1 0 53952 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_544
timestamp 1621261055
transform 1 0 53376 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_548
timestamp 1621261055
transform 1 0 53760 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_551
timestamp 1621261055
transform 1 0 54048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_559
timestamp 1621261055
transform 1 0 54816 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_567
timestamp 1621261055
transform 1 0 55584 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_575
timestamp 1621261055
transform 1 0 56352 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_583
timestamp 1621261055
transform 1 0 57120 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_591
timestamp 1621261055
transform 1 0 57888 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_103
timestamp 1621261055
transform -1 0 58848 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_595
timestamp 1621261055
transform 1 0 58272 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_104
timestamp 1621261055
transform 1 0 1152 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_4
timestamp 1621261055
transform 1 0 1536 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_12
timestamp 1621261055
transform 1 0 2304 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_20
timestamp 1621261055
transform 1 0 3072 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_720
timestamp 1621261055
transform 1 0 3840 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_29
timestamp 1621261055
transform 1 0 3936 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_37
timestamp 1621261055
transform 1 0 4704 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_45
timestamp 1621261055
transform 1 0 5472 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_53
timestamp 1621261055
transform 1 0 6240 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_61
timestamp 1621261055
transform 1 0 7008 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_69
timestamp 1621261055
transform 1 0 7776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_77
timestamp 1621261055
transform 1 0 8544 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_81
timestamp 1621261055
transform 1 0 8928 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_88
timestamp 1621261055
transform 1 0 9600 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_52_84
timestamp 1621261055
transform 1 0 9216 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_721
timestamp 1621261055
transform 1 0 9120 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_96
timestamp 1621261055
transform 1 0 10368 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_52_90
timestamp 1621261055
transform 1 0 9792 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_159
timestamp 1621261055
transform 1 0 9888 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _097_
timestamp 1621261055
transform 1 0 10080 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_52_104
timestamp 1621261055
transform 1 0 11136 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _044_
timestamp 1621261055
transform 1 0 11232 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_52_108
timestamp 1621261055
transform 1 0 11520 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_116
timestamp 1621261055
transform 1 0 12288 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_124
timestamp 1621261055
transform 1 0 13056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_132
timestamp 1621261055
transform 1 0 13824 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_722
timestamp 1621261055
transform 1 0 14400 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_136
timestamp 1621261055
transform 1 0 14208 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_139
timestamp 1621261055
transform 1 0 14496 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_147
timestamp 1621261055
transform 1 0 15264 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_155
timestamp 1621261055
transform 1 0 16032 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_163
timestamp 1621261055
transform 1 0 16800 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_171
timestamp 1621261055
transform 1 0 17568 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_179
timestamp 1621261055
transform 1 0 18336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_187
timestamp 1621261055
transform 1 0 19104 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_723
timestamp 1621261055
transform 1 0 19680 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_191
timestamp 1621261055
transform 1 0 19488 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_194
timestamp 1621261055
transform 1 0 19776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_202
timestamp 1621261055
transform 1 0 20544 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_210
timestamp 1621261055
transform 1 0 21312 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_218
timestamp 1621261055
transform 1 0 22080 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_226
timestamp 1621261055
transform 1 0 22848 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_234
timestamp 1621261055
transform 1 0 23616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_242
timestamp 1621261055
transform 1 0 24384 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_724
timestamp 1621261055
transform 1 0 24960 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_246
timestamp 1621261055
transform 1 0 24768 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_249
timestamp 1621261055
transform 1 0 25056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_257
timestamp 1621261055
transform 1 0 25824 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_265
timestamp 1621261055
transform 1 0 26592 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _095_
timestamp 1621261055
transform -1 0 29856 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_155
timestamp 1621261055
transform -1 0 29568 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_273
timestamp 1621261055
transform 1 0 27360 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_281
timestamp 1621261055
transform 1 0 28128 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_289
timestamp 1621261055
transform 1 0 28896 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_52_293
timestamp 1621261055
transform 1 0 29280 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_725
timestamp 1621261055
transform 1 0 30240 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_299
timestamp 1621261055
transform 1 0 29856 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_52_304
timestamp 1621261055
transform 1 0 30336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_312
timestamp 1621261055
transform 1 0 31104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_320
timestamp 1621261055
transform 1 0 31872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_328
timestamp 1621261055
transform 1 0 32640 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_336
timestamp 1621261055
transform 1 0 33408 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_344
timestamp 1621261055
transform 1 0 34176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_726
timestamp 1621261055
transform 1 0 35520 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_352
timestamp 1621261055
transform 1 0 34944 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_356
timestamp 1621261055
transform 1 0 35328 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_359
timestamp 1621261055
transform 1 0 35616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_367
timestamp 1621261055
transform 1 0 36384 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_375
timestamp 1621261055
transform 1 0 37152 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_383
timestamp 1621261055
transform 1 0 37920 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_391
timestamp 1621261055
transform 1 0 38688 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_399
timestamp 1621261055
transform 1 0 39456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_727
timestamp 1621261055
transform 1 0 40800 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_407
timestamp 1621261055
transform 1 0 40224 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_411
timestamp 1621261055
transform 1 0 40608 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_414
timestamp 1621261055
transform 1 0 40896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_422
timestamp 1621261055
transform 1 0 41664 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_430
timestamp 1621261055
transform 1 0 42432 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_438
timestamp 1621261055
transform 1 0 43200 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_446
timestamp 1621261055
transform 1 0 43968 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_454
timestamp 1621261055
transform 1 0 44736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_728
timestamp 1621261055
transform 1 0 46080 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_462
timestamp 1621261055
transform 1 0 45504 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_466
timestamp 1621261055
transform 1 0 45888 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_469
timestamp 1621261055
transform 1 0 46176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_477
timestamp 1621261055
transform 1 0 46944 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_485
timestamp 1621261055
transform 1 0 47712 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_493
timestamp 1621261055
transform 1 0 48480 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_501
timestamp 1621261055
transform 1 0 49248 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_509
timestamp 1621261055
transform 1 0 50016 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_729
timestamp 1621261055
transform 1 0 51360 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_517
timestamp 1621261055
transform 1 0 50784 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_521
timestamp 1621261055
transform 1 0 51168 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_524
timestamp 1621261055
transform 1 0 51456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_532
timestamp 1621261055
transform 1 0 52224 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_540
timestamp 1621261055
transform 1 0 52992 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_548
timestamp 1621261055
transform 1 0 53760 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_556
timestamp 1621261055
transform 1 0 54528 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_564
timestamp 1621261055
transform 1 0 55296 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_730
timestamp 1621261055
transform 1 0 56640 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_52_572
timestamp 1621261055
transform 1 0 56064 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_576
timestamp 1621261055
transform 1 0 56448 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_579
timestamp 1621261055
transform 1 0 56736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_587
timestamp 1621261055
transform 1 0 57504 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_105
timestamp 1621261055
transform -1 0 58848 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_595
timestamp 1621261055
transform 1 0 58272 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_106
timestamp 1621261055
transform 1 0 1152 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_4
timestamp 1621261055
transform 1 0 1536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_12
timestamp 1621261055
transform 1 0 2304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_20
timestamp 1621261055
transform 1 0 3072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_28
timestamp 1621261055
transform 1 0 3840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_36
timestamp 1621261055
transform 1 0 4608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_44
timestamp 1621261055
transform 1 0 5376 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_52
timestamp 1621261055
transform 1 0 6144 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_54
timestamp 1621261055
transform 1 0 6336 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_731
timestamp 1621261055
transform 1 0 6432 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_56
timestamp 1621261055
transform 1 0 6528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_64
timestamp 1621261055
transform 1 0 7296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_72
timestamp 1621261055
transform 1 0 8064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_80
timestamp 1621261055
transform 1 0 8832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _188_
timestamp 1621261055
transform -1 0 11136 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_247
timestamp 1621261055
transform -1 0 10848 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_88
timestamp 1621261055
transform 1 0 9600 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_96
timestamp 1621261055
transform 1 0 10368 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_98
timestamp 1621261055
transform 1 0 10560 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_104
timestamp 1621261055
transform 1 0 11136 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_108
timestamp 1621261055
transform 1 0 11520 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _155_
timestamp 1621261055
transform 1 0 12864 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_732
timestamp 1621261055
transform 1 0 11712 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_99
timestamp 1621261055
transform 1 0 12672 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_111
timestamp 1621261055
transform 1 0 11808 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_53_119
timestamp 1621261055
transform 1 0 12576 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_125
timestamp 1621261055
transform 1 0 13152 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_133
timestamp 1621261055
transform 1 0 13920 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_141
timestamp 1621261055
transform 1 0 14688 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_149
timestamp 1621261055
transform 1 0 15456 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_157
timestamp 1621261055
transform 1 0 16224 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_733
timestamp 1621261055
transform 1 0 16992 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_166
timestamp 1621261055
transform 1 0 17088 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_174
timestamp 1621261055
transform 1 0 17856 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_182
timestamp 1621261055
transform 1 0 18624 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_190
timestamp 1621261055
transform 1 0 19392 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_198
timestamp 1621261055
transform 1 0 20160 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_206
timestamp 1621261055
transform 1 0 20928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_214
timestamp 1621261055
transform 1 0 21696 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_734
timestamp 1621261055
transform 1 0 22272 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_218
timestamp 1621261055
transform 1 0 22080 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_221
timestamp 1621261055
transform 1 0 22368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_229
timestamp 1621261055
transform 1 0 23136 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_237
timestamp 1621261055
transform 1 0 23904 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_245
timestamp 1621261055
transform 1 0 24672 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_253
timestamp 1621261055
transform 1 0 25440 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_261
timestamp 1621261055
transform 1 0 26208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_269
timestamp 1621261055
transform 1 0 26976 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_735
timestamp 1621261055
transform 1 0 27552 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_273
timestamp 1621261055
transform 1 0 27360 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_276
timestamp 1621261055
transform 1 0 27648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_284
timestamp 1621261055
transform 1 0 28416 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_292
timestamp 1621261055
transform 1 0 29184 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_300
timestamp 1621261055
transform 1 0 29952 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_308
timestamp 1621261055
transform 1 0 30720 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_316
timestamp 1621261055
transform 1 0 31488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_324
timestamp 1621261055
transform 1 0 32256 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_736
timestamp 1621261055
transform 1 0 32832 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_328
timestamp 1621261055
transform 1 0 32640 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_331
timestamp 1621261055
transform 1 0 32928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_339
timestamp 1621261055
transform 1 0 33696 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_347
timestamp 1621261055
transform 1 0 34464 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_355
timestamp 1621261055
transform 1 0 35232 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_363
timestamp 1621261055
transform 1 0 36000 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_371
timestamp 1621261055
transform 1 0 36768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_737
timestamp 1621261055
transform 1 0 38112 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_379
timestamp 1621261055
transform 1 0 37536 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_383
timestamp 1621261055
transform 1 0 37920 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_386
timestamp 1621261055
transform 1 0 38208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_394
timestamp 1621261055
transform 1 0 38976 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_402
timestamp 1621261055
transform 1 0 39744 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_410
timestamp 1621261055
transform 1 0 40512 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_418
timestamp 1621261055
transform 1 0 41280 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_426
timestamp 1621261055
transform 1 0 42048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_738
timestamp 1621261055
transform 1 0 43392 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_434
timestamp 1621261055
transform 1 0 42816 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_438
timestamp 1621261055
transform 1 0 43200 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_441
timestamp 1621261055
transform 1 0 43488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_449
timestamp 1621261055
transform 1 0 44256 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_457
timestamp 1621261055
transform 1 0 45024 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_465
timestamp 1621261055
transform 1 0 45792 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_473
timestamp 1621261055
transform 1 0 46560 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_481
timestamp 1621261055
transform 1 0 47328 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_739
timestamp 1621261055
transform 1 0 48672 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_489
timestamp 1621261055
transform 1 0 48096 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_493
timestamp 1621261055
transform 1 0 48480 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_496
timestamp 1621261055
transform 1 0 48768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_504
timestamp 1621261055
transform 1 0 49536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_512
timestamp 1621261055
transform 1 0 50304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_520
timestamp 1621261055
transform 1 0 51072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_528
timestamp 1621261055
transform 1 0 51840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_536
timestamp 1621261055
transform 1 0 52608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_740
timestamp 1621261055
transform 1 0 53952 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_544
timestamp 1621261055
transform 1 0 53376 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_548
timestamp 1621261055
transform 1 0 53760 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_551
timestamp 1621261055
transform 1 0 54048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_559
timestamp 1621261055
transform 1 0 54816 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_567
timestamp 1621261055
transform 1 0 55584 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_575
timestamp 1621261055
transform 1 0 56352 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_583
timestamp 1621261055
transform 1 0 57120 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_591
timestamp 1621261055
transform 1 0 57888 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_107
timestamp 1621261055
transform -1 0 58848 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_595
timestamp 1621261055
transform 1 0 58272 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_108
timestamp 1621261055
transform 1 0 1152 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_110
timestamp 1621261055
transform 1 0 1152 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_4
timestamp 1621261055
transform 1 0 1536 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_12
timestamp 1621261055
transform 1 0 2304 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_20
timestamp 1621261055
transform 1 0 3072 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_4
timestamp 1621261055
transform 1 0 1536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_12
timestamp 1621261055
transform 1 0 2304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_20
timestamp 1621261055
transform 1 0 3072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_28
timestamp 1621261055
transform 1 0 3840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_29
timestamp 1621261055
transform 1 0 3936 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_741
timestamp 1621261055
transform 1 0 3840 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_44
timestamp 1621261055
transform 1 0 5376 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_36
timestamp 1621261055
transform 1 0 4608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_37
timestamp 1621261055
transform 1 0 4704 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_52
timestamp 1621261055
transform 1 0 6144 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_53
timestamp 1621261055
transform 1 0 6240 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_45
timestamp 1621261055
transform 1 0 5472 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_55_54
timestamp 1621261055
transform 1 0 6336 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_752
timestamp 1621261055
transform 1 0 6432 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_61
timestamp 1621261055
transform 1 0 7008 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_69
timestamp 1621261055
transform 1 0 7776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_77
timestamp 1621261055
transform 1 0 8544 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_81
timestamp 1621261055
transform 1 0 8928 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_56
timestamp 1621261055
transform 1 0 6528 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_64
timestamp 1621261055
transform 1 0 7296 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_72
timestamp 1621261055
transform 1 0 8064 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_80
timestamp 1621261055
transform 1 0 8832 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_742
timestamp 1621261055
transform 1 0 9120 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_84
timestamp 1621261055
transform 1 0 9216 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_92
timestamp 1621261055
transform 1 0 9984 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_100
timestamp 1621261055
transform 1 0 10752 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_108
timestamp 1621261055
transform 1 0 11520 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_88
timestamp 1621261055
transform 1 0 9600 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_96
timestamp 1621261055
transform 1 0 10368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_104
timestamp 1621261055
transform 1 0 11136 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_108
timestamp 1621261055
transform 1 0 11520 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_111
timestamp 1621261055
transform 1 0 11808 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_114
timestamp 1621261055
transform 1 0 12096 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_112
timestamp 1621261055
transform 1 0 11904 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_128
timestamp 1621261055
transform 1 0 12192 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_753
timestamp 1621261055
transform 1 0 11712 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_119
timestamp 1621261055
transform 1 0 12576 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_120
timestamp 1621261055
transform 1 0 12672 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _177_
timestamp 1621261055
transform 1 0 12384 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_127
timestamp 1621261055
transform 1 0 13344 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_128
timestamp 1621261055
transform 1 0 13440 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_135
timestamp 1621261055
transform 1 0 14112 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_743
timestamp 1621261055
transform 1 0 14400 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_136
timestamp 1621261055
transform 1 0 14208 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_139
timestamp 1621261055
transform 1 0 14496 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_147
timestamp 1621261055
transform 1 0 15264 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_155
timestamp 1621261055
transform 1 0 16032 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_143
timestamp 1621261055
transform 1 0 14880 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_151
timestamp 1621261055
transform 1 0 15648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_159
timestamp 1621261055
transform 1 0 16416 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_754
timestamp 1621261055
transform 1 0 16992 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_163
timestamp 1621261055
transform 1 0 16800 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_171
timestamp 1621261055
transform 1 0 17568 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_179
timestamp 1621261055
transform 1 0 18336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_187
timestamp 1621261055
transform 1 0 19104 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_163
timestamp 1621261055
transform 1 0 16800 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_166
timestamp 1621261055
transform 1 0 17088 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_174
timestamp 1621261055
transform 1 0 17856 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_182
timestamp 1621261055
transform 1 0 18624 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_744
timestamp 1621261055
transform 1 0 19680 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_191
timestamp 1621261055
transform 1 0 19488 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_194
timestamp 1621261055
transform 1 0 19776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_202
timestamp 1621261055
transform 1 0 20544 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_210
timestamp 1621261055
transform 1 0 21312 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_190
timestamp 1621261055
transform 1 0 19392 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_198
timestamp 1621261055
transform 1 0 20160 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_206
timestamp 1621261055
transform 1 0 20928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_214
timestamp 1621261055
transform 1 0 21696 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_221
timestamp 1621261055
transform 1 0 22368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_218
timestamp 1621261055
transform 1 0 22080 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_218
timestamp 1621261055
transform 1 0 22080 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_755
timestamp 1621261055
transform 1 0 22272 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_229
timestamp 1621261055
transform 1 0 23136 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_226
timestamp 1621261055
transform 1 0 22848 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_237
timestamp 1621261055
transform 1 0 23904 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_240
timestamp 1621261055
transform 1 0 24192 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_236
timestamp 1621261055
transform 1 0 23808 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_234
timestamp 1621261055
transform 1 0 23616 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _174_
timestamp 1621261055
transform 1 0 23904 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_745
timestamp 1621261055
transform 1 0 24960 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_249
timestamp 1621261055
transform 1 0 25056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_257
timestamp 1621261055
transform 1 0 25824 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_265
timestamp 1621261055
transform 1 0 26592 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_245
timestamp 1621261055
transform 1 0 24672 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_253
timestamp 1621261055
transform 1 0 25440 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_261
timestamp 1621261055
transform 1 0 26208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_269
timestamp 1621261055
transform 1 0 26976 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_756
timestamp 1621261055
transform 1 0 27552 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_273
timestamp 1621261055
transform 1 0 27360 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_281
timestamp 1621261055
transform 1 0 28128 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_289
timestamp 1621261055
transform 1 0 28896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_297
timestamp 1621261055
transform 1 0 29664 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_273
timestamp 1621261055
transform 1 0 27360 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_276
timestamp 1621261055
transform 1 0 27648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_284
timestamp 1621261055
transform 1 0 28416 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_292
timestamp 1621261055
transform 1 0 29184 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_746
timestamp 1621261055
transform 1 0 30240 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_301
timestamp 1621261055
transform 1 0 30048 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_304
timestamp 1621261055
transform 1 0 30336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_312
timestamp 1621261055
transform 1 0 31104 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_320
timestamp 1621261055
transform 1 0 31872 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_300
timestamp 1621261055
transform 1 0 29952 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_308
timestamp 1621261055
transform 1 0 30720 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_316
timestamp 1621261055
transform 1 0 31488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_324
timestamp 1621261055
transform 1 0 32256 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_757
timestamp 1621261055
transform 1 0 32832 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_328
timestamp 1621261055
transform 1 0 32640 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_336
timestamp 1621261055
transform 1 0 33408 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_344
timestamp 1621261055
transform 1 0 34176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_328
timestamp 1621261055
transform 1 0 32640 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_331
timestamp 1621261055
transform 1 0 32928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_339
timestamp 1621261055
transform 1 0 33696 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_347
timestamp 1621261055
transform 1 0 34464 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_747
timestamp 1621261055
transform 1 0 35520 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_352
timestamp 1621261055
transform 1 0 34944 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_356
timestamp 1621261055
transform 1 0 35328 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_359
timestamp 1621261055
transform 1 0 35616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_367
timestamp 1621261055
transform 1 0 36384 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_375
timestamp 1621261055
transform 1 0 37152 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_355
timestamp 1621261055
transform 1 0 35232 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_363
timestamp 1621261055
transform 1 0 36000 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_371
timestamp 1621261055
transform 1 0 36768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_758
timestamp 1621261055
transform 1 0 38112 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_383
timestamp 1621261055
transform 1 0 37920 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_391
timestamp 1621261055
transform 1 0 38688 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_399
timestamp 1621261055
transform 1 0 39456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_379
timestamp 1621261055
transform 1 0 37536 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_383
timestamp 1621261055
transform 1 0 37920 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_386
timestamp 1621261055
transform 1 0 38208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_394
timestamp 1621261055
transform 1 0 38976 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_402
timestamp 1621261055
transform 1 0 39744 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_748
timestamp 1621261055
transform 1 0 40800 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_407
timestamp 1621261055
transform 1 0 40224 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_411
timestamp 1621261055
transform 1 0 40608 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_414
timestamp 1621261055
transform 1 0 40896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_422
timestamp 1621261055
transform 1 0 41664 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_430
timestamp 1621261055
transform 1 0 42432 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_410
timestamp 1621261055
transform 1 0 40512 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_418
timestamp 1621261055
transform 1 0 41280 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_426
timestamp 1621261055
transform 1 0 42048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_759
timestamp 1621261055
transform 1 0 43392 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_438
timestamp 1621261055
transform 1 0 43200 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_446
timestamp 1621261055
transform 1 0 43968 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_454
timestamp 1621261055
transform 1 0 44736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_434
timestamp 1621261055
transform 1 0 42816 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_438
timestamp 1621261055
transform 1 0 43200 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_441
timestamp 1621261055
transform 1 0 43488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_449
timestamp 1621261055
transform 1 0 44256 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_457
timestamp 1621261055
transform 1 0 45024 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_749
timestamp 1621261055
transform 1 0 46080 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_462
timestamp 1621261055
transform 1 0 45504 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_466
timestamp 1621261055
transform 1 0 45888 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_469
timestamp 1621261055
transform 1 0 46176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_477
timestamp 1621261055
transform 1 0 46944 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_485
timestamp 1621261055
transform 1 0 47712 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_465
timestamp 1621261055
transform 1 0 45792 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_473
timestamp 1621261055
transform 1 0 46560 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_481
timestamp 1621261055
transform 1 0 47328 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_493
timestamp 1621261055
transform 1 0 48480 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_489
timestamp 1621261055
transform 1 0 48096 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_493
timestamp 1621261055
transform 1 0 48480 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_503
timestamp 1621261055
transform 1 0 49440 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_496
timestamp 1621261055
transform 1 0 48768 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_501
timestamp 1621261055
transform 1 0 49248 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_149
timestamp 1621261055
transform -1 0 49152 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_760
timestamp 1621261055
transform 1 0 48672 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _083_
timestamp 1621261055
transform -1 0 49440 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_511
timestamp 1621261055
transform 1 0 50208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_509
timestamp 1621261055
transform 1 0 50016 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_519
timestamp 1621261055
transform 1 0 50976 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_521
timestamp 1621261055
transform 1 0 51168 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_517
timestamp 1621261055
transform 1 0 50784 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_527
timestamp 1621261055
transform 1 0 51744 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_524
timestamp 1621261055
transform 1 0 51456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_750
timestamp 1621261055
transform 1 0 51360 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_535
timestamp 1621261055
transform 1 0 52512 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_538
timestamp 1621261055
transform 1 0 52800 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_532
timestamp 1621261055
transform 1 0 52224 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_243
timestamp 1621261055
transform -1 0 52512 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _208_
timestamp 1621261055
transform -1 0 52800 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_55_549
timestamp 1621261055
transform 1 0 53856 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_547
timestamp 1621261055
transform 1 0 53664 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_543
timestamp 1621261055
transform 1 0 53280 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_546
timestamp 1621261055
transform 1 0 53568 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_551
timestamp 1621261055
transform 1 0 54048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_554
timestamp 1621261055
transform 1 0 54336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_761
timestamp 1621261055
transform 1 0 53952 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_559
timestamp 1621261055
transform 1 0 54816 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_562
timestamp 1621261055
transform 1 0 55104 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_567
timestamp 1621261055
transform 1 0 55584 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_575
timestamp 1621261055
transform 1 0 56352 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_570
timestamp 1621261055
transform 1 0 55872 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_583
timestamp 1621261055
transform 1 0 57120 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_579
timestamp 1621261055
transform 1 0 56736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_751
timestamp 1621261055
transform 1 0 56640 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_55_591
timestamp 1621261055
transform 1 0 57888 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_54_593
timestamp 1621261055
transform 1 0 58080 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_54_589
timestamp 1621261055
transform 1 0 57696 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_587
timestamp 1621261055
transform 1 0 57504 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _039_
timestamp 1621261055
transform 1 0 57792 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_109
timestamp 1621261055
transform -1 0 58848 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_111
timestamp 1621261055
transform -1 0 58848 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_595
timestamp 1621261055
transform 1 0 58272 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _014_
timestamp 1621261055
transform 1 0 2784 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_112
timestamp 1621261055
transform 1 0 1152 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_56_4
timestamp 1621261055
transform 1 0 1536 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_12
timestamp 1621261055
transform 1 0 2304 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_56_16
timestamp 1621261055
transform 1 0 2688 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_20
timestamp 1621261055
transform 1 0 3072 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_762
timestamp 1621261055
transform 1 0 3840 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_29
timestamp 1621261055
transform 1 0 3936 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_37
timestamp 1621261055
transform 1 0 4704 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_45
timestamp 1621261055
transform 1 0 5472 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_53
timestamp 1621261055
transform 1 0 6240 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_61
timestamp 1621261055
transform 1 0 7008 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_69
timestamp 1621261055
transform 1 0 7776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_77
timestamp 1621261055
transform 1 0 8544 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_81
timestamp 1621261055
transform 1 0 8928 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_763
timestamp 1621261055
transform 1 0 9120 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_84
timestamp 1621261055
transform 1 0 9216 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_92
timestamp 1621261055
transform 1 0 9984 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_100
timestamp 1621261055
transform 1 0 10752 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_108
timestamp 1621261055
transform 1 0 11520 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_116
timestamp 1621261055
transform 1 0 12288 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_124
timestamp 1621261055
transform 1 0 13056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_132
timestamp 1621261055
transform 1 0 13824 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_764
timestamp 1621261055
transform 1 0 14400 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_136
timestamp 1621261055
transform 1 0 14208 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_139
timestamp 1621261055
transform 1 0 14496 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_147
timestamp 1621261055
transform 1 0 15264 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_155
timestamp 1621261055
transform 1 0 16032 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_163
timestamp 1621261055
transform 1 0 16800 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_171
timestamp 1621261055
transform 1 0 17568 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_179
timestamp 1621261055
transform 1 0 18336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_187
timestamp 1621261055
transform 1 0 19104 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_765
timestamp 1621261055
transform 1 0 19680 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_191
timestamp 1621261055
transform 1 0 19488 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_194
timestamp 1621261055
transform 1 0 19776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_202
timestamp 1621261055
transform 1 0 20544 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_210
timestamp 1621261055
transform 1 0 21312 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_218
timestamp 1621261055
transform 1 0 22080 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_226
timestamp 1621261055
transform 1 0 22848 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_234
timestamp 1621261055
transform 1 0 23616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_242
timestamp 1621261055
transform 1 0 24384 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_766
timestamp 1621261055
transform 1 0 24960 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_246
timestamp 1621261055
transform 1 0 24768 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_249
timestamp 1621261055
transform 1 0 25056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_257
timestamp 1621261055
transform 1 0 25824 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_265
timestamp 1621261055
transform 1 0 26592 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_273
timestamp 1621261055
transform 1 0 27360 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_281
timestamp 1621261055
transform 1 0 28128 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_289
timestamp 1621261055
transform 1 0 28896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_297
timestamp 1621261055
transform 1 0 29664 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_767
timestamp 1621261055
transform 1 0 30240 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_301
timestamp 1621261055
transform 1 0 30048 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_304
timestamp 1621261055
transform 1 0 30336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_312
timestamp 1621261055
transform 1 0 31104 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_320
timestamp 1621261055
transform 1 0 31872 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _059_
timestamp 1621261055
transform -1 0 33408 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_97
timestamp 1621261055
transform -1 0 33120 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_328
timestamp 1621261055
transform 1 0 32640 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_330
timestamp 1621261055
transform 1 0 32832 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_336
timestamp 1621261055
transform 1 0 33408 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_344
timestamp 1621261055
transform 1 0 34176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_768
timestamp 1621261055
transform 1 0 35520 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_352
timestamp 1621261055
transform 1 0 34944 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_356
timestamp 1621261055
transform 1 0 35328 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_359
timestamp 1621261055
transform 1 0 35616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_367
timestamp 1621261055
transform 1 0 36384 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_375
timestamp 1621261055
transform 1 0 37152 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_383
timestamp 1621261055
transform 1 0 37920 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_391
timestamp 1621261055
transform 1 0 38688 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_399
timestamp 1621261055
transform 1 0 39456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_769
timestamp 1621261055
transform 1 0 40800 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_407
timestamp 1621261055
transform 1 0 40224 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_411
timestamp 1621261055
transform 1 0 40608 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_414
timestamp 1621261055
transform 1 0 40896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_422
timestamp 1621261055
transform 1 0 41664 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_430
timestamp 1621261055
transform 1 0 42432 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_438
timestamp 1621261055
transform 1 0 43200 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_446
timestamp 1621261055
transform 1 0 43968 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_454
timestamp 1621261055
transform 1 0 44736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_770
timestamp 1621261055
transform 1 0 46080 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_462
timestamp 1621261055
transform 1 0 45504 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_466
timestamp 1621261055
transform 1 0 45888 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_469
timestamp 1621261055
transform 1 0 46176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_477
timestamp 1621261055
transform 1 0 46944 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_485
timestamp 1621261055
transform 1 0 47712 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_493
timestamp 1621261055
transform 1 0 48480 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_501
timestamp 1621261055
transform 1 0 49248 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_509
timestamp 1621261055
transform 1 0 50016 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_771
timestamp 1621261055
transform 1 0 51360 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_517
timestamp 1621261055
transform 1 0 50784 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_521
timestamp 1621261055
transform 1 0 51168 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_524
timestamp 1621261055
transform 1 0 51456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_532
timestamp 1621261055
transform 1 0 52224 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_540
timestamp 1621261055
transform 1 0 52992 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_548
timestamp 1621261055
transform 1 0 53760 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_556
timestamp 1621261055
transform 1 0 54528 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_564
timestamp 1621261055
transform 1 0 55296 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_772
timestamp 1621261055
transform 1 0 56640 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_56_572
timestamp 1621261055
transform 1 0 56064 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_576
timestamp 1621261055
transform 1 0 56448 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_579
timestamp 1621261055
transform 1 0 56736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_587
timestamp 1621261055
transform 1 0 57504 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_113
timestamp 1621261055
transform -1 0 58848 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_595
timestamp 1621261055
transform 1 0 58272 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _139_
timestamp 1621261055
transform 1 0 1536 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_114
timestamp 1621261055
transform 1 0 1152 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_199
timestamp 1621261055
transform 1 0 1824 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_9
timestamp 1621261055
transform 1 0 2016 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_17
timestamp 1621261055
transform 1 0 2784 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_25
timestamp 1621261055
transform 1 0 3552 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_33
timestamp 1621261055
transform 1 0 4320 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_41
timestamp 1621261055
transform 1 0 5088 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_49
timestamp 1621261055
transform 1 0 5856 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_53
timestamp 1621261055
transform 1 0 6240 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_773
timestamp 1621261055
transform 1 0 6432 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_56
timestamp 1621261055
transform 1 0 6528 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_64
timestamp 1621261055
transform 1 0 7296 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_72
timestamp 1621261055
transform 1 0 8064 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_80
timestamp 1621261055
transform 1 0 8832 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_88
timestamp 1621261055
transform 1 0 9600 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_96
timestamp 1621261055
transform 1 0 10368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_104
timestamp 1621261055
transform 1 0 11136 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_108
timestamp 1621261055
transform 1 0 11520 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_774
timestamp 1621261055
transform 1 0 11712 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_111
timestamp 1621261055
transform 1 0 11808 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_119
timestamp 1621261055
transform 1 0 12576 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_127
timestamp 1621261055
transform 1 0 13344 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_135
timestamp 1621261055
transform 1 0 14112 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _096_
timestamp 1621261055
transform 1 0 15456 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_157
timestamp 1621261055
transform 1 0 15264 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_57_143
timestamp 1621261055
transform 1 0 14880 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_57_152
timestamp 1621261055
transform 1 0 15744 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_160
timestamp 1621261055
transform 1 0 16512 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _129_
timestamp 1621261055
transform 1 0 17472 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_775
timestamp 1621261055
transform 1 0 16992 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_188
timestamp 1621261055
transform 1 0 17280 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_164
timestamp 1621261055
transform 1 0 16896 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_166
timestamp 1621261055
transform 1 0 17088 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_173
timestamp 1621261055
transform 1 0 17760 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_181
timestamp 1621261055
transform 1 0 18528 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_189
timestamp 1621261055
transform 1 0 19296 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_197
timestamp 1621261055
transform 1 0 20064 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_205
timestamp 1621261055
transform 1 0 20832 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_213
timestamp 1621261055
transform 1 0 21600 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_776
timestamp 1621261055
transform 1 0 22272 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_217
timestamp 1621261055
transform 1 0 21984 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_219
timestamp 1621261055
transform 1 0 22176 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_221
timestamp 1621261055
transform 1 0 22368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_229
timestamp 1621261055
transform 1 0 23136 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_237
timestamp 1621261055
transform 1 0 23904 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_245
timestamp 1621261055
transform 1 0 24672 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_253
timestamp 1621261055
transform 1 0 25440 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_261
timestamp 1621261055
transform 1 0 26208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_269
timestamp 1621261055
transform 1 0 26976 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_777
timestamp 1621261055
transform 1 0 27552 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_273
timestamp 1621261055
transform 1 0 27360 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_276
timestamp 1621261055
transform 1 0 27648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_284
timestamp 1621261055
transform 1 0 28416 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_292
timestamp 1621261055
transform 1 0 29184 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_300
timestamp 1621261055
transform 1 0 29952 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_308
timestamp 1621261055
transform 1 0 30720 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_316
timestamp 1621261055
transform 1 0 31488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_324
timestamp 1621261055
transform 1 0 32256 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_778
timestamp 1621261055
transform 1 0 32832 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_328
timestamp 1621261055
transform 1 0 32640 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_331
timestamp 1621261055
transform 1 0 32928 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_339
timestamp 1621261055
transform 1 0 33696 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_347
timestamp 1621261055
transform 1 0 34464 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_355
timestamp 1621261055
transform 1 0 35232 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_363
timestamp 1621261055
transform 1 0 36000 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_371
timestamp 1621261055
transform 1 0 36768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_779
timestamp 1621261055
transform 1 0 38112 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_379
timestamp 1621261055
transform 1 0 37536 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_383
timestamp 1621261055
transform 1 0 37920 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_386
timestamp 1621261055
transform 1 0 38208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_394
timestamp 1621261055
transform 1 0 38976 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_402
timestamp 1621261055
transform 1 0 39744 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_410
timestamp 1621261055
transform 1 0 40512 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_418
timestamp 1621261055
transform 1 0 41280 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_426
timestamp 1621261055
transform 1 0 42048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_780
timestamp 1621261055
transform 1 0 43392 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_434
timestamp 1621261055
transform 1 0 42816 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_438
timestamp 1621261055
transform 1 0 43200 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_441
timestamp 1621261055
transform 1 0 43488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_449
timestamp 1621261055
transform 1 0 44256 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_457
timestamp 1621261055
transform 1 0 45024 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_465
timestamp 1621261055
transform 1 0 45792 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_473
timestamp 1621261055
transform 1 0 46560 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_481
timestamp 1621261055
transform 1 0 47328 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_781
timestamp 1621261055
transform 1 0 48672 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_489
timestamp 1621261055
transform 1 0 48096 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_493
timestamp 1621261055
transform 1 0 48480 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_496
timestamp 1621261055
transform 1 0 48768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_504
timestamp 1621261055
transform 1 0 49536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_512
timestamp 1621261055
transform 1 0 50304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_520
timestamp 1621261055
transform 1 0 51072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_528
timestamp 1621261055
transform 1 0 51840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_536
timestamp 1621261055
transform 1 0 52608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_782
timestamp 1621261055
transform 1 0 53952 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_544
timestamp 1621261055
transform 1 0 53376 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_548
timestamp 1621261055
transform 1 0 53760 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_551
timestamp 1621261055
transform 1 0 54048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_559
timestamp 1621261055
transform 1 0 54816 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_567
timestamp 1621261055
transform 1 0 55584 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_575
timestamp 1621261055
transform 1 0 56352 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_583
timestamp 1621261055
transform 1 0 57120 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_591
timestamp 1621261055
transform 1 0 57888 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_115
timestamp 1621261055
transform -1 0 58848 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_595
timestamp 1621261055
transform 1 0 58272 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_116
timestamp 1621261055
transform 1 0 1152 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_58_4
timestamp 1621261055
transform 1 0 1536 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_12
timestamp 1621261055
transform 1 0 2304 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_20
timestamp 1621261055
transform 1 0 3072 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_783
timestamp 1621261055
transform 1 0 3840 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_29
timestamp 1621261055
transform 1 0 3936 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_37
timestamp 1621261055
transform 1 0 4704 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_45
timestamp 1621261055
transform 1 0 5472 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_53
timestamp 1621261055
transform 1 0 6240 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_61
timestamp 1621261055
transform 1 0 7008 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_69
timestamp 1621261055
transform 1 0 7776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_77
timestamp 1621261055
transform 1 0 8544 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_81
timestamp 1621261055
transform 1 0 8928 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_784
timestamp 1621261055
transform 1 0 9120 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_84
timestamp 1621261055
transform 1 0 9216 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_92
timestamp 1621261055
transform 1 0 9984 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_100
timestamp 1621261055
transform 1 0 10752 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_108
timestamp 1621261055
transform 1 0 11520 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_116
timestamp 1621261055
transform 1 0 12288 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_124
timestamp 1621261055
transform 1 0 13056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_132
timestamp 1621261055
transform 1 0 13824 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_785
timestamp 1621261055
transform 1 0 14400 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_136
timestamp 1621261055
transform 1 0 14208 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_139
timestamp 1621261055
transform 1 0 14496 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_147
timestamp 1621261055
transform 1 0 15264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_155
timestamp 1621261055
transform 1 0 16032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_163
timestamp 1621261055
transform 1 0 16800 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_171
timestamp 1621261055
transform 1 0 17568 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_179
timestamp 1621261055
transform 1 0 18336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_187
timestamp 1621261055
transform 1 0 19104 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_786
timestamp 1621261055
transform 1 0 19680 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_191
timestamp 1621261055
transform 1 0 19488 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_194
timestamp 1621261055
transform 1 0 19776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_202
timestamp 1621261055
transform 1 0 20544 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_210
timestamp 1621261055
transform 1 0 21312 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_218
timestamp 1621261055
transform 1 0 22080 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_226
timestamp 1621261055
transform 1 0 22848 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_234
timestamp 1621261055
transform 1 0 23616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_242
timestamp 1621261055
transform 1 0 24384 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _143_
timestamp 1621261055
transform 1 0 25440 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_787
timestamp 1621261055
transform 1 0 24960 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_205
timestamp 1621261055
transform 1 0 25248 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_246
timestamp 1621261055
transform 1 0 24768 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_249
timestamp 1621261055
transform 1 0 25056 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_256
timestamp 1621261055
transform 1 0 25728 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_264
timestamp 1621261055
transform 1 0 26496 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_272
timestamp 1621261055
transform 1 0 27264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_280
timestamp 1621261055
transform 1 0 28032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_288
timestamp 1621261055
transform 1 0 28800 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_296
timestamp 1621261055
transform 1 0 29568 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_788
timestamp 1621261055
transform 1 0 30240 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_300
timestamp 1621261055
transform 1 0 29952 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_302
timestamp 1621261055
transform 1 0 30144 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_304
timestamp 1621261055
transform 1 0 30336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_312
timestamp 1621261055
transform 1 0 31104 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_320
timestamp 1621261055
transform 1 0 31872 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_328
timestamp 1621261055
transform 1 0 32640 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_336
timestamp 1621261055
transform 1 0 33408 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_344
timestamp 1621261055
transform 1 0 34176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_789
timestamp 1621261055
transform 1 0 35520 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_352
timestamp 1621261055
transform 1 0 34944 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_356
timestamp 1621261055
transform 1 0 35328 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_359
timestamp 1621261055
transform 1 0 35616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_367
timestamp 1621261055
transform 1 0 36384 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_375
timestamp 1621261055
transform 1 0 37152 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_383
timestamp 1621261055
transform 1 0 37920 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_391
timestamp 1621261055
transform 1 0 38688 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_399
timestamp 1621261055
transform 1 0 39456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_790
timestamp 1621261055
transform 1 0 40800 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_407
timestamp 1621261055
transform 1 0 40224 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_411
timestamp 1621261055
transform 1 0 40608 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_414
timestamp 1621261055
transform 1 0 40896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_422
timestamp 1621261055
transform 1 0 41664 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_430
timestamp 1621261055
transform 1 0 42432 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_438
timestamp 1621261055
transform 1 0 43200 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_446
timestamp 1621261055
transform 1 0 43968 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_454
timestamp 1621261055
transform 1 0 44736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_791
timestamp 1621261055
transform 1 0 46080 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_462
timestamp 1621261055
transform 1 0 45504 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_466
timestamp 1621261055
transform 1 0 45888 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_469
timestamp 1621261055
transform 1 0 46176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_477
timestamp 1621261055
transform 1 0 46944 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_485
timestamp 1621261055
transform 1 0 47712 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _042_
timestamp 1621261055
transform 1 0 48096 0 -1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_58_492
timestamp 1621261055
transform 1 0 48384 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_500
timestamp 1621261055
transform 1 0 49152 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_508
timestamp 1621261055
transform 1 0 49920 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_792
timestamp 1621261055
transform 1 0 51360 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_516
timestamp 1621261055
transform 1 0 50688 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_520
timestamp 1621261055
transform 1 0 51072 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_58_522
timestamp 1621261055
transform 1 0 51264 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_524
timestamp 1621261055
transform 1 0 51456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_532
timestamp 1621261055
transform 1 0 52224 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_540
timestamp 1621261055
transform 1 0 52992 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_548
timestamp 1621261055
transform 1 0 53760 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_556
timestamp 1621261055
transform 1 0 54528 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_564
timestamp 1621261055
transform 1 0 55296 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_793
timestamp 1621261055
transform 1 0 56640 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_58_572
timestamp 1621261055
transform 1 0 56064 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_576
timestamp 1621261055
transform 1 0 56448 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_579
timestamp 1621261055
transform 1 0 56736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_587
timestamp 1621261055
transform 1 0 57504 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_117
timestamp 1621261055
transform -1 0 58848 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_595
timestamp 1621261055
transform 1 0 58272 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_118
timestamp 1621261055
transform 1 0 1152 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_4
timestamp 1621261055
transform 1 0 1536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_12
timestamp 1621261055
transform 1 0 2304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_20
timestamp 1621261055
transform 1 0 3072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_28
timestamp 1621261055
transform 1 0 3840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_36
timestamp 1621261055
transform 1 0 4608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_44
timestamp 1621261055
transform 1 0 5376 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_52
timestamp 1621261055
transform 1 0 6144 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_54
timestamp 1621261055
transform 1 0 6336 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_794
timestamp 1621261055
transform 1 0 6432 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_56
timestamp 1621261055
transform 1 0 6528 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_64
timestamp 1621261055
transform 1 0 7296 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_72
timestamp 1621261055
transform 1 0 8064 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_80
timestamp 1621261055
transform 1 0 8832 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_88
timestamp 1621261055
transform 1 0 9600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_96
timestamp 1621261055
transform 1 0 10368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_104
timestamp 1621261055
transform 1 0 11136 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_108
timestamp 1621261055
transform 1 0 11520 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_795
timestamp 1621261055
transform 1 0 11712 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_111
timestamp 1621261055
transform 1 0 11808 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_119
timestamp 1621261055
transform 1 0 12576 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_127
timestamp 1621261055
transform 1 0 13344 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_135
timestamp 1621261055
transform 1 0 14112 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_143
timestamp 1621261055
transform 1 0 14880 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_151
timestamp 1621261055
transform 1 0 15648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_159
timestamp 1621261055
transform 1 0 16416 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_796
timestamp 1621261055
transform 1 0 16992 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_163
timestamp 1621261055
transform 1 0 16800 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_166
timestamp 1621261055
transform 1 0 17088 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_174
timestamp 1621261055
transform 1 0 17856 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_182
timestamp 1621261055
transform 1 0 18624 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_190
timestamp 1621261055
transform 1 0 19392 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_198
timestamp 1621261055
transform 1 0 20160 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_206
timestamp 1621261055
transform 1 0 20928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_214
timestamp 1621261055
transform 1 0 21696 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_797
timestamp 1621261055
transform 1 0 22272 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_218
timestamp 1621261055
transform 1 0 22080 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_221
timestamp 1621261055
transform 1 0 22368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_229
timestamp 1621261055
transform 1 0 23136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_237
timestamp 1621261055
transform 1 0 23904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_245
timestamp 1621261055
transform 1 0 24672 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_253
timestamp 1621261055
transform 1 0 25440 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_261
timestamp 1621261055
transform 1 0 26208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_269
timestamp 1621261055
transform 1 0 26976 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_798
timestamp 1621261055
transform 1 0 27552 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_273
timestamp 1621261055
transform 1 0 27360 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_276
timestamp 1621261055
transform 1 0 27648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_284
timestamp 1621261055
transform 1 0 28416 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_292
timestamp 1621261055
transform 1 0 29184 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _023_
timestamp 1621261055
transform 1 0 30912 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_59_300
timestamp 1621261055
transform 1 0 29952 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_308
timestamp 1621261055
transform 1 0 30720 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_313
timestamp 1621261055
transform 1 0 31200 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_321
timestamp 1621261055
transform 1 0 31968 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _123_
timestamp 1621261055
transform 1 0 33312 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_799
timestamp 1621261055
transform 1 0 32832 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_182
timestamp 1621261055
transform 1 0 33120 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_329
timestamp 1621261055
transform 1 0 32736 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_331
timestamp 1621261055
transform 1 0 32928 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_338
timestamp 1621261055
transform 1 0 33600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_346
timestamp 1621261055
transform 1 0 34368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_354
timestamp 1621261055
transform 1 0 35136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_362
timestamp 1621261055
transform 1 0 35904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_370
timestamp 1621261055
transform 1 0 36672 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_378
timestamp 1621261055
transform 1 0 37440 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_800
timestamp 1621261055
transform 1 0 38112 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_382
timestamp 1621261055
transform 1 0 37824 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_384
timestamp 1621261055
transform 1 0 38016 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_386
timestamp 1621261055
transform 1 0 38208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_394
timestamp 1621261055
transform 1 0 38976 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_402
timestamp 1621261055
transform 1 0 39744 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _017_
timestamp 1621261055
transform 1 0 40128 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_59_409
timestamp 1621261055
transform 1 0 40416 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_417
timestamp 1621261055
transform 1 0 41184 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_425
timestamp 1621261055
transform 1 0 41952 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_801
timestamp 1621261055
transform 1 0 43392 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_433
timestamp 1621261055
transform 1 0 42720 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_437
timestamp 1621261055
transform 1 0 43104 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_439
timestamp 1621261055
transform 1 0 43296 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_441
timestamp 1621261055
transform 1 0 43488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_449
timestamp 1621261055
transform 1 0 44256 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_457
timestamp 1621261055
transform 1 0 45024 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _193_
timestamp 1621261055
transform -1 0 46752 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_222
timestamp 1621261055
transform -1 0 46464 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_59_465
timestamp 1621261055
transform 1 0 45792 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_59_469
timestamp 1621261055
transform 1 0 46176 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_475
timestamp 1621261055
transform 1 0 46752 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_483
timestamp 1621261055
transform 1 0 47520 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_802
timestamp 1621261055
transform 1 0 48672 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_491
timestamp 1621261055
transform 1 0 48288 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_496
timestamp 1621261055
transform 1 0 48768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_504
timestamp 1621261055
transform 1 0 49536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_512
timestamp 1621261055
transform 1 0 50304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_520
timestamp 1621261055
transform 1 0 51072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_528
timestamp 1621261055
transform 1 0 51840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_536
timestamp 1621261055
transform 1 0 52608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_803
timestamp 1621261055
transform 1 0 53952 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_544
timestamp 1621261055
transform 1 0 53376 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_548
timestamp 1621261055
transform 1 0 53760 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_551
timestamp 1621261055
transform 1 0 54048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_559
timestamp 1621261055
transform 1 0 54816 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_567
timestamp 1621261055
transform 1 0 55584 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_575
timestamp 1621261055
transform 1 0 56352 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_583
timestamp 1621261055
transform 1 0 57120 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_591
timestamp 1621261055
transform 1 0 57888 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_119
timestamp 1621261055
transform -1 0 58848 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_595
timestamp 1621261055
transform 1 0 58272 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _182_
timestamp 1621261055
transform -1 0 2592 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_120
timestamp 1621261055
transform 1 0 1152 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_218
timestamp 1621261055
transform -1 0 2304 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_60_4
timestamp 1621261055
transform 1 0 1536 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_8
timestamp 1621261055
transform 1 0 1920 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_15
timestamp 1621261055
transform 1 0 2592 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_23
timestamp 1621261055
transform 1 0 3360 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_60_27
timestamp 1621261055
transform 1 0 3744 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_804
timestamp 1621261055
transform 1 0 3840 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_29
timestamp 1621261055
transform 1 0 3936 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_37
timestamp 1621261055
transform 1 0 4704 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_45
timestamp 1621261055
transform 1 0 5472 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_53
timestamp 1621261055
transform 1 0 6240 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_61
timestamp 1621261055
transform 1 0 7008 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_69
timestamp 1621261055
transform 1 0 7776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_77
timestamp 1621261055
transform 1 0 8544 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_81
timestamp 1621261055
transform 1 0 8928 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_805
timestamp 1621261055
transform 1 0 9120 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_84
timestamp 1621261055
transform 1 0 9216 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_92
timestamp 1621261055
transform 1 0 9984 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_100
timestamp 1621261055
transform 1 0 10752 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_108
timestamp 1621261055
transform 1 0 11520 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_116
timestamp 1621261055
transform 1 0 12288 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_124
timestamp 1621261055
transform 1 0 13056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_132
timestamp 1621261055
transform 1 0 13824 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_806
timestamp 1621261055
transform 1 0 14400 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_136
timestamp 1621261055
transform 1 0 14208 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_139
timestamp 1621261055
transform 1 0 14496 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_147
timestamp 1621261055
transform 1 0 15264 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_155
timestamp 1621261055
transform 1 0 16032 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_163
timestamp 1621261055
transform 1 0 16800 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_171
timestamp 1621261055
transform 1 0 17568 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_179
timestamp 1621261055
transform 1 0 18336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_187
timestamp 1621261055
transform 1 0 19104 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_807
timestamp 1621261055
transform 1 0 19680 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_191
timestamp 1621261055
transform 1 0 19488 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_194
timestamp 1621261055
transform 1 0 19776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_202
timestamp 1621261055
transform 1 0 20544 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_210
timestamp 1621261055
transform 1 0 21312 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_218
timestamp 1621261055
transform 1 0 22080 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_226
timestamp 1621261055
transform 1 0 22848 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_234
timestamp 1621261055
transform 1 0 23616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_242
timestamp 1621261055
transform 1 0 24384 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_808
timestamp 1621261055
transform 1 0 24960 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_246
timestamp 1621261055
transform 1 0 24768 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_249
timestamp 1621261055
transform 1 0 25056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_257
timestamp 1621261055
transform 1 0 25824 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_265
timestamp 1621261055
transform 1 0 26592 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_273
timestamp 1621261055
transform 1 0 27360 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_281
timestamp 1621261055
transform 1 0 28128 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_289
timestamp 1621261055
transform 1 0 28896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_297
timestamp 1621261055
transform 1 0 29664 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_809
timestamp 1621261055
transform 1 0 30240 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_301
timestamp 1621261055
transform 1 0 30048 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_304
timestamp 1621261055
transform 1 0 30336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_312
timestamp 1621261055
transform 1 0 31104 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_320
timestamp 1621261055
transform 1 0 31872 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_328
timestamp 1621261055
transform 1 0 32640 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_336
timestamp 1621261055
transform 1 0 33408 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_344
timestamp 1621261055
transform 1 0 34176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_810
timestamp 1621261055
transform 1 0 35520 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_352
timestamp 1621261055
transform 1 0 34944 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_356
timestamp 1621261055
transform 1 0 35328 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_359
timestamp 1621261055
transform 1 0 35616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_367
timestamp 1621261055
transform 1 0 36384 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_375
timestamp 1621261055
transform 1 0 37152 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_383
timestamp 1621261055
transform 1 0 37920 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_391
timestamp 1621261055
transform 1 0 38688 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_399
timestamp 1621261055
transform 1 0 39456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_811
timestamp 1621261055
transform 1 0 40800 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_407
timestamp 1621261055
transform 1 0 40224 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_411
timestamp 1621261055
transform 1 0 40608 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_414
timestamp 1621261055
transform 1 0 40896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_422
timestamp 1621261055
transform 1 0 41664 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_430
timestamp 1621261055
transform 1 0 42432 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_438
timestamp 1621261055
transform 1 0 43200 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_446
timestamp 1621261055
transform 1 0 43968 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_454
timestamp 1621261055
transform 1 0 44736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_812
timestamp 1621261055
transform 1 0 46080 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_462
timestamp 1621261055
transform 1 0 45504 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_466
timestamp 1621261055
transform 1 0 45888 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_469
timestamp 1621261055
transform 1 0 46176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_477
timestamp 1621261055
transform 1 0 46944 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_485
timestamp 1621261055
transform 1 0 47712 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_493
timestamp 1621261055
transform 1 0 48480 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_501
timestamp 1621261055
transform 1 0 49248 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_509
timestamp 1621261055
transform 1 0 50016 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_813
timestamp 1621261055
transform 1 0 51360 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_517
timestamp 1621261055
transform 1 0 50784 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_521
timestamp 1621261055
transform 1 0 51168 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_524
timestamp 1621261055
transform 1 0 51456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_532
timestamp 1621261055
transform 1 0 52224 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_540
timestamp 1621261055
transform 1 0 52992 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_548
timestamp 1621261055
transform 1 0 53760 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_556
timestamp 1621261055
transform 1 0 54528 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_564
timestamp 1621261055
transform 1 0 55296 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_814
timestamp 1621261055
transform 1 0 56640 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_60_572
timestamp 1621261055
transform 1 0 56064 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_576
timestamp 1621261055
transform 1 0 56448 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_579
timestamp 1621261055
transform 1 0 56736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_587
timestamp 1621261055
transform 1 0 57504 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_121
timestamp 1621261055
transform -1 0 58848 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_595
timestamp 1621261055
transform 1 0 58272 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_122
timestamp 1621261055
transform 1 0 1152 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_124
timestamp 1621261055
transform 1 0 1152 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_4
timestamp 1621261055
transform 1 0 1536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_12
timestamp 1621261055
transform 1 0 2304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_20
timestamp 1621261055
transform 1 0 3072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_4
timestamp 1621261055
transform 1 0 1536 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_12
timestamp 1621261055
transform 1 0 2304 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_20
timestamp 1621261055
transform 1 0 3072 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_29
timestamp 1621261055
transform 1 0 3936 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_28
timestamp 1621261055
transform 1 0 3840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_825
timestamp 1621261055
transform 1 0 3840 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_37
timestamp 1621261055
transform 1 0 4704 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_44
timestamp 1621261055
transform 1 0 5376 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_36
timestamp 1621261055
transform 1 0 4608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_53
timestamp 1621261055
transform 1 0 6240 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_45
timestamp 1621261055
transform 1 0 5472 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_52
timestamp 1621261055
transform 1 0 6144 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_61_54
timestamp 1621261055
transform 1 0 6336 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_815
timestamp 1621261055
transform 1 0 6432 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_56
timestamp 1621261055
transform 1 0 6528 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_64
timestamp 1621261055
transform 1 0 7296 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_72
timestamp 1621261055
transform 1 0 8064 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_80
timestamp 1621261055
transform 1 0 8832 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_61
timestamp 1621261055
transform 1 0 7008 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_69
timestamp 1621261055
transform 1 0 7776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_77
timestamp 1621261055
transform 1 0 8544 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_81
timestamp 1621261055
transform 1 0 8928 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_826
timestamp 1621261055
transform 1 0 9120 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_88
timestamp 1621261055
transform 1 0 9600 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_96
timestamp 1621261055
transform 1 0 10368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_104
timestamp 1621261055
transform 1 0 11136 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_108
timestamp 1621261055
transform 1 0 11520 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_84
timestamp 1621261055
transform 1 0 9216 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_92
timestamp 1621261055
transform 1 0 9984 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_100
timestamp 1621261055
transform 1 0 10752 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_108
timestamp 1621261055
transform 1 0 11520 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_114
timestamp 1621261055
transform 1 0 12096 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_62_110
timestamp 1621261055
transform 1 0 11712 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_111
timestamp 1621261055
transform 1 0 11808 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_816
timestamp 1621261055
transform 1 0 11712 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _025_
timestamp 1621261055
transform 1 0 11808 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_122
timestamp 1621261055
transform 1 0 12864 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_119
timestamp 1621261055
transform 1 0 12576 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_130
timestamp 1621261055
transform 1 0 13632 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_127
timestamp 1621261055
transform 1 0 13344 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_135
timestamp 1621261055
transform 1 0 14112 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_827
timestamp 1621261055
transform 1 0 14400 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_143
timestamp 1621261055
transform 1 0 14880 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_151
timestamp 1621261055
transform 1 0 15648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_159
timestamp 1621261055
transform 1 0 16416 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_139
timestamp 1621261055
transform 1 0 14496 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_147
timestamp 1621261055
transform 1 0 15264 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_155
timestamp 1621261055
transform 1 0 16032 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_62_165
timestamp 1621261055
transform 1 0 16992 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_163
timestamp 1621261055
transform 1 0 16800 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_166
timestamp 1621261055
transform 1 0 17088 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_163
timestamp 1621261055
transform 1 0 16800 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_233
timestamp 1621261055
transform -1 0 17280 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_817
timestamp 1621261055
transform 1 0 16992 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _202_
timestamp 1621261055
transform -1 0 17568 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_179
timestamp 1621261055
transform 1 0 18336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_171
timestamp 1621261055
transform 1 0 17568 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_174
timestamp 1621261055
transform 1 0 17856 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_187
timestamp 1621261055
transform 1 0 19104 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_182
timestamp 1621261055
transform 1 0 18624 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_194
timestamp 1621261055
transform 1 0 19776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_191
timestamp 1621261055
transform 1 0 19488 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_190
timestamp 1621261055
transform 1 0 19392 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_828
timestamp 1621261055
transform 1 0 19680 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_202
timestamp 1621261055
transform 1 0 20544 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_206
timestamp 1621261055
transform 1 0 20928 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_198
timestamp 1621261055
transform 1 0 20160 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_210
timestamp 1621261055
transform 1 0 21312 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_210
timestamp 1621261055
transform 1 0 21312 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_239
timestamp 1621261055
transform -1 0 21600 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _206_
timestamp 1621261055
transform -1 0 21888 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_61_216
timestamp 1621261055
transform 1 0 21888 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_818
timestamp 1621261055
transform 1 0 22272 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_221
timestamp 1621261055
transform 1 0 22368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_229
timestamp 1621261055
transform 1 0 23136 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_237
timestamp 1621261055
transform 1 0 23904 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_218
timestamp 1621261055
transform 1 0 22080 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_226
timestamp 1621261055
transform 1 0 22848 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_234
timestamp 1621261055
transform 1 0 23616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_242
timestamp 1621261055
transform 1 0 24384 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_829
timestamp 1621261055
transform 1 0 24960 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_245
timestamp 1621261055
transform 1 0 24672 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_253
timestamp 1621261055
transform 1 0 25440 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_261
timestamp 1621261055
transform 1 0 26208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_269
timestamp 1621261055
transform 1 0 26976 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_246
timestamp 1621261055
transform 1 0 24768 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_249
timestamp 1621261055
transform 1 0 25056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_257
timestamp 1621261055
transform 1 0 25824 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_265
timestamp 1621261055
transform 1 0 26592 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_819
timestamp 1621261055
transform 1 0 27552 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_273
timestamp 1621261055
transform 1 0 27360 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_276
timestamp 1621261055
transform 1 0 27648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_284
timestamp 1621261055
transform 1 0 28416 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_292
timestamp 1621261055
transform 1 0 29184 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_273
timestamp 1621261055
transform 1 0 27360 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_281
timestamp 1621261055
transform 1 0 28128 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_289
timestamp 1621261055
transform 1 0 28896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_297
timestamp 1621261055
transform 1 0 29664 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_830
timestamp 1621261055
transform 1 0 30240 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_300
timestamp 1621261055
transform 1 0 29952 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_308
timestamp 1621261055
transform 1 0 30720 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_316
timestamp 1621261055
transform 1 0 31488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_324
timestamp 1621261055
transform 1 0 32256 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_301
timestamp 1621261055
transform 1 0 30048 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_304
timestamp 1621261055
transform 1 0 30336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_312
timestamp 1621261055
transform 1 0 31104 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_320
timestamp 1621261055
transform 1 0 31872 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_820
timestamp 1621261055
transform 1 0 32832 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_328
timestamp 1621261055
transform 1 0 32640 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_331
timestamp 1621261055
transform 1 0 32928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_339
timestamp 1621261055
transform 1 0 33696 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_347
timestamp 1621261055
transform 1 0 34464 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_328
timestamp 1621261055
transform 1 0 32640 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_336
timestamp 1621261055
transform 1 0 33408 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_344
timestamp 1621261055
transform 1 0 34176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_831
timestamp 1621261055
transform 1 0 35520 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_355
timestamp 1621261055
transform 1 0 35232 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_363
timestamp 1621261055
transform 1 0 36000 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_371
timestamp 1621261055
transform 1 0 36768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_352
timestamp 1621261055
transform 1 0 34944 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_356
timestamp 1621261055
transform 1 0 35328 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_359
timestamp 1621261055
transform 1 0 35616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_367
timestamp 1621261055
transform 1 0 36384 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_375
timestamp 1621261055
transform 1 0 37152 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_821
timestamp 1621261055
transform 1 0 38112 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_379
timestamp 1621261055
transform 1 0 37536 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_383
timestamp 1621261055
transform 1 0 37920 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_386
timestamp 1621261055
transform 1 0 38208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_394
timestamp 1621261055
transform 1 0 38976 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_402
timestamp 1621261055
transform 1 0 39744 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_383
timestamp 1621261055
transform 1 0 37920 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_391
timestamp 1621261055
transform 1 0 38688 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_399
timestamp 1621261055
transform 1 0 39456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_832
timestamp 1621261055
transform 1 0 40800 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_410
timestamp 1621261055
transform 1 0 40512 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_418
timestamp 1621261055
transform 1 0 41280 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_426
timestamp 1621261055
transform 1 0 42048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_407
timestamp 1621261055
transform 1 0 40224 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_411
timestamp 1621261055
transform 1 0 40608 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_414
timestamp 1621261055
transform 1 0 40896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_422
timestamp 1621261055
transform 1 0 41664 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_430
timestamp 1621261055
transform 1 0 42432 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_822
timestamp 1621261055
transform 1 0 43392 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_434
timestamp 1621261055
transform 1 0 42816 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_438
timestamp 1621261055
transform 1 0 43200 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_441
timestamp 1621261055
transform 1 0 43488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_449
timestamp 1621261055
transform 1 0 44256 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_457
timestamp 1621261055
transform 1 0 45024 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_438
timestamp 1621261055
transform 1 0 43200 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_446
timestamp 1621261055
transform 1 0 43968 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_454
timestamp 1621261055
transform 1 0 44736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_833
timestamp 1621261055
transform 1 0 46080 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_465
timestamp 1621261055
transform 1 0 45792 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_473
timestamp 1621261055
transform 1 0 46560 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_481
timestamp 1621261055
transform 1 0 47328 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_462
timestamp 1621261055
transform 1 0 45504 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_466
timestamp 1621261055
transform 1 0 45888 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_469
timestamp 1621261055
transform 1 0 46176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_477
timestamp 1621261055
transform 1 0 46944 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_485
timestamp 1621261055
transform 1 0 47712 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_823
timestamp 1621261055
transform 1 0 48672 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_489
timestamp 1621261055
transform 1 0 48096 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_493
timestamp 1621261055
transform 1 0 48480 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_496
timestamp 1621261055
transform 1 0 48768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_504
timestamp 1621261055
transform 1 0 49536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_512
timestamp 1621261055
transform 1 0 50304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_493
timestamp 1621261055
transform 1 0 48480 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_501
timestamp 1621261055
transform 1 0 49248 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_509
timestamp 1621261055
transform 1 0 50016 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_834
timestamp 1621261055
transform 1 0 51360 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_520
timestamp 1621261055
transform 1 0 51072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_528
timestamp 1621261055
transform 1 0 51840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_536
timestamp 1621261055
transform 1 0 52608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_517
timestamp 1621261055
transform 1 0 50784 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_521
timestamp 1621261055
transform 1 0 51168 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_524
timestamp 1621261055
transform 1 0 51456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_532
timestamp 1621261055
transform 1 0 52224 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_540
timestamp 1621261055
transform 1 0 52992 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_824
timestamp 1621261055
transform 1 0 53952 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_61_544
timestamp 1621261055
transform 1 0 53376 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_548
timestamp 1621261055
transform 1 0 53760 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_551
timestamp 1621261055
transform 1 0 54048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_559
timestamp 1621261055
transform 1 0 54816 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_567
timestamp 1621261055
transform 1 0 55584 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_548
timestamp 1621261055
transform 1 0 53760 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_556
timestamp 1621261055
transform 1 0 54528 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_564
timestamp 1621261055
transform 1 0 55296 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_835
timestamp 1621261055
transform 1 0 56640 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_575
timestamp 1621261055
transform 1 0 56352 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_583
timestamp 1621261055
transform 1 0 57120 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_591
timestamp 1621261055
transform 1 0 57888 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_62_572
timestamp 1621261055
transform 1 0 56064 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_576
timestamp 1621261055
transform 1 0 56448 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_579
timestamp 1621261055
transform 1 0 56736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_587
timestamp 1621261055
transform 1 0 57504 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_123
timestamp 1621261055
transform -1 0 58848 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_125
timestamp 1621261055
transform -1 0 58848 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_595
timestamp 1621261055
transform 1 0 58272 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_595
timestamp 1621261055
transform 1 0 58272 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_126
timestamp 1621261055
transform 1 0 1152 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_4
timestamp 1621261055
transform 1 0 1536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_12
timestamp 1621261055
transform 1 0 2304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_20
timestamp 1621261055
transform 1 0 3072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_28
timestamp 1621261055
transform 1 0 3840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_36
timestamp 1621261055
transform 1 0 4608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_44
timestamp 1621261055
transform 1 0 5376 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_52
timestamp 1621261055
transform 1 0 6144 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_54
timestamp 1621261055
transform 1 0 6336 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_836
timestamp 1621261055
transform 1 0 6432 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_56
timestamp 1621261055
transform 1 0 6528 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_64
timestamp 1621261055
transform 1 0 7296 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_72
timestamp 1621261055
transform 1 0 8064 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_80
timestamp 1621261055
transform 1 0 8832 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_88
timestamp 1621261055
transform 1 0 9600 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_96
timestamp 1621261055
transform 1 0 10368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_104
timestamp 1621261055
transform 1 0 11136 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_108
timestamp 1621261055
transform 1 0 11520 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_837
timestamp 1621261055
transform 1 0 11712 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_111
timestamp 1621261055
transform 1 0 11808 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_119
timestamp 1621261055
transform 1 0 12576 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_127
timestamp 1621261055
transform 1 0 13344 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_135
timestamp 1621261055
transform 1 0 14112 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_143
timestamp 1621261055
transform 1 0 14880 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_151
timestamp 1621261055
transform 1 0 15648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_159
timestamp 1621261055
transform 1 0 16416 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_838
timestamp 1621261055
transform 1 0 16992 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_163
timestamp 1621261055
transform 1 0 16800 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_166
timestamp 1621261055
transform 1 0 17088 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_174
timestamp 1621261055
transform 1 0 17856 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_182
timestamp 1621261055
transform 1 0 18624 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_190
timestamp 1621261055
transform 1 0 19392 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_198
timestamp 1621261055
transform 1 0 20160 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_206
timestamp 1621261055
transform 1 0 20928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_214
timestamp 1621261055
transform 1 0 21696 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_839
timestamp 1621261055
transform 1 0 22272 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_218
timestamp 1621261055
transform 1 0 22080 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_221
timestamp 1621261055
transform 1 0 22368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_229
timestamp 1621261055
transform 1 0 23136 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_237
timestamp 1621261055
transform 1 0 23904 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_245
timestamp 1621261055
transform 1 0 24672 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_253
timestamp 1621261055
transform 1 0 25440 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_261
timestamp 1621261055
transform 1 0 26208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_269
timestamp 1621261055
transform 1 0 26976 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_840
timestamp 1621261055
transform 1 0 27552 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_273
timestamp 1621261055
transform 1 0 27360 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_276
timestamp 1621261055
transform 1 0 27648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_284
timestamp 1621261055
transform 1 0 28416 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_292
timestamp 1621261055
transform 1 0 29184 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_300
timestamp 1621261055
transform 1 0 29952 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_308
timestamp 1621261055
transform 1 0 30720 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_316
timestamp 1621261055
transform 1 0 31488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_324
timestamp 1621261055
transform 1 0 32256 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_841
timestamp 1621261055
transform 1 0 32832 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_328
timestamp 1621261055
transform 1 0 32640 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_331
timestamp 1621261055
transform 1 0 32928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_339
timestamp 1621261055
transform 1 0 33696 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_347
timestamp 1621261055
transform 1 0 34464 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_355
timestamp 1621261055
transform 1 0 35232 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_363
timestamp 1621261055
transform 1 0 36000 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_371
timestamp 1621261055
transform 1 0 36768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_842
timestamp 1621261055
transform 1 0 38112 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_379
timestamp 1621261055
transform 1 0 37536 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_383
timestamp 1621261055
transform 1 0 37920 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_386
timestamp 1621261055
transform 1 0 38208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_394
timestamp 1621261055
transform 1 0 38976 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_402
timestamp 1621261055
transform 1 0 39744 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_410
timestamp 1621261055
transform 1 0 40512 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_418
timestamp 1621261055
transform 1 0 41280 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_426
timestamp 1621261055
transform 1 0 42048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _119_
timestamp 1621261055
transform -1 0 44352 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_843
timestamp 1621261055
transform 1 0 43392 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_180
timestamp 1621261055
transform -1 0 44064 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_63_434
timestamp 1621261055
transform 1 0 42816 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_438
timestamp 1621261055
transform 1 0 43200 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_63_441
timestamp 1621261055
transform 1 0 43488 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_450
timestamp 1621261055
transform 1 0 44352 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_458
timestamp 1621261055
transform 1 0 45120 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _140_
timestamp 1621261055
transform -1 0 47904 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_201
timestamp 1621261055
transform -1 0 47616 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_466
timestamp 1621261055
transform 1 0 45888 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_474
timestamp 1621261055
transform 1 0 46656 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_844
timestamp 1621261055
transform 1 0 48672 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_487
timestamp 1621261055
transform 1 0 47904 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_496
timestamp 1621261055
transform 1 0 48768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_504
timestamp 1621261055
transform 1 0 49536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_512
timestamp 1621261055
transform 1 0 50304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_520
timestamp 1621261055
transform 1 0 51072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_528
timestamp 1621261055
transform 1 0 51840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_536
timestamp 1621261055
transform 1 0 52608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_845
timestamp 1621261055
transform 1 0 53952 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_544
timestamp 1621261055
transform 1 0 53376 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_548
timestamp 1621261055
transform 1 0 53760 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_551
timestamp 1621261055
transform 1 0 54048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_559
timestamp 1621261055
transform 1 0 54816 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_567
timestamp 1621261055
transform 1 0 55584 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_575
timestamp 1621261055
transform 1 0 56352 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_583
timestamp 1621261055
transform 1 0 57120 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_591
timestamp 1621261055
transform 1 0 57888 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_127
timestamp 1621261055
transform -1 0 58848 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_595
timestamp 1621261055
transform 1 0 58272 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_128
timestamp 1621261055
transform 1 0 1152 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_64_4
timestamp 1621261055
transform 1 0 1536 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_12
timestamp 1621261055
transform 1 0 2304 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_20
timestamp 1621261055
transform 1 0 3072 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _163_
timestamp 1621261055
transform 1 0 6336 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_846
timestamp 1621261055
transform 1 0 3840 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_109
timestamp 1621261055
transform 1 0 6144 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_29
timestamp 1621261055
transform 1 0 3936 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_37
timestamp 1621261055
transform 1 0 4704 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_45
timestamp 1621261055
transform 1 0 5472 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_49
timestamp 1621261055
transform 1 0 5856 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_51
timestamp 1621261055
transform 1 0 6048 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_57
timestamp 1621261055
transform 1 0 6624 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_65
timestamp 1621261055
transform 1 0 7392 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_73
timestamp 1621261055
transform 1 0 8160 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_81
timestamp 1621261055
transform 1 0 8928 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_847
timestamp 1621261055
transform 1 0 9120 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_84
timestamp 1621261055
transform 1 0 9216 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_92
timestamp 1621261055
transform 1 0 9984 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_100
timestamp 1621261055
transform 1 0 10752 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_108
timestamp 1621261055
transform 1 0 11520 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_116
timestamp 1621261055
transform 1 0 12288 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_124
timestamp 1621261055
transform 1 0 13056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_132
timestamp 1621261055
transform 1 0 13824 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_848
timestamp 1621261055
transform 1 0 14400 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_136
timestamp 1621261055
transform 1 0 14208 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_139
timestamp 1621261055
transform 1 0 14496 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_147
timestamp 1621261055
transform 1 0 15264 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_155
timestamp 1621261055
transform 1 0 16032 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_163
timestamp 1621261055
transform 1 0 16800 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_171
timestamp 1621261055
transform 1 0 17568 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_179
timestamp 1621261055
transform 1 0 18336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_187
timestamp 1621261055
transform 1 0 19104 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_849
timestamp 1621261055
transform 1 0 19680 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_191
timestamp 1621261055
transform 1 0 19488 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_194
timestamp 1621261055
transform 1 0 19776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_202
timestamp 1621261055
transform 1 0 20544 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_210
timestamp 1621261055
transform 1 0 21312 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_218
timestamp 1621261055
transform 1 0 22080 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_226
timestamp 1621261055
transform 1 0 22848 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_234
timestamp 1621261055
transform 1 0 23616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_242
timestamp 1621261055
transform 1 0 24384 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_850
timestamp 1621261055
transform 1 0 24960 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_246
timestamp 1621261055
transform 1 0 24768 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_249
timestamp 1621261055
transform 1 0 25056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_257
timestamp 1621261055
transform 1 0 25824 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_265
timestamp 1621261055
transform 1 0 26592 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_273
timestamp 1621261055
transform 1 0 27360 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_281
timestamp 1621261055
transform 1 0 28128 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_289
timestamp 1621261055
transform 1 0 28896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_297
timestamp 1621261055
transform 1 0 29664 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_851
timestamp 1621261055
transform 1 0 30240 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_301
timestamp 1621261055
transform 1 0 30048 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_304
timestamp 1621261055
transform 1 0 30336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_312
timestamp 1621261055
transform 1 0 31104 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_320
timestamp 1621261055
transform 1 0 31872 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_328
timestamp 1621261055
transform 1 0 32640 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_336
timestamp 1621261055
transform 1 0 33408 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_344
timestamp 1621261055
transform 1 0 34176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_852
timestamp 1621261055
transform 1 0 35520 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_352
timestamp 1621261055
transform 1 0 34944 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_356
timestamp 1621261055
transform 1 0 35328 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_359
timestamp 1621261055
transform 1 0 35616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_367
timestamp 1621261055
transform 1 0 36384 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_375
timestamp 1621261055
transform 1 0 37152 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_383
timestamp 1621261055
transform 1 0 37920 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_391
timestamp 1621261055
transform 1 0 38688 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_399
timestamp 1621261055
transform 1 0 39456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _128_
timestamp 1621261055
transform -1 0 41568 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_853
timestamp 1621261055
transform 1 0 40800 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_186
timestamp 1621261055
transform -1 0 41280 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_64_407
timestamp 1621261055
transform 1 0 40224 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_411
timestamp 1621261055
transform 1 0 40608 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_414
timestamp 1621261055
transform 1 0 40896 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_421
timestamp 1621261055
transform 1 0 41568 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_429
timestamp 1621261055
transform 1 0 42336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_437
timestamp 1621261055
transform 1 0 43104 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_445
timestamp 1621261055
transform 1 0 43872 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_453
timestamp 1621261055
transform 1 0 44640 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_854
timestamp 1621261055
transform 1 0 46080 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_461
timestamp 1621261055
transform 1 0 45408 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_465
timestamp 1621261055
transform 1 0 45792 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_467
timestamp 1621261055
transform 1 0 45984 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_469
timestamp 1621261055
transform 1 0 46176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_477
timestamp 1621261055
transform 1 0 46944 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_485
timestamp 1621261055
transform 1 0 47712 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_493
timestamp 1621261055
transform 1 0 48480 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_501
timestamp 1621261055
transform 1 0 49248 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_509
timestamp 1621261055
transform 1 0 50016 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_855
timestamp 1621261055
transform 1 0 51360 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_517
timestamp 1621261055
transform 1 0 50784 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_521
timestamp 1621261055
transform 1 0 51168 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_524
timestamp 1621261055
transform 1 0 51456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_532
timestamp 1621261055
transform 1 0 52224 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_540
timestamp 1621261055
transform 1 0 52992 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_548
timestamp 1621261055
transform 1 0 53760 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_556
timestamp 1621261055
transform 1 0 54528 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_564
timestamp 1621261055
transform 1 0 55296 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_856
timestamp 1621261055
transform 1 0 56640 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_572
timestamp 1621261055
transform 1 0 56064 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_576
timestamp 1621261055
transform 1 0 56448 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_579
timestamp 1621261055
transform 1 0 56736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_587
timestamp 1621261055
transform 1 0 57504 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_129
timestamp 1621261055
transform -1 0 58848 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_595
timestamp 1621261055
transform 1 0 58272 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_130
timestamp 1621261055
transform 1 0 1152 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_4
timestamp 1621261055
transform 1 0 1536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_12
timestamp 1621261055
transform 1 0 2304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_20
timestamp 1621261055
transform 1 0 3072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_28
timestamp 1621261055
transform 1 0 3840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_36
timestamp 1621261055
transform 1 0 4608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_44
timestamp 1621261055
transform 1 0 5376 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_52
timestamp 1621261055
transform 1 0 6144 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_54
timestamp 1621261055
transform 1 0 6336 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_857
timestamp 1621261055
transform 1 0 6432 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_56
timestamp 1621261055
transform 1 0 6528 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_64
timestamp 1621261055
transform 1 0 7296 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_72
timestamp 1621261055
transform 1 0 8064 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_80
timestamp 1621261055
transform 1 0 8832 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _058_
timestamp 1621261055
transform 1 0 10656 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_65_88
timestamp 1621261055
transform 1 0 9600 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_96
timestamp 1621261055
transform 1 0 10368 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_98
timestamp 1621261055
transform 1 0 10560 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_102
timestamp 1621261055
transform 1 0 10944 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_858
timestamp 1621261055
transform 1 0 11712 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_111
timestamp 1621261055
transform 1 0 11808 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_119
timestamp 1621261055
transform 1 0 12576 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_127
timestamp 1621261055
transform 1 0 13344 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_135
timestamp 1621261055
transform 1 0 14112 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_143
timestamp 1621261055
transform 1 0 14880 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_151
timestamp 1621261055
transform 1 0 15648 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_159
timestamp 1621261055
transform 1 0 16416 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_859
timestamp 1621261055
transform 1 0 16992 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_163
timestamp 1621261055
transform 1 0 16800 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_166
timestamp 1621261055
transform 1 0 17088 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_174
timestamp 1621261055
transform 1 0 17856 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_182
timestamp 1621261055
transform 1 0 18624 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_190
timestamp 1621261055
transform 1 0 19392 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_198
timestamp 1621261055
transform 1 0 20160 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_206
timestamp 1621261055
transform 1 0 20928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_214
timestamp 1621261055
transform 1 0 21696 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_860
timestamp 1621261055
transform 1 0 22272 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_218
timestamp 1621261055
transform 1 0 22080 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_221
timestamp 1621261055
transform 1 0 22368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_229
timestamp 1621261055
transform 1 0 23136 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_237
timestamp 1621261055
transform 1 0 23904 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_241
timestamp 1621261055
transform 1 0 24288 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_243
timestamp 1621261055
transform 1 0 24480 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _030_
timestamp 1621261055
transform 1 0 24576 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_65_247
timestamp 1621261055
transform 1 0 24864 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_255
timestamp 1621261055
transform 1 0 25632 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_263
timestamp 1621261055
transform 1 0 26400 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _127_
timestamp 1621261055
transform 1 0 28032 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_861
timestamp 1621261055
transform 1 0 27552 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_184
timestamp 1621261055
transform 1 0 27840 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_65_271
timestamp 1621261055
transform 1 0 27168 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_276
timestamp 1621261055
transform 1 0 27648 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_283
timestamp 1621261055
transform 1 0 28320 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_291
timestamp 1621261055
transform 1 0 29088 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _018_
timestamp 1621261055
transform 1 0 31392 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_65_299
timestamp 1621261055
transform 1 0 29856 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_307
timestamp 1621261055
transform 1 0 30624 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_318
timestamp 1621261055
transform 1 0 31680 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_862
timestamp 1621261055
transform 1 0 32832 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_326
timestamp 1621261055
transform 1 0 32448 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_331
timestamp 1621261055
transform 1 0 32928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_339
timestamp 1621261055
transform 1 0 33696 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_347
timestamp 1621261055
transform 1 0 34464 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_355
timestamp 1621261055
transform 1 0 35232 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_363
timestamp 1621261055
transform 1 0 36000 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_371
timestamp 1621261055
transform 1 0 36768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_863
timestamp 1621261055
transform 1 0 38112 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_379
timestamp 1621261055
transform 1 0 37536 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_383
timestamp 1621261055
transform 1 0 37920 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_386
timestamp 1621261055
transform 1 0 38208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_394
timestamp 1621261055
transform 1 0 38976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_402
timestamp 1621261055
transform 1 0 39744 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_410
timestamp 1621261055
transform 1 0 40512 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_418
timestamp 1621261055
transform 1 0 41280 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_426
timestamp 1621261055
transform 1 0 42048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _081_
timestamp 1621261055
transform -1 0 44160 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_864
timestamp 1621261055
transform 1 0 43392 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_145
timestamp 1621261055
transform -1 0 43872 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_65_434
timestamp 1621261055
transform 1 0 42816 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_438
timestamp 1621261055
transform 1 0 43200 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_441
timestamp 1621261055
transform 1 0 43488 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_448
timestamp 1621261055
transform 1 0 44160 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_456
timestamp 1621261055
transform 1 0 44928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_464
timestamp 1621261055
transform 1 0 45696 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_472
timestamp 1621261055
transform 1 0 46464 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_480
timestamp 1621261055
transform 1 0 47232 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_865
timestamp 1621261055
transform 1 0 48672 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_488
timestamp 1621261055
transform 1 0 48000 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_492
timestamp 1621261055
transform 1 0 48384 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_494
timestamp 1621261055
transform 1 0 48576 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_496
timestamp 1621261055
transform 1 0 48768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_504
timestamp 1621261055
transform 1 0 49536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_512
timestamp 1621261055
transform 1 0 50304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_520
timestamp 1621261055
transform 1 0 51072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_528
timestamp 1621261055
transform 1 0 51840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_536
timestamp 1621261055
transform 1 0 52608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_866
timestamp 1621261055
transform 1 0 53952 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_544
timestamp 1621261055
transform 1 0 53376 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_548
timestamp 1621261055
transform 1 0 53760 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_551
timestamp 1621261055
transform 1 0 54048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_559
timestamp 1621261055
transform 1 0 54816 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_567
timestamp 1621261055
transform 1 0 55584 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_575
timestamp 1621261055
transform 1 0 56352 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_583
timestamp 1621261055
transform 1 0 57120 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_591
timestamp 1621261055
transform 1 0 57888 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_131
timestamp 1621261055
transform -1 0 58848 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_595
timestamp 1621261055
transform 1 0 58272 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _069_
timestamp 1621261055
transform 1 0 2784 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_132
timestamp 1621261055
transform 1 0 1152 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_133
timestamp 1621261055
transform 1 0 2592 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_4
timestamp 1621261055
transform 1 0 1536 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_12
timestamp 1621261055
transform 1 0 2304 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_66_14
timestamp 1621261055
transform 1 0 2496 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_20
timestamp 1621261055
transform 1 0 3072 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_867
timestamp 1621261055
transform 1 0 3840 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_29
timestamp 1621261055
transform 1 0 3936 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_37
timestamp 1621261055
transform 1 0 4704 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_45
timestamp 1621261055
transform 1 0 5472 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_53
timestamp 1621261055
transform 1 0 6240 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _016_
timestamp 1621261055
transform 1 0 6624 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_66_60
timestamp 1621261055
transform 1 0 6912 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_68
timestamp 1621261055
transform 1 0 7680 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_76
timestamp 1621261055
transform 1 0 8448 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_80
timestamp 1621261055
transform 1 0 8832 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_868
timestamp 1621261055
transform 1 0 9120 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_66_82
timestamp 1621261055
transform 1 0 9024 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_84
timestamp 1621261055
transform 1 0 9216 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_92
timestamp 1621261055
transform 1 0 9984 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_100
timestamp 1621261055
transform 1 0 10752 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_108
timestamp 1621261055
transform 1 0 11520 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _195_
timestamp 1621261055
transform -1 0 13536 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_226
timestamp 1621261055
transform -1 0 13248 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_116
timestamp 1621261055
transform 1 0 12288 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_129
timestamp 1621261055
transform 1 0 13536 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_869
timestamp 1621261055
transform 1 0 14400 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_66_137
timestamp 1621261055
transform 1 0 14304 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_139
timestamp 1621261055
transform 1 0 14496 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_147
timestamp 1621261055
transform 1 0 15264 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_155
timestamp 1621261055
transform 1 0 16032 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_163
timestamp 1621261055
transform 1 0 16800 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_171
timestamp 1621261055
transform 1 0 17568 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_179
timestamp 1621261055
transform 1 0 18336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_187
timestamp 1621261055
transform 1 0 19104 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_870
timestamp 1621261055
transform 1 0 19680 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_191
timestamp 1621261055
transform 1 0 19488 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_194
timestamp 1621261055
transform 1 0 19776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_202
timestamp 1621261055
transform 1 0 20544 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_210
timestamp 1621261055
transform 1 0 21312 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_218
timestamp 1621261055
transform 1 0 22080 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_226
timestamp 1621261055
transform 1 0 22848 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_234
timestamp 1621261055
transform 1 0 23616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_242
timestamp 1621261055
transform 1 0 24384 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_871
timestamp 1621261055
transform 1 0 24960 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_246
timestamp 1621261055
transform 1 0 24768 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_249
timestamp 1621261055
transform 1 0 25056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_257
timestamp 1621261055
transform 1 0 25824 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_265
timestamp 1621261055
transform 1 0 26592 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_273
timestamp 1621261055
transform 1 0 27360 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_281
timestamp 1621261055
transform 1 0 28128 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_289
timestamp 1621261055
transform 1 0 28896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_297
timestamp 1621261055
transform 1 0 29664 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_872
timestamp 1621261055
transform 1 0 30240 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_301
timestamp 1621261055
transform 1 0 30048 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_304
timestamp 1621261055
transform 1 0 30336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_312
timestamp 1621261055
transform 1 0 31104 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_320
timestamp 1621261055
transform 1 0 31872 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_328
timestamp 1621261055
transform 1 0 32640 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_336
timestamp 1621261055
transform 1 0 33408 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_344
timestamp 1621261055
transform 1 0 34176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_873
timestamp 1621261055
transform 1 0 35520 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_352
timestamp 1621261055
transform 1 0 34944 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_356
timestamp 1621261055
transform 1 0 35328 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_359
timestamp 1621261055
transform 1 0 35616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_367
timestamp 1621261055
transform 1 0 36384 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_375
timestamp 1621261055
transform 1 0 37152 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_383
timestamp 1621261055
transform 1 0 37920 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_391
timestamp 1621261055
transform 1 0 38688 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_399
timestamp 1621261055
transform 1 0 39456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_874
timestamp 1621261055
transform 1 0 40800 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_407
timestamp 1621261055
transform 1 0 40224 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_411
timestamp 1621261055
transform 1 0 40608 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_414
timestamp 1621261055
transform 1 0 40896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_422
timestamp 1621261055
transform 1 0 41664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_430
timestamp 1621261055
transform 1 0 42432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_438
timestamp 1621261055
transform 1 0 43200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_446
timestamp 1621261055
transform 1 0 43968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_454
timestamp 1621261055
transform 1 0 44736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_875
timestamp 1621261055
transform 1 0 46080 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_462
timestamp 1621261055
transform 1 0 45504 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_466
timestamp 1621261055
transform 1 0 45888 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_469
timestamp 1621261055
transform 1 0 46176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_477
timestamp 1621261055
transform 1 0 46944 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_485
timestamp 1621261055
transform 1 0 47712 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_493
timestamp 1621261055
transform 1 0 48480 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_501
timestamp 1621261055
transform 1 0 49248 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_509
timestamp 1621261055
transform 1 0 50016 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_876
timestamp 1621261055
transform 1 0 51360 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_517
timestamp 1621261055
transform 1 0 50784 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_521
timestamp 1621261055
transform 1 0 51168 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_524
timestamp 1621261055
transform 1 0 51456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_532
timestamp 1621261055
transform 1 0 52224 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_540
timestamp 1621261055
transform 1 0 52992 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_548
timestamp 1621261055
transform 1 0 53760 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_556
timestamp 1621261055
transform 1 0 54528 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_564
timestamp 1621261055
transform 1 0 55296 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_877
timestamp 1621261055
transform 1 0 56640 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_66_572
timestamp 1621261055
transform 1 0 56064 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_576
timestamp 1621261055
transform 1 0 56448 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_579
timestamp 1621261055
transform 1 0 56736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_587
timestamp 1621261055
transform 1 0 57504 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_133
timestamp 1621261055
transform -1 0 58848 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_595
timestamp 1621261055
transform 1 0 58272 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_134
timestamp 1621261055
transform 1 0 1152 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_4
timestamp 1621261055
transform 1 0 1536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_12
timestamp 1621261055
transform 1 0 2304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_20
timestamp 1621261055
transform 1 0 3072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_28
timestamp 1621261055
transform 1 0 3840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_36
timestamp 1621261055
transform 1 0 4608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_44
timestamp 1621261055
transform 1 0 5376 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_52
timestamp 1621261055
transform 1 0 6144 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_54
timestamp 1621261055
transform 1 0 6336 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_878
timestamp 1621261055
transform 1 0 6432 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_56
timestamp 1621261055
transform 1 0 6528 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_64
timestamp 1621261055
transform 1 0 7296 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_72
timestamp 1621261055
transform 1 0 8064 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_80
timestamp 1621261055
transform 1 0 8832 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_88
timestamp 1621261055
transform 1 0 9600 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_96
timestamp 1621261055
transform 1 0 10368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_104
timestamp 1621261055
transform 1 0 11136 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_108
timestamp 1621261055
transform 1 0 11520 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_879
timestamp 1621261055
transform 1 0 11712 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_111
timestamp 1621261055
transform 1 0 11808 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_119
timestamp 1621261055
transform 1 0 12576 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_127
timestamp 1621261055
transform 1 0 13344 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_135
timestamp 1621261055
transform 1 0 14112 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_143
timestamp 1621261055
transform 1 0 14880 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_151
timestamp 1621261055
transform 1 0 15648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_159
timestamp 1621261055
transform 1 0 16416 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_880
timestamp 1621261055
transform 1 0 16992 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_163
timestamp 1621261055
transform 1 0 16800 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_166
timestamp 1621261055
transform 1 0 17088 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_174
timestamp 1621261055
transform 1 0 17856 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_182
timestamp 1621261055
transform 1 0 18624 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_190
timestamp 1621261055
transform 1 0 19392 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_198
timestamp 1621261055
transform 1 0 20160 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_206
timestamp 1621261055
transform 1 0 20928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_214
timestamp 1621261055
transform 1 0 21696 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_881
timestamp 1621261055
transform 1 0 22272 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_218
timestamp 1621261055
transform 1 0 22080 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_221
timestamp 1621261055
transform 1 0 22368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_229
timestamp 1621261055
transform 1 0 23136 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_237
timestamp 1621261055
transform 1 0 23904 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_245
timestamp 1621261055
transform 1 0 24672 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_253
timestamp 1621261055
transform 1 0 25440 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_261
timestamp 1621261055
transform 1 0 26208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_269
timestamp 1621261055
transform 1 0 26976 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _107_
timestamp 1621261055
transform 1 0 28032 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_882
timestamp 1621261055
transform 1 0 27552 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_169
timestamp 1621261055
transform 1 0 27840 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_273
timestamp 1621261055
transform 1 0 27360 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_276
timestamp 1621261055
transform 1 0 27648 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_283
timestamp 1621261055
transform 1 0 28320 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_291
timestamp 1621261055
transform 1 0 29088 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _043_
timestamp 1621261055
transform 1 0 31200 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_67_299
timestamp 1621261055
transform 1 0 29856 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_307
timestamp 1621261055
transform 1 0 30624 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_311
timestamp 1621261055
transform 1 0 31008 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_316
timestamp 1621261055
transform 1 0 31488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_324
timestamp 1621261055
transform 1 0 32256 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_883
timestamp 1621261055
transform 1 0 32832 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_328
timestamp 1621261055
transform 1 0 32640 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_331
timestamp 1621261055
transform 1 0 32928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_339
timestamp 1621261055
transform 1 0 33696 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_347
timestamp 1621261055
transform 1 0 34464 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_355
timestamp 1621261055
transform 1 0 35232 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_363
timestamp 1621261055
transform 1 0 36000 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_371
timestamp 1621261055
transform 1 0 36768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_884
timestamp 1621261055
transform 1 0 38112 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_379
timestamp 1621261055
transform 1 0 37536 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_383
timestamp 1621261055
transform 1 0 37920 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_386
timestamp 1621261055
transform 1 0 38208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_394
timestamp 1621261055
transform 1 0 38976 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_402
timestamp 1621261055
transform 1 0 39744 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_410
timestamp 1621261055
transform 1 0 40512 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_418
timestamp 1621261055
transform 1 0 41280 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_426
timestamp 1621261055
transform 1 0 42048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_885
timestamp 1621261055
transform 1 0 43392 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_434
timestamp 1621261055
transform 1 0 42816 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_438
timestamp 1621261055
transform 1 0 43200 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_441
timestamp 1621261055
transform 1 0 43488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_449
timestamp 1621261055
transform 1 0 44256 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_457
timestamp 1621261055
transform 1 0 45024 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_465
timestamp 1621261055
transform 1 0 45792 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_473
timestamp 1621261055
transform 1 0 46560 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_481
timestamp 1621261055
transform 1 0 47328 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_886
timestamp 1621261055
transform 1 0 48672 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_489
timestamp 1621261055
transform 1 0 48096 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_493
timestamp 1621261055
transform 1 0 48480 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_496
timestamp 1621261055
transform 1 0 48768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_504
timestamp 1621261055
transform 1 0 49536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_512
timestamp 1621261055
transform 1 0 50304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_520
timestamp 1621261055
transform 1 0 51072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_528
timestamp 1621261055
transform 1 0 51840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_536
timestamp 1621261055
transform 1 0 52608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _213_
timestamp 1621261055
transform -1 0 54720 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_887
timestamp 1621261055
transform 1 0 53952 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_245
timestamp 1621261055
transform -1 0 54432 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_67_544
timestamp 1621261055
transform 1 0 53376 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_548
timestamp 1621261055
transform 1 0 53760 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_551
timestamp 1621261055
transform 1 0 54048 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_558
timestamp 1621261055
transform 1 0 54720 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_566
timestamp 1621261055
transform 1 0 55488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_574
timestamp 1621261055
transform 1 0 56256 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_582
timestamp 1621261055
transform 1 0 57024 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_590
timestamp 1621261055
transform 1 0 57792 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_594
timestamp 1621261055
transform 1 0 58176 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_135
timestamp 1621261055
transform -1 0 58848 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_67_596
timestamp 1621261055
transform 1 0 58368 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_136
timestamp 1621261055
transform 1 0 1152 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_4
timestamp 1621261055
transform 1 0 1536 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_12
timestamp 1621261055
transform 1 0 2304 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_20
timestamp 1621261055
transform 1 0 3072 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_888
timestamp 1621261055
transform 1 0 3840 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_29
timestamp 1621261055
transform 1 0 3936 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_37
timestamp 1621261055
transform 1 0 4704 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_45
timestamp 1621261055
transform 1 0 5472 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_53
timestamp 1621261055
transform 1 0 6240 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_61
timestamp 1621261055
transform 1 0 7008 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_69
timestamp 1621261055
transform 1 0 7776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_77
timestamp 1621261055
transform 1 0 8544 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_81
timestamp 1621261055
transform 1 0 8928 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_889
timestamp 1621261055
transform 1 0 9120 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_84
timestamp 1621261055
transform 1 0 9216 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_92
timestamp 1621261055
transform 1 0 9984 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_100
timestamp 1621261055
transform 1 0 10752 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_108
timestamp 1621261055
transform 1 0 11520 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_116
timestamp 1621261055
transform 1 0 12288 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_124
timestamp 1621261055
transform 1 0 13056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_132
timestamp 1621261055
transform 1 0 13824 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_890
timestamp 1621261055
transform 1 0 14400 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_136
timestamp 1621261055
transform 1 0 14208 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_139
timestamp 1621261055
transform 1 0 14496 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_147
timestamp 1621261055
transform 1 0 15264 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_155
timestamp 1621261055
transform 1 0 16032 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_163
timestamp 1621261055
transform 1 0 16800 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_171
timestamp 1621261055
transform 1 0 17568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_179
timestamp 1621261055
transform 1 0 18336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_187
timestamp 1621261055
transform 1 0 19104 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_891
timestamp 1621261055
transform 1 0 19680 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_191
timestamp 1621261055
transform 1 0 19488 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_194
timestamp 1621261055
transform 1 0 19776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_202
timestamp 1621261055
transform 1 0 20544 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_210
timestamp 1621261055
transform 1 0 21312 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_218
timestamp 1621261055
transform 1 0 22080 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_226
timestamp 1621261055
transform 1 0 22848 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_234
timestamp 1621261055
transform 1 0 23616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_242
timestamp 1621261055
transform 1 0 24384 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_892
timestamp 1621261055
transform 1 0 24960 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_246
timestamp 1621261055
transform 1 0 24768 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_249
timestamp 1621261055
transform 1 0 25056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_257
timestamp 1621261055
transform 1 0 25824 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_265
timestamp 1621261055
transform 1 0 26592 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_273
timestamp 1621261055
transform 1 0 27360 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_281
timestamp 1621261055
transform 1 0 28128 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_289
timestamp 1621261055
transform 1 0 28896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_297
timestamp 1621261055
transform 1 0 29664 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_893
timestamp 1621261055
transform 1 0 30240 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_301
timestamp 1621261055
transform 1 0 30048 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_304
timestamp 1621261055
transform 1 0 30336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_312
timestamp 1621261055
transform 1 0 31104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_320
timestamp 1621261055
transform 1 0 31872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_328
timestamp 1621261055
transform 1 0 32640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_336
timestamp 1621261055
transform 1 0 33408 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_344
timestamp 1621261055
transform 1 0 34176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_894
timestamp 1621261055
transform 1 0 35520 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_352
timestamp 1621261055
transform 1 0 34944 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_356
timestamp 1621261055
transform 1 0 35328 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_359
timestamp 1621261055
transform 1 0 35616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_367
timestamp 1621261055
transform 1 0 36384 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_375
timestamp 1621261055
transform 1 0 37152 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_383
timestamp 1621261055
transform 1 0 37920 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_391
timestamp 1621261055
transform 1 0 38688 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_399
timestamp 1621261055
transform 1 0 39456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_895
timestamp 1621261055
transform 1 0 40800 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_407
timestamp 1621261055
transform 1 0 40224 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_411
timestamp 1621261055
transform 1 0 40608 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_414
timestamp 1621261055
transform 1 0 40896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_422
timestamp 1621261055
transform 1 0 41664 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_430
timestamp 1621261055
transform 1 0 42432 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_438
timestamp 1621261055
transform 1 0 43200 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_446
timestamp 1621261055
transform 1 0 43968 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_454
timestamp 1621261055
transform 1 0 44736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_896
timestamp 1621261055
transform 1 0 46080 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_462
timestamp 1621261055
transform 1 0 45504 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_466
timestamp 1621261055
transform 1 0 45888 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_469
timestamp 1621261055
transform 1 0 46176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_477
timestamp 1621261055
transform 1 0 46944 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_485
timestamp 1621261055
transform 1 0 47712 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_493
timestamp 1621261055
transform 1 0 48480 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_501
timestamp 1621261055
transform 1 0 49248 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_509
timestamp 1621261055
transform 1 0 50016 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_897
timestamp 1621261055
transform 1 0 51360 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_517
timestamp 1621261055
transform 1 0 50784 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_521
timestamp 1621261055
transform 1 0 51168 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_524
timestamp 1621261055
transform 1 0 51456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_532
timestamp 1621261055
transform 1 0 52224 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_540
timestamp 1621261055
transform 1 0 52992 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _200_
timestamp 1621261055
transform -1 0 55392 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_231
timestamp 1621261055
transform -1 0 55104 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_548
timestamp 1621261055
transform 1 0 53760 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_556
timestamp 1621261055
transform 1 0 54528 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_68_565
timestamp 1621261055
transform 1 0 55392 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_898
timestamp 1621261055
transform 1 0 56640 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_68_573
timestamp 1621261055
transform 1 0 56160 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_68_577
timestamp 1621261055
transform 1 0 56544 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_579
timestamp 1621261055
transform 1 0 56736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_587
timestamp 1621261055
transform 1 0 57504 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_137
timestamp 1621261055
transform -1 0 58848 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_595
timestamp 1621261055
transform 1 0 58272 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_138
timestamp 1621261055
transform 1 0 1152 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_140
timestamp 1621261055
transform 1 0 1152 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_4
timestamp 1621261055
transform 1 0 1536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_12
timestamp 1621261055
transform 1 0 2304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_20
timestamp 1621261055
transform 1 0 3072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_4
timestamp 1621261055
transform 1 0 1536 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_12
timestamp 1621261055
transform 1 0 2304 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_20
timestamp 1621261055
transform 1 0 3072 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_29
timestamp 1621261055
transform 1 0 3936 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_28
timestamp 1621261055
transform 1 0 3840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_909
timestamp 1621261055
transform 1 0 3840 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_37
timestamp 1621261055
transform 1 0 4704 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_44
timestamp 1621261055
transform 1 0 5376 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_36
timestamp 1621261055
transform 1 0 4608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_53
timestamp 1621261055
transform 1 0 6240 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_45
timestamp 1621261055
transform 1 0 5472 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_52
timestamp 1621261055
transform 1 0 6144 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_69_54
timestamp 1621261055
transform 1 0 6336 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_899
timestamp 1621261055
transform 1 0 6432 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_56
timestamp 1621261055
transform 1 0 6528 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_64
timestamp 1621261055
transform 1 0 7296 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_72
timestamp 1621261055
transform 1 0 8064 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_80
timestamp 1621261055
transform 1 0 8832 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_61
timestamp 1621261055
transform 1 0 7008 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_69
timestamp 1621261055
transform 1 0 7776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_77
timestamp 1621261055
transform 1 0 8544 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_81
timestamp 1621261055
transform 1 0 8928 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_910
timestamp 1621261055
transform 1 0 9120 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_88
timestamp 1621261055
transform 1 0 9600 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_96
timestamp 1621261055
transform 1 0 10368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_104
timestamp 1621261055
transform 1 0 11136 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_108
timestamp 1621261055
transform 1 0 11520 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_84
timestamp 1621261055
transform 1 0 9216 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_92
timestamp 1621261055
transform 1 0 9984 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_100
timestamp 1621261055
transform 1 0 10752 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_108
timestamp 1621261055
transform 1 0 11520 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_900
timestamp 1621261055
transform 1 0 11712 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_111
timestamp 1621261055
transform 1 0 11808 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_119
timestamp 1621261055
transform 1 0 12576 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_127
timestamp 1621261055
transform 1 0 13344 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_135
timestamp 1621261055
transform 1 0 14112 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_116
timestamp 1621261055
transform 1 0 12288 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_124
timestamp 1621261055
transform 1 0 13056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_132
timestamp 1621261055
transform 1 0 13824 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_911
timestamp 1621261055
transform 1 0 14400 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_143
timestamp 1621261055
transform 1 0 14880 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_151
timestamp 1621261055
transform 1 0 15648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_159
timestamp 1621261055
transform 1 0 16416 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_136
timestamp 1621261055
transform 1 0 14208 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_139
timestamp 1621261055
transform 1 0 14496 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_147
timestamp 1621261055
transform 1 0 15264 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_155
timestamp 1621261055
transform 1 0 16032 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_163
timestamp 1621261055
transform 1 0 16800 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_166
timestamp 1621261055
transform 1 0 17088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_163
timestamp 1621261055
transform 1 0 16800 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_901
timestamp 1621261055
transform 1 0 16992 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_179
timestamp 1621261055
transform 1 0 18336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_171
timestamp 1621261055
transform 1 0 17568 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_174
timestamp 1621261055
transform 1 0 17856 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_187
timestamp 1621261055
transform 1 0 19104 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_69_182
timestamp 1621261055
transform 1 0 18624 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_114
timestamp 1621261055
transform 1 0 19008 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _167_
timestamp 1621261055
transform 1 0 19200 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_912
timestamp 1621261055
transform 1 0 19680 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_191
timestamp 1621261055
transform 1 0 19488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_199
timestamp 1621261055
transform 1 0 20256 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_207
timestamp 1621261055
transform 1 0 21024 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_215
timestamp 1621261055
transform 1 0 21792 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_191
timestamp 1621261055
transform 1 0 19488 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_194
timestamp 1621261055
transform 1 0 19776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_202
timestamp 1621261055
transform 1 0 20544 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_210
timestamp 1621261055
transform 1 0 21312 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_902
timestamp 1621261055
transform 1 0 22272 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_69_219
timestamp 1621261055
transform 1 0 22176 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_221
timestamp 1621261055
transform 1 0 22368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_229
timestamp 1621261055
transform 1 0 23136 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_237
timestamp 1621261055
transform 1 0 23904 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_218
timestamp 1621261055
transform 1 0 22080 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_226
timestamp 1621261055
transform 1 0 22848 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_234
timestamp 1621261055
transform 1 0 23616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_242
timestamp 1621261055
transform 1 0 24384 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_913
timestamp 1621261055
transform 1 0 24960 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_245
timestamp 1621261055
transform 1 0 24672 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_253
timestamp 1621261055
transform 1 0 25440 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_261
timestamp 1621261055
transform 1 0 26208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_269
timestamp 1621261055
transform 1 0 26976 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_246
timestamp 1621261055
transform 1 0 24768 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_249
timestamp 1621261055
transform 1 0 25056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_257
timestamp 1621261055
transform 1 0 25824 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_265
timestamp 1621261055
transform 1 0 26592 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_903
timestamp 1621261055
transform 1 0 27552 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_273
timestamp 1621261055
transform 1 0 27360 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_276
timestamp 1621261055
transform 1 0 27648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_284
timestamp 1621261055
transform 1 0 28416 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_292
timestamp 1621261055
transform 1 0 29184 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_273
timestamp 1621261055
transform 1 0 27360 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_281
timestamp 1621261055
transform 1 0 28128 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_289
timestamp 1621261055
transform 1 0 28896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_297
timestamp 1621261055
transform 1 0 29664 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_914
timestamp 1621261055
transform 1 0 30240 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_300
timestamp 1621261055
transform 1 0 29952 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_308
timestamp 1621261055
transform 1 0 30720 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_316
timestamp 1621261055
transform 1 0 31488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_324
timestamp 1621261055
transform 1 0 32256 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_301
timestamp 1621261055
transform 1 0 30048 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_304
timestamp 1621261055
transform 1 0 30336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_312
timestamp 1621261055
transform 1 0 31104 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_320
timestamp 1621261055
transform 1 0 31872 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_904
timestamp 1621261055
transform 1 0 32832 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_328
timestamp 1621261055
transform 1 0 32640 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_331
timestamp 1621261055
transform 1 0 32928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_339
timestamp 1621261055
transform 1 0 33696 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_347
timestamp 1621261055
transform 1 0 34464 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_328
timestamp 1621261055
transform 1 0 32640 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_336
timestamp 1621261055
transform 1 0 33408 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_344
timestamp 1621261055
transform 1 0 34176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_915
timestamp 1621261055
transform 1 0 35520 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_355
timestamp 1621261055
transform 1 0 35232 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_363
timestamp 1621261055
transform 1 0 36000 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_371
timestamp 1621261055
transform 1 0 36768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_352
timestamp 1621261055
transform 1 0 34944 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_356
timestamp 1621261055
transform 1 0 35328 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_359
timestamp 1621261055
transform 1 0 35616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_367
timestamp 1621261055
transform 1 0 36384 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_375
timestamp 1621261055
transform 1 0 37152 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_70_383
timestamp 1621261055
transform 1 0 37920 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_386
timestamp 1621261055
transform 1 0 38208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_383
timestamp 1621261055
transform 1 0 37920 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_379
timestamp 1621261055
transform 1 0 37536 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_212
timestamp 1621261055
transform 1 0 38016 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_905
timestamp 1621261055
transform 1 0 38112 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _150_
timestamp 1621261055
transform 1 0 38208 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_389
timestamp 1621261055
transform 1 0 38496 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_394
timestamp 1621261055
transform 1 0 38976 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_397
timestamp 1621261055
transform 1 0 39264 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_402
timestamp 1621261055
transform 1 0 39744 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_405
timestamp 1621261055
transform 1 0 40032 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _026_
timestamp 1621261055
transform 1 0 40320 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_916
timestamp 1621261055
transform 1 0 40800 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_406
timestamp 1621261055
transform 1 0 40128 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_411
timestamp 1621261055
transform 1 0 40608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_419
timestamp 1621261055
transform 1 0 41376 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_427
timestamp 1621261055
transform 1 0 42144 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_414
timestamp 1621261055
transform 1 0 40896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_422
timestamp 1621261055
transform 1 0 41664 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_430
timestamp 1621261055
transform 1 0 42432 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_906
timestamp 1621261055
transform 1 0 43392 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_435
timestamp 1621261055
transform 1 0 42912 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_69_439
timestamp 1621261055
transform 1 0 43296 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_441
timestamp 1621261055
transform 1 0 43488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_449
timestamp 1621261055
transform 1 0 44256 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_457
timestamp 1621261055
transform 1 0 45024 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_438
timestamp 1621261055
transform 1 0 43200 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_446
timestamp 1621261055
transform 1 0 43968 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_454
timestamp 1621261055
transform 1 0 44736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_466
timestamp 1621261055
transform 1 0 45888 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_462
timestamp 1621261055
transform 1 0 45504 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_465
timestamp 1621261055
transform 1 0 45792 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_469
timestamp 1621261055
transform 1 0 46176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_473
timestamp 1621261055
transform 1 0 46560 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_917
timestamp 1621261055
transform 1 0 46080 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_485
timestamp 1621261055
transform 1 0 47712 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_477
timestamp 1621261055
transform 1 0 46944 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_483
timestamp 1621261055
transform 1 0 47520 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_481
timestamp 1621261055
transform 1 0 47328 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_197
timestamp 1621261055
transform -1 0 47808 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _137_
timestamp 1621261055
transform -1 0 48096 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_493
timestamp 1621261055
transform 1 0 48480 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_493
timestamp 1621261055
transform 1 0 48480 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_489
timestamp 1621261055
transform 1 0 48096 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_501
timestamp 1621261055
transform 1 0 49248 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_496
timestamp 1621261055
transform 1 0 48768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_907
timestamp 1621261055
transform 1 0 48672 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_509
timestamp 1621261055
transform 1 0 50016 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_512
timestamp 1621261055
transform 1 0 50304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_504
timestamp 1621261055
transform 1 0 49536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_101
timestamp 1621261055
transform 1 0 50208 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _156_
timestamp 1621261055
transform 1 0 50400 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_520
timestamp 1621261055
transform 1 0 51072 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_516
timestamp 1621261055
transform 1 0 50688 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_520
timestamp 1621261055
transform 1 0 51072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_524
timestamp 1621261055
transform 1 0 51456 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_70_522
timestamp 1621261055
transform 1 0 51264 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_528
timestamp 1621261055
transform 1 0 51840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_918
timestamp 1621261055
transform 1 0 51360 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _100_
timestamp 1621261055
transform 1 0 51840 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_539
timestamp 1621261055
transform 1 0 52896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_531
timestamp 1621261055
transform 1 0 52128 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_536
timestamp 1621261055
transform 1 0 52608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_908
timestamp 1621261055
transform 1 0 53952 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_69_544
timestamp 1621261055
transform 1 0 53376 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_548
timestamp 1621261055
transform 1 0 53760 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_551
timestamp 1621261055
transform 1 0 54048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_559
timestamp 1621261055
transform 1 0 54816 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_567
timestamp 1621261055
transform 1 0 55584 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_547
timestamp 1621261055
transform 1 0 53664 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_555
timestamp 1621261055
transform 1 0 54432 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_563
timestamp 1621261055
transform 1 0 55200 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_919
timestamp 1621261055
transform 1 0 56640 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_575
timestamp 1621261055
transform 1 0 56352 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_583
timestamp 1621261055
transform 1 0 57120 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_591
timestamp 1621261055
transform 1 0 57888 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_70_571
timestamp 1621261055
transform 1 0 55968 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_575
timestamp 1621261055
transform 1 0 56352 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_70_577
timestamp 1621261055
transform 1 0 56544 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_579
timestamp 1621261055
transform 1 0 56736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_587
timestamp 1621261055
transform 1 0 57504 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_139
timestamp 1621261055
transform -1 0 58848 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_141
timestamp 1621261055
transform -1 0 58848 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_595
timestamp 1621261055
transform 1 0 58272 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_595
timestamp 1621261055
transform 1 0 58272 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_142
timestamp 1621261055
transform 1 0 1152 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_4
timestamp 1621261055
transform 1 0 1536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_12
timestamp 1621261055
transform 1 0 2304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_20
timestamp 1621261055
transform 1 0 3072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_28
timestamp 1621261055
transform 1 0 3840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_36
timestamp 1621261055
transform 1 0 4608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_44
timestamp 1621261055
transform 1 0 5376 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_52
timestamp 1621261055
transform 1 0 6144 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_54
timestamp 1621261055
transform 1 0 6336 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_920
timestamp 1621261055
transform 1 0 6432 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_56
timestamp 1621261055
transform 1 0 6528 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_64
timestamp 1621261055
transform 1 0 7296 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_72
timestamp 1621261055
transform 1 0 8064 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_80
timestamp 1621261055
transform 1 0 8832 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_88
timestamp 1621261055
transform 1 0 9600 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_96
timestamp 1621261055
transform 1 0 10368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_104
timestamp 1621261055
transform 1 0 11136 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_108
timestamp 1621261055
transform 1 0 11520 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_921
timestamp 1621261055
transform 1 0 11712 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_111
timestamp 1621261055
transform 1 0 11808 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_119
timestamp 1621261055
transform 1 0 12576 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_127
timestamp 1621261055
transform 1 0 13344 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_135
timestamp 1621261055
transform 1 0 14112 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_143
timestamp 1621261055
transform 1 0 14880 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_151
timestamp 1621261055
transform 1 0 15648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_159
timestamp 1621261055
transform 1 0 16416 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_922
timestamp 1621261055
transform 1 0 16992 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_163
timestamp 1621261055
transform 1 0 16800 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_166
timestamp 1621261055
transform 1 0 17088 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_174
timestamp 1621261055
transform 1 0 17856 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_182
timestamp 1621261055
transform 1 0 18624 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_190
timestamp 1621261055
transform 1 0 19392 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_198
timestamp 1621261055
transform 1 0 20160 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_206
timestamp 1621261055
transform 1 0 20928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_214
timestamp 1621261055
transform 1 0 21696 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_923
timestamp 1621261055
transform 1 0 22272 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_218
timestamp 1621261055
transform 1 0 22080 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_221
timestamp 1621261055
transform 1 0 22368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_229
timestamp 1621261055
transform 1 0 23136 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_237
timestamp 1621261055
transform 1 0 23904 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_245
timestamp 1621261055
transform 1 0 24672 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_253
timestamp 1621261055
transform 1 0 25440 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_261
timestamp 1621261055
transform 1 0 26208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_269
timestamp 1621261055
transform 1 0 26976 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_924
timestamp 1621261055
transform 1 0 27552 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_118
timestamp 1621261055
transform 1 0 29664 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_273
timestamp 1621261055
transform 1 0 27360 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_276
timestamp 1621261055
transform 1 0 27648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_284
timestamp 1621261055
transform 1 0 28416 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_292
timestamp 1621261055
transform 1 0 29184 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_71_296
timestamp 1621261055
transform 1 0 29568 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _171_
timestamp 1621261055
transform 1 0 29856 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_71_302
timestamp 1621261055
transform 1 0 30144 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_310
timestamp 1621261055
transform 1 0 30912 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_318
timestamp 1621261055
transform 1 0 31680 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_925
timestamp 1621261055
transform 1 0 32832 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_326
timestamp 1621261055
transform 1 0 32448 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_331
timestamp 1621261055
transform 1 0 32928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_339
timestamp 1621261055
transform 1 0 33696 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_347
timestamp 1621261055
transform 1 0 34464 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_355
timestamp 1621261055
transform 1 0 35232 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_363
timestamp 1621261055
transform 1 0 36000 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_371
timestamp 1621261055
transform 1 0 36768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_926
timestamp 1621261055
transform 1 0 38112 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_379
timestamp 1621261055
transform 1 0 37536 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_383
timestamp 1621261055
transform 1 0 37920 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_386
timestamp 1621261055
transform 1 0 38208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_394
timestamp 1621261055
transform 1 0 38976 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_402
timestamp 1621261055
transform 1 0 39744 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_410
timestamp 1621261055
transform 1 0 40512 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_418
timestamp 1621261055
transform 1 0 41280 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_426
timestamp 1621261055
transform 1 0 42048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_927
timestamp 1621261055
transform 1 0 43392 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_434
timestamp 1621261055
transform 1 0 42816 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_438
timestamp 1621261055
transform 1 0 43200 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_441
timestamp 1621261055
transform 1 0 43488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_449
timestamp 1621261055
transform 1 0 44256 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_457
timestamp 1621261055
transform 1 0 45024 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_465
timestamp 1621261055
transform 1 0 45792 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_473
timestamp 1621261055
transform 1 0 46560 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_481
timestamp 1621261055
transform 1 0 47328 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _066_
timestamp 1621261055
transform -1 0 49440 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_928
timestamp 1621261055
transform 1 0 48672 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_111
timestamp 1621261055
transform -1 0 49152 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_71_489
timestamp 1621261055
transform 1 0 48096 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_493
timestamp 1621261055
transform 1 0 48480 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_496
timestamp 1621261055
transform 1 0 48768 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_503
timestamp 1621261055
transform 1 0 49440 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_511
timestamp 1621261055
transform 1 0 50208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_519
timestamp 1621261055
transform 1 0 50976 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_527
timestamp 1621261055
transform 1 0 51744 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_535
timestamp 1621261055
transform 1 0 52512 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_929
timestamp 1621261055
transform 1 0 53952 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_543
timestamp 1621261055
transform 1 0 53280 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_547
timestamp 1621261055
transform 1 0 53664 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_549
timestamp 1621261055
transform 1 0 53856 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_551
timestamp 1621261055
transform 1 0 54048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_559
timestamp 1621261055
transform 1 0 54816 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_567
timestamp 1621261055
transform 1 0 55584 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _101_
timestamp 1621261055
transform -1 0 58080 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_163
timestamp 1621261055
transform -1 0 57792 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_575
timestamp 1621261055
transform 1 0 56352 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_583
timestamp 1621261055
transform 1 0 57120 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_71_587
timestamp 1621261055
transform 1 0 57504 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_593
timestamp 1621261055
transform 1 0 58080 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_143
timestamp 1621261055
transform -1 0 58848 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_144
timestamp 1621261055
transform 1 0 1152 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_72_4
timestamp 1621261055
transform 1 0 1536 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_12
timestamp 1621261055
transform 1 0 2304 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_20
timestamp 1621261055
transform 1 0 3072 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_930
timestamp 1621261055
transform 1 0 3840 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_29
timestamp 1621261055
transform 1 0 3936 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_37
timestamp 1621261055
transform 1 0 4704 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_45
timestamp 1621261055
transform 1 0 5472 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_53
timestamp 1621261055
transform 1 0 6240 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_61
timestamp 1621261055
transform 1 0 7008 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_69
timestamp 1621261055
transform 1 0 7776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_77
timestamp 1621261055
transform 1 0 8544 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_81
timestamp 1621261055
transform 1 0 8928 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_931
timestamp 1621261055
transform 1 0 9120 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_84
timestamp 1621261055
transform 1 0 9216 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_92
timestamp 1621261055
transform 1 0 9984 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_100
timestamp 1621261055
transform 1 0 10752 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_108
timestamp 1621261055
transform 1 0 11520 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_116
timestamp 1621261055
transform 1 0 12288 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_124
timestamp 1621261055
transform 1 0 13056 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_132
timestamp 1621261055
transform 1 0 13824 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_932
timestamp 1621261055
transform 1 0 14400 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_136
timestamp 1621261055
transform 1 0 14208 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_139
timestamp 1621261055
transform 1 0 14496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_147
timestamp 1621261055
transform 1 0 15264 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_155
timestamp 1621261055
transform 1 0 16032 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_163
timestamp 1621261055
transform 1 0 16800 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_171
timestamp 1621261055
transform 1 0 17568 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_179
timestamp 1621261055
transform 1 0 18336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_187
timestamp 1621261055
transform 1 0 19104 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_933
timestamp 1621261055
transform 1 0 19680 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_191
timestamp 1621261055
transform 1 0 19488 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_194
timestamp 1621261055
transform 1 0 19776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_202
timestamp 1621261055
transform 1 0 20544 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_210
timestamp 1621261055
transform 1 0 21312 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_218
timestamp 1621261055
transform 1 0 22080 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_226
timestamp 1621261055
transform 1 0 22848 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_234
timestamp 1621261055
transform 1 0 23616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_242
timestamp 1621261055
transform 1 0 24384 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _134_
timestamp 1621261055
transform 1 0 25440 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_934
timestamp 1621261055
transform 1 0 24960 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_193
timestamp 1621261055
transform 1 0 25248 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_246
timestamp 1621261055
transform 1 0 24768 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_249
timestamp 1621261055
transform 1 0 25056 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_256
timestamp 1621261055
transform 1 0 25728 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_264
timestamp 1621261055
transform 1 0 26496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_272
timestamp 1621261055
transform 1 0 27264 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_280
timestamp 1621261055
transform 1 0 28032 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_288
timestamp 1621261055
transform 1 0 28800 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_296
timestamp 1621261055
transform 1 0 29568 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _082_
timestamp 1621261055
transform -1 0 31968 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_935
timestamp 1621261055
transform 1 0 30240 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_147
timestamp 1621261055
transform -1 0 31680 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_300
timestamp 1621261055
transform 1 0 29952 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_72_302
timestamp 1621261055
transform 1 0 30144 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_304
timestamp 1621261055
transform 1 0 30336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_312
timestamp 1621261055
transform 1 0 31104 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_72_321
timestamp 1621261055
transform 1 0 31968 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_329
timestamp 1621261055
transform 1 0 32736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_337
timestamp 1621261055
transform 1 0 33504 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_345
timestamp 1621261055
transform 1 0 34272 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_936
timestamp 1621261055
transform 1 0 35520 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_353
timestamp 1621261055
transform 1 0 35040 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_72_357
timestamp 1621261055
transform 1 0 35424 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_359
timestamp 1621261055
transform 1 0 35616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_367
timestamp 1621261055
transform 1 0 36384 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_375
timestamp 1621261055
transform 1 0 37152 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_383
timestamp 1621261055
transform 1 0 37920 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_391
timestamp 1621261055
transform 1 0 38688 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_399
timestamp 1621261055
transform 1 0 39456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_937
timestamp 1621261055
transform 1 0 40800 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_407
timestamp 1621261055
transform 1 0 40224 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_411
timestamp 1621261055
transform 1 0 40608 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_414
timestamp 1621261055
transform 1 0 40896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_422
timestamp 1621261055
transform 1 0 41664 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_430
timestamp 1621261055
transform 1 0 42432 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_438
timestamp 1621261055
transform 1 0 43200 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_446
timestamp 1621261055
transform 1 0 43968 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_454
timestamp 1621261055
transform 1 0 44736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_938
timestamp 1621261055
transform 1 0 46080 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_462
timestamp 1621261055
transform 1 0 45504 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_466
timestamp 1621261055
transform 1 0 45888 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_469
timestamp 1621261055
transform 1 0 46176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_477
timestamp 1621261055
transform 1 0 46944 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_485
timestamp 1621261055
transform 1 0 47712 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_493
timestamp 1621261055
transform 1 0 48480 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_501
timestamp 1621261055
transform 1 0 49248 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_509
timestamp 1621261055
transform 1 0 50016 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_939
timestamp 1621261055
transform 1 0 51360 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_517
timestamp 1621261055
transform 1 0 50784 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_521
timestamp 1621261055
transform 1 0 51168 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_524
timestamp 1621261055
transform 1 0 51456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_532
timestamp 1621261055
transform 1 0 52224 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_540
timestamp 1621261055
transform 1 0 52992 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_548
timestamp 1621261055
transform 1 0 53760 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_556
timestamp 1621261055
transform 1 0 54528 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_564
timestamp 1621261055
transform 1 0 55296 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_940
timestamp 1621261055
transform 1 0 56640 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_572
timestamp 1621261055
transform 1 0 56064 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_576
timestamp 1621261055
transform 1 0 56448 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_579
timestamp 1621261055
transform 1 0 56736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_587
timestamp 1621261055
transform 1 0 57504 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_145
timestamp 1621261055
transform -1 0 58848 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_595
timestamp 1621261055
transform 1 0 58272 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _104_
timestamp 1621261055
transform 1 0 1728 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_146
timestamp 1621261055
transform 1 0 1152 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_165
timestamp 1621261055
transform 1 0 1536 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_9
timestamp 1621261055
transform 1 0 2016 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_17
timestamp 1621261055
transform 1 0 2784 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_25
timestamp 1621261055
transform 1 0 3552 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _162_
timestamp 1621261055
transform 1 0 5760 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_107
timestamp 1621261055
transform 1 0 5568 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_33
timestamp 1621261055
transform 1 0 4320 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_41
timestamp 1621261055
transform 1 0 5088 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_73_45
timestamp 1621261055
transform 1 0 5472 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_51
timestamp 1621261055
transform 1 0 6048 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_941
timestamp 1621261055
transform 1 0 6432 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_56
timestamp 1621261055
transform 1 0 6528 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_64
timestamp 1621261055
transform 1 0 7296 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_72
timestamp 1621261055
transform 1 0 8064 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_80
timestamp 1621261055
transform 1 0 8832 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_88
timestamp 1621261055
transform 1 0 9600 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_96
timestamp 1621261055
transform 1 0 10368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_104
timestamp 1621261055
transform 1 0 11136 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_108
timestamp 1621261055
transform 1 0 11520 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_942
timestamp 1621261055
transform 1 0 11712 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_111
timestamp 1621261055
transform 1 0 11808 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_119
timestamp 1621261055
transform 1 0 12576 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_127
timestamp 1621261055
transform 1 0 13344 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_135
timestamp 1621261055
transform 1 0 14112 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_143
timestamp 1621261055
transform 1 0 14880 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_151
timestamp 1621261055
transform 1 0 15648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_159
timestamp 1621261055
transform 1 0 16416 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_943
timestamp 1621261055
transform 1 0 16992 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_163
timestamp 1621261055
transform 1 0 16800 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_166
timestamp 1621261055
transform 1 0 17088 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_174
timestamp 1621261055
transform 1 0 17856 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_182
timestamp 1621261055
transform 1 0 18624 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _151_
timestamp 1621261055
transform 1 0 19872 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_214
timestamp 1621261055
transform 1 0 19680 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_190
timestamp 1621261055
transform 1 0 19392 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_192
timestamp 1621261055
transform 1 0 19584 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_198
timestamp 1621261055
transform 1 0 20160 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_206
timestamp 1621261055
transform 1 0 20928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_214
timestamp 1621261055
transform 1 0 21696 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_944
timestamp 1621261055
transform 1 0 22272 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_218
timestamp 1621261055
transform 1 0 22080 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_221
timestamp 1621261055
transform 1 0 22368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_229
timestamp 1621261055
transform 1 0 23136 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_237
timestamp 1621261055
transform 1 0 23904 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_245
timestamp 1621261055
transform 1 0 24672 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_253
timestamp 1621261055
transform 1 0 25440 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_261
timestamp 1621261055
transform 1 0 26208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_269
timestamp 1621261055
transform 1 0 26976 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_945
timestamp 1621261055
transform 1 0 27552 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_273
timestamp 1621261055
transform 1 0 27360 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_276
timestamp 1621261055
transform 1 0 27648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_284
timestamp 1621261055
transform 1 0 28416 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_292
timestamp 1621261055
transform 1 0 29184 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_300
timestamp 1621261055
transform 1 0 29952 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_308
timestamp 1621261055
transform 1 0 30720 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_316
timestamp 1621261055
transform 1 0 31488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_324
timestamp 1621261055
transform 1 0 32256 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_946
timestamp 1621261055
transform 1 0 32832 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_328
timestamp 1621261055
transform 1 0 32640 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_331
timestamp 1621261055
transform 1 0 32928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_339
timestamp 1621261055
transform 1 0 33696 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_347
timestamp 1621261055
transform 1 0 34464 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_355
timestamp 1621261055
transform 1 0 35232 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_363
timestamp 1621261055
transform 1 0 36000 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_371
timestamp 1621261055
transform 1 0 36768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_947
timestamp 1621261055
transform 1 0 38112 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_379
timestamp 1621261055
transform 1 0 37536 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_383
timestamp 1621261055
transform 1 0 37920 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_386
timestamp 1621261055
transform 1 0 38208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_394
timestamp 1621261055
transform 1 0 38976 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_402
timestamp 1621261055
transform 1 0 39744 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_410
timestamp 1621261055
transform 1 0 40512 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_418
timestamp 1621261055
transform 1 0 41280 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_426
timestamp 1621261055
transform 1 0 42048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_948
timestamp 1621261055
transform 1 0 43392 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_434
timestamp 1621261055
transform 1 0 42816 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_438
timestamp 1621261055
transform 1 0 43200 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_441
timestamp 1621261055
transform 1 0 43488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_449
timestamp 1621261055
transform 1 0 44256 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_457
timestamp 1621261055
transform 1 0 45024 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_465
timestamp 1621261055
transform 1 0 45792 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_473
timestamp 1621261055
transform 1 0 46560 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_481
timestamp 1621261055
transform 1 0 47328 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_949
timestamp 1621261055
transform 1 0 48672 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_489
timestamp 1621261055
transform 1 0 48096 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_493
timestamp 1621261055
transform 1 0 48480 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_496
timestamp 1621261055
transform 1 0 48768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_504
timestamp 1621261055
transform 1 0 49536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_512
timestamp 1621261055
transform 1 0 50304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_520
timestamp 1621261055
transform 1 0 51072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_528
timestamp 1621261055
transform 1 0 51840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_536
timestamp 1621261055
transform 1 0 52608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_950
timestamp 1621261055
transform 1 0 53952 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_544
timestamp 1621261055
transform 1 0 53376 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_548
timestamp 1621261055
transform 1 0 53760 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_551
timestamp 1621261055
transform 1 0 54048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_559
timestamp 1621261055
transform 1 0 54816 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_567
timestamp 1621261055
transform 1 0 55584 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_575
timestamp 1621261055
transform 1 0 56352 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_583
timestamp 1621261055
transform 1 0 57120 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_591
timestamp 1621261055
transform 1 0 57888 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_147
timestamp 1621261055
transform -1 0 58848 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_595
timestamp 1621261055
transform 1 0 58272 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_148
timestamp 1621261055
transform 1 0 1152 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_4
timestamp 1621261055
transform 1 0 1536 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_12
timestamp 1621261055
transform 1 0 2304 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_20
timestamp 1621261055
transform 1 0 3072 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_951
timestamp 1621261055
transform 1 0 3840 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_29
timestamp 1621261055
transform 1 0 3936 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_37
timestamp 1621261055
transform 1 0 4704 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_45
timestamp 1621261055
transform 1 0 5472 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_53
timestamp 1621261055
transform 1 0 6240 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_61
timestamp 1621261055
transform 1 0 7008 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_69
timestamp 1621261055
transform 1 0 7776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_77
timestamp 1621261055
transform 1 0 8544 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_81
timestamp 1621261055
transform 1 0 8928 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_952
timestamp 1621261055
transform 1 0 9120 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_84
timestamp 1621261055
transform 1 0 9216 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_92
timestamp 1621261055
transform 1 0 9984 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_100
timestamp 1621261055
transform 1 0 10752 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_108
timestamp 1621261055
transform 1 0 11520 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_116
timestamp 1621261055
transform 1 0 12288 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_124
timestamp 1621261055
transform 1 0 13056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_132
timestamp 1621261055
transform 1 0 13824 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_953
timestamp 1621261055
transform 1 0 14400 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_136
timestamp 1621261055
transform 1 0 14208 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_139
timestamp 1621261055
transform 1 0 14496 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_147
timestamp 1621261055
transform 1 0 15264 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_155
timestamp 1621261055
transform 1 0 16032 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_163
timestamp 1621261055
transform 1 0 16800 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_171
timestamp 1621261055
transform 1 0 17568 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_179
timestamp 1621261055
transform 1 0 18336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_187
timestamp 1621261055
transform 1 0 19104 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_954
timestamp 1621261055
transform 1 0 19680 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_191
timestamp 1621261055
transform 1 0 19488 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_194
timestamp 1621261055
transform 1 0 19776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_202
timestamp 1621261055
transform 1 0 20544 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_210
timestamp 1621261055
transform 1 0 21312 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_218
timestamp 1621261055
transform 1 0 22080 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_226
timestamp 1621261055
transform 1 0 22848 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_234
timestamp 1621261055
transform 1 0 23616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_242
timestamp 1621261055
transform 1 0 24384 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_955
timestamp 1621261055
transform 1 0 24960 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_246
timestamp 1621261055
transform 1 0 24768 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_249
timestamp 1621261055
transform 1 0 25056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_257
timestamp 1621261055
transform 1 0 25824 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_265
timestamp 1621261055
transform 1 0 26592 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_273
timestamp 1621261055
transform 1 0 27360 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_281
timestamp 1621261055
transform 1 0 28128 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_289
timestamp 1621261055
transform 1 0 28896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_297
timestamp 1621261055
transform 1 0 29664 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_956
timestamp 1621261055
transform 1 0 30240 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_301
timestamp 1621261055
transform 1 0 30048 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_304
timestamp 1621261055
transform 1 0 30336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_312
timestamp 1621261055
transform 1 0 31104 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_320
timestamp 1621261055
transform 1 0 31872 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_328
timestamp 1621261055
transform 1 0 32640 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_336
timestamp 1621261055
transform 1 0 33408 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_344
timestamp 1621261055
transform 1 0 34176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _009_
timestamp 1621261055
transform 1 0 37056 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_957
timestamp 1621261055
transform 1 0 35520 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_352
timestamp 1621261055
transform 1 0 34944 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_356
timestamp 1621261055
transform 1 0 35328 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_359
timestamp 1621261055
transform 1 0 35616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_367
timestamp 1621261055
transform 1 0 36384 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_371
timestamp 1621261055
transform 1 0 36768 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_74_373
timestamp 1621261055
transform 1 0 36960 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_377
timestamp 1621261055
transform 1 0 37344 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_385
timestamp 1621261055
transform 1 0 38112 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_393
timestamp 1621261055
transform 1 0 38880 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_401
timestamp 1621261055
transform 1 0 39648 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_958
timestamp 1621261055
transform 1 0 40800 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_409
timestamp 1621261055
transform 1 0 40416 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_414
timestamp 1621261055
transform 1 0 40896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_422
timestamp 1621261055
transform 1 0 41664 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_430
timestamp 1621261055
transform 1 0 42432 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _072_
timestamp 1621261055
transform -1 0 43296 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_137
timestamp 1621261055
transform -1 0 43008 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_439
timestamp 1621261055
transform 1 0 43296 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_447
timestamp 1621261055
transform 1 0 44064 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_455
timestamp 1621261055
transform 1 0 44832 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_959
timestamp 1621261055
transform 1 0 46080 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_463
timestamp 1621261055
transform 1 0 45600 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_74_467
timestamp 1621261055
transform 1 0 45984 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_469
timestamp 1621261055
transform 1 0 46176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_477
timestamp 1621261055
transform 1 0 46944 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_485
timestamp 1621261055
transform 1 0 47712 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_493
timestamp 1621261055
transform 1 0 48480 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_501
timestamp 1621261055
transform 1 0 49248 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_509
timestamp 1621261055
transform 1 0 50016 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_960
timestamp 1621261055
transform 1 0 51360 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_517
timestamp 1621261055
transform 1 0 50784 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_521
timestamp 1621261055
transform 1 0 51168 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_524
timestamp 1621261055
transform 1 0 51456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_532
timestamp 1621261055
transform 1 0 52224 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_540
timestamp 1621261055
transform 1 0 52992 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_548
timestamp 1621261055
transform 1 0 53760 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_556
timestamp 1621261055
transform 1 0 54528 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_564
timestamp 1621261055
transform 1 0 55296 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_961
timestamp 1621261055
transform 1 0 56640 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_74_572
timestamp 1621261055
transform 1 0 56064 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_576
timestamp 1621261055
transform 1 0 56448 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_579
timestamp 1621261055
transform 1 0 56736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_587
timestamp 1621261055
transform 1 0 57504 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_149
timestamp 1621261055
transform -1 0 58848 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_595
timestamp 1621261055
transform 1 0 58272 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_150
timestamp 1621261055
transform 1 0 1152 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_75_4
timestamp 1621261055
transform 1 0 1536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_12
timestamp 1621261055
transform 1 0 2304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_20
timestamp 1621261055
transform 1 0 3072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_28
timestamp 1621261055
transform 1 0 3840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_36
timestamp 1621261055
transform 1 0 4608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_44
timestamp 1621261055
transform 1 0 5376 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_52
timestamp 1621261055
transform 1 0 6144 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_54
timestamp 1621261055
transform 1 0 6336 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_962
timestamp 1621261055
transform 1 0 6432 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_56
timestamp 1621261055
transform 1 0 6528 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_64
timestamp 1621261055
transform 1 0 7296 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_72
timestamp 1621261055
transform 1 0 8064 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_80
timestamp 1621261055
transform 1 0 8832 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_88
timestamp 1621261055
transform 1 0 9600 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_96
timestamp 1621261055
transform 1 0 10368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_104
timestamp 1621261055
transform 1 0 11136 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_108
timestamp 1621261055
transform 1 0 11520 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_963
timestamp 1621261055
transform 1 0 11712 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_111
timestamp 1621261055
transform 1 0 11808 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_119
timestamp 1621261055
transform 1 0 12576 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_127
timestamp 1621261055
transform 1 0 13344 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_135
timestamp 1621261055
transform 1 0 14112 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_143
timestamp 1621261055
transform 1 0 14880 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_151
timestamp 1621261055
transform 1 0 15648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_159
timestamp 1621261055
transform 1 0 16416 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_964
timestamp 1621261055
transform 1 0 16992 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_163
timestamp 1621261055
transform 1 0 16800 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_166
timestamp 1621261055
transform 1 0 17088 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_174
timestamp 1621261055
transform 1 0 17856 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_182
timestamp 1621261055
transform 1 0 18624 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _004_
timestamp 1621261055
transform 1 0 21312 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_75_190
timestamp 1621261055
transform 1 0 19392 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_198
timestamp 1621261055
transform 1 0 20160 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_206
timestamp 1621261055
transform 1 0 20928 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_75_213
timestamp 1621261055
transform 1 0 21600 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _078_
timestamp 1621261055
transform -1 0 24480 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_965
timestamp 1621261055
transform 1 0 22272 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_143
timestamp 1621261055
transform -1 0 24192 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_217
timestamp 1621261055
transform 1 0 21984 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_219
timestamp 1621261055
transform 1 0 22176 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_221
timestamp 1621261055
transform 1 0 22368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_229
timestamp 1621261055
transform 1 0 23136 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_75_237
timestamp 1621261055
transform 1 0 23904 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_243
timestamp 1621261055
transform 1 0 24480 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_251
timestamp 1621261055
transform 1 0 25248 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_259
timestamp 1621261055
transform 1 0 26016 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_267
timestamp 1621261055
transform 1 0 26784 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_966
timestamp 1621261055
transform 1 0 27552 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_276
timestamp 1621261055
transform 1 0 27648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_284
timestamp 1621261055
transform 1 0 28416 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_292
timestamp 1621261055
transform 1 0 29184 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_300
timestamp 1621261055
transform 1 0 29952 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_308
timestamp 1621261055
transform 1 0 30720 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_316
timestamp 1621261055
transform 1 0 31488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_324
timestamp 1621261055
transform 1 0 32256 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_967
timestamp 1621261055
transform 1 0 32832 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_328
timestamp 1621261055
transform 1 0 32640 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_331
timestamp 1621261055
transform 1 0 32928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_339
timestamp 1621261055
transform 1 0 33696 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_347
timestamp 1621261055
transform 1 0 34464 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_355
timestamp 1621261055
transform 1 0 35232 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_363
timestamp 1621261055
transform 1 0 36000 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_371
timestamp 1621261055
transform 1 0 36768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_968
timestamp 1621261055
transform 1 0 38112 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_379
timestamp 1621261055
transform 1 0 37536 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_383
timestamp 1621261055
transform 1 0 37920 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_386
timestamp 1621261055
transform 1 0 38208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_394
timestamp 1621261055
transform 1 0 38976 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_402
timestamp 1621261055
transform 1 0 39744 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _148_
timestamp 1621261055
transform 1 0 40896 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_209
timestamp 1621261055
transform 1 0 40704 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_410
timestamp 1621261055
transform 1 0 40512 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_417
timestamp 1621261055
transform 1 0 41184 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_425
timestamp 1621261055
transform 1 0 41952 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_969
timestamp 1621261055
transform 1 0 43392 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_433
timestamp 1621261055
transform 1 0 42720 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_437
timestamp 1621261055
transform 1 0 43104 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_439
timestamp 1621261055
transform 1 0 43296 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_441
timestamp 1621261055
transform 1 0 43488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_449
timestamp 1621261055
transform 1 0 44256 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_457
timestamp 1621261055
transform 1 0 45024 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_465
timestamp 1621261055
transform 1 0 45792 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_473
timestamp 1621261055
transform 1 0 46560 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_481
timestamp 1621261055
transform 1 0 47328 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_970
timestamp 1621261055
transform 1 0 48672 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_489
timestamp 1621261055
transform 1 0 48096 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_493
timestamp 1621261055
transform 1 0 48480 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_496
timestamp 1621261055
transform 1 0 48768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_504
timestamp 1621261055
transform 1 0 49536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_512
timestamp 1621261055
transform 1 0 50304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_520
timestamp 1621261055
transform 1 0 51072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_528
timestamp 1621261055
transform 1 0 51840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_536
timestamp 1621261055
transform 1 0 52608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_971
timestamp 1621261055
transform 1 0 53952 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_544
timestamp 1621261055
transform 1 0 53376 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_548
timestamp 1621261055
transform 1 0 53760 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_551
timestamp 1621261055
transform 1 0 54048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_559
timestamp 1621261055
transform 1 0 54816 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_567
timestamp 1621261055
transform 1 0 55584 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_575
timestamp 1621261055
transform 1 0 56352 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_583
timestamp 1621261055
transform 1 0 57120 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_591
timestamp 1621261055
transform 1 0 57888 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_151
timestamp 1621261055
transform -1 0 58848 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_595
timestamp 1621261055
transform 1 0 58272 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_152
timestamp 1621261055
transform 1 0 1152 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_76_4
timestamp 1621261055
transform 1 0 1536 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_12
timestamp 1621261055
transform 1 0 2304 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_20
timestamp 1621261055
transform 1 0 3072 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_972
timestamp 1621261055
transform 1 0 3840 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_29
timestamp 1621261055
transform 1 0 3936 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_37
timestamp 1621261055
transform 1 0 4704 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_45
timestamp 1621261055
transform 1 0 5472 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_53
timestamp 1621261055
transform 1 0 6240 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_61
timestamp 1621261055
transform 1 0 7008 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_69
timestamp 1621261055
transform 1 0 7776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_77
timestamp 1621261055
transform 1 0 8544 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_81
timestamp 1621261055
transform 1 0 8928 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_973
timestamp 1621261055
transform 1 0 9120 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_84
timestamp 1621261055
transform 1 0 9216 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_92
timestamp 1621261055
transform 1 0 9984 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_100
timestamp 1621261055
transform 1 0 10752 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_108
timestamp 1621261055
transform 1 0 11520 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_116
timestamp 1621261055
transform 1 0 12288 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_124
timestamp 1621261055
transform 1 0 13056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_132
timestamp 1621261055
transform 1 0 13824 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_974
timestamp 1621261055
transform 1 0 14400 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_136
timestamp 1621261055
transform 1 0 14208 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_139
timestamp 1621261055
transform 1 0 14496 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_147
timestamp 1621261055
transform 1 0 15264 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_155
timestamp 1621261055
transform 1 0 16032 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_163
timestamp 1621261055
transform 1 0 16800 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_171
timestamp 1621261055
transform 1 0 17568 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_179
timestamp 1621261055
transform 1 0 18336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_187
timestamp 1621261055
transform 1 0 19104 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_975
timestamp 1621261055
transform 1 0 19680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_191
timestamp 1621261055
transform 1 0 19488 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_194
timestamp 1621261055
transform 1 0 19776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_202
timestamp 1621261055
transform 1 0 20544 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_210
timestamp 1621261055
transform 1 0 21312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_218
timestamp 1621261055
transform 1 0 22080 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_226
timestamp 1621261055
transform 1 0 22848 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_234
timestamp 1621261055
transform 1 0 23616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_242
timestamp 1621261055
transform 1 0 24384 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _189_
timestamp 1621261055
transform -1 0 27264 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_976
timestamp 1621261055
transform 1 0 24960 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_249
timestamp 1621261055
transform -1 0 26976 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_246
timestamp 1621261055
transform 1 0 24768 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_249
timestamp 1621261055
transform 1 0 25056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_257
timestamp 1621261055
transform 1 0 25824 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_265
timestamp 1621261055
transform 1 0 26592 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_272
timestamp 1621261055
transform 1 0 27264 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_280
timestamp 1621261055
transform 1 0 28032 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_288
timestamp 1621261055
transform 1 0 28800 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_296
timestamp 1621261055
transform 1 0 29568 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_977
timestamp 1621261055
transform 1 0 30240 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_300
timestamp 1621261055
transform 1 0 29952 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_76_302
timestamp 1621261055
transform 1 0 30144 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_304
timestamp 1621261055
transform 1 0 30336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_312
timestamp 1621261055
transform 1 0 31104 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_320
timestamp 1621261055
transform 1 0 31872 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_328
timestamp 1621261055
transform 1 0 32640 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_336
timestamp 1621261055
transform 1 0 33408 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_344
timestamp 1621261055
transform 1 0 34176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_978
timestamp 1621261055
transform 1 0 35520 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_352
timestamp 1621261055
transform 1 0 34944 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_356
timestamp 1621261055
transform 1 0 35328 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_359
timestamp 1621261055
transform 1 0 35616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_367
timestamp 1621261055
transform 1 0 36384 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_375
timestamp 1621261055
transform 1 0 37152 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_383
timestamp 1621261055
transform 1 0 37920 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_391
timestamp 1621261055
transform 1 0 38688 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_399
timestamp 1621261055
transform 1 0 39456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_979
timestamp 1621261055
transform 1 0 40800 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_407
timestamp 1621261055
transform 1 0 40224 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_411
timestamp 1621261055
transform 1 0 40608 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_414
timestamp 1621261055
transform 1 0 40896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_422
timestamp 1621261055
transform 1 0 41664 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_430
timestamp 1621261055
transform 1 0 42432 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_438
timestamp 1621261055
transform 1 0 43200 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_446
timestamp 1621261055
transform 1 0 43968 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_454
timestamp 1621261055
transform 1 0 44736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_980
timestamp 1621261055
transform 1 0 46080 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_462
timestamp 1621261055
transform 1 0 45504 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_466
timestamp 1621261055
transform 1 0 45888 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_469
timestamp 1621261055
transform 1 0 46176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_477
timestamp 1621261055
transform 1 0 46944 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_485
timestamp 1621261055
transform 1 0 47712 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_493
timestamp 1621261055
transform 1 0 48480 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_501
timestamp 1621261055
transform 1 0 49248 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_509
timestamp 1621261055
transform 1 0 50016 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_981
timestamp 1621261055
transform 1 0 51360 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_76_517
timestamp 1621261055
transform 1 0 50784 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_521
timestamp 1621261055
transform 1 0 51168 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_524
timestamp 1621261055
transform 1 0 51456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_532
timestamp 1621261055
transform 1 0 52224 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_540
timestamp 1621261055
transform 1 0 52992 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_548
timestamp 1621261055
transform 1 0 53760 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_556
timestamp 1621261055
transform 1 0 54528 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_564
timestamp 1621261055
transform 1 0 55296 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_982
timestamp 1621261055
transform 1 0 56640 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output436
timestamp 1621261055
transform -1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_88
timestamp 1621261055
transform -1 0 57696 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_76_572
timestamp 1621261055
transform 1 0 56064 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_576
timestamp 1621261055
transform 1 0 56448 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_579
timestamp 1621261055
transform 1 0 56736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_593
timestamp 1621261055
transform 1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_153
timestamp 1621261055
transform -1 0 58848 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_154
timestamp 1621261055
transform 1 0 1152 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_156
timestamp 1621261055
transform 1 0 1152 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_4
timestamp 1621261055
transform 1 0 1536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_12
timestamp 1621261055
transform 1 0 2304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_20
timestamp 1621261055
transform 1 0 3072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_4
timestamp 1621261055
transform 1 0 1536 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_12
timestamp 1621261055
transform 1 0 2304 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_20
timestamp 1621261055
transform 1 0 3072 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_29
timestamp 1621261055
transform 1 0 3936 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_28
timestamp 1621261055
transform 1 0 3840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_993
timestamp 1621261055
transform 1 0 3840 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_37
timestamp 1621261055
transform 1 0 4704 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_44
timestamp 1621261055
transform 1 0 5376 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_36
timestamp 1621261055
transform 1 0 4608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_53
timestamp 1621261055
transform 1 0 6240 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_45
timestamp 1621261055
transform 1 0 5472 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_52
timestamp 1621261055
transform 1 0 6144 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_77_54
timestamp 1621261055
transform 1 0 6336 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_983
timestamp 1621261055
transform 1 0 6432 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_56
timestamp 1621261055
transform 1 0 6528 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_64
timestamp 1621261055
transform 1 0 7296 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_72
timestamp 1621261055
transform 1 0 8064 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_80
timestamp 1621261055
transform 1 0 8832 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_61
timestamp 1621261055
transform 1 0 7008 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_69
timestamp 1621261055
transform 1 0 7776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_77
timestamp 1621261055
transform 1 0 8544 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_81
timestamp 1621261055
transform 1 0 8928 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_994
timestamp 1621261055
transform 1 0 9120 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_88
timestamp 1621261055
transform 1 0 9600 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_96
timestamp 1621261055
transform 1 0 10368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_104
timestamp 1621261055
transform 1 0 11136 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_108
timestamp 1621261055
transform 1 0 11520 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_84
timestamp 1621261055
transform 1 0 9216 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_92
timestamp 1621261055
transform 1 0 9984 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_100
timestamp 1621261055
transform 1 0 10752 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_108
timestamp 1621261055
transform 1 0 11520 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_114
timestamp 1621261055
transform 1 0 12096 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_110
timestamp 1621261055
transform 1 0 11712 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_111
timestamp 1621261055
transform 1 0 11808 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_984
timestamp 1621261055
transform 1 0 11712 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _215_
timestamp 1621261055
transform 1 0 11808 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_122
timestamp 1621261055
transform 1 0 12864 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_119
timestamp 1621261055
transform 1 0 12576 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_130
timestamp 1621261055
transform 1 0 13632 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_127
timestamp 1621261055
transform 1 0 13344 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_178
timestamp 1621261055
transform 1 0 13728 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _118_
timestamp 1621261055
transform 1 0 13920 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_995
timestamp 1621261055
transform 1 0 14400 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_136
timestamp 1621261055
transform 1 0 14208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_144
timestamp 1621261055
transform 1 0 14976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_152
timestamp 1621261055
transform 1 0 15744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_160
timestamp 1621261055
transform 1 0 16512 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_139
timestamp 1621261055
transform 1 0 14496 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_147
timestamp 1621261055
transform 1 0 15264 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_155
timestamp 1621261055
transform 1 0 16032 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_985
timestamp 1621261055
transform 1 0 16992 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_77_164
timestamp 1621261055
transform 1 0 16896 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_166
timestamp 1621261055
transform 1 0 17088 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_174
timestamp 1621261055
transform 1 0 17856 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_182
timestamp 1621261055
transform 1 0 18624 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_163
timestamp 1621261055
transform 1 0 16800 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_171
timestamp 1621261055
transform 1 0 17568 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_179
timestamp 1621261055
transform 1 0 18336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_187
timestamp 1621261055
transform 1 0 19104 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_996
timestamp 1621261055
transform 1 0 19680 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_190
timestamp 1621261055
transform 1 0 19392 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_198
timestamp 1621261055
transform 1 0 20160 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_206
timestamp 1621261055
transform 1 0 20928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_214
timestamp 1621261055
transform 1 0 21696 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_191
timestamp 1621261055
transform 1 0 19488 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_194
timestamp 1621261055
transform 1 0 19776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_202
timestamp 1621261055
transform 1 0 20544 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_210
timestamp 1621261055
transform 1 0 21312 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_986
timestamp 1621261055
transform 1 0 22272 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_218
timestamp 1621261055
transform 1 0 22080 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_221
timestamp 1621261055
transform 1 0 22368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_229
timestamp 1621261055
transform 1 0 23136 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_237
timestamp 1621261055
transform 1 0 23904 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_218
timestamp 1621261055
transform 1 0 22080 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_226
timestamp 1621261055
transform 1 0 22848 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_234
timestamp 1621261055
transform 1 0 23616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_242
timestamp 1621261055
transform 1 0 24384 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_78_249
timestamp 1621261055
transform 1 0 25056 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_246
timestamp 1621261055
transform 1 0 24768 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_245
timestamp 1621261055
transform 1 0 24672 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_997
timestamp 1621261055
transform 1 0 24960 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_78_255
timestamp 1621261055
transform 1 0 25632 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_253
timestamp 1621261055
transform 1 0 25440 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_253
timestamp 1621261055
transform 1 0 25440 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_161
timestamp 1621261055
transform 1 0 25728 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _099_
timestamp 1621261055
transform 1 0 25920 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_269
timestamp 1621261055
transform 1 0 26976 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_261
timestamp 1621261055
transform 1 0 26208 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_269
timestamp 1621261055
transform 1 0 26976 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_261
timestamp 1621261055
transform 1 0 26208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_987
timestamp 1621261055
transform 1 0 27552 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_273
timestamp 1621261055
transform 1 0 27360 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_276
timestamp 1621261055
transform 1 0 27648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_284
timestamp 1621261055
transform 1 0 28416 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_292
timestamp 1621261055
transform 1 0 29184 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_277
timestamp 1621261055
transform 1 0 27744 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_285
timestamp 1621261055
transform 1 0 28512 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_293
timestamp 1621261055
transform 1 0 29280 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_998
timestamp 1621261055
transform 1 0 30240 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_300
timestamp 1621261055
transform 1 0 29952 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_308
timestamp 1621261055
transform 1 0 30720 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_316
timestamp 1621261055
transform 1 0 31488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_324
timestamp 1621261055
transform 1 0 32256 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_301
timestamp 1621261055
transform 1 0 30048 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_304
timestamp 1621261055
transform 1 0 30336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_312
timestamp 1621261055
transform 1 0 31104 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_320
timestamp 1621261055
transform 1 0 31872 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_988
timestamp 1621261055
transform 1 0 32832 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_328
timestamp 1621261055
transform 1 0 32640 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_331
timestamp 1621261055
transform 1 0 32928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_339
timestamp 1621261055
transform 1 0 33696 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_347
timestamp 1621261055
transform 1 0 34464 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_328
timestamp 1621261055
transform 1 0 32640 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_336
timestamp 1621261055
transform 1 0 33408 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_344
timestamp 1621261055
transform 1 0 34176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_999
timestamp 1621261055
transform 1 0 35520 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_355
timestamp 1621261055
transform 1 0 35232 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_363
timestamp 1621261055
transform 1 0 36000 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_371
timestamp 1621261055
transform 1 0 36768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_352
timestamp 1621261055
transform 1 0 34944 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_356
timestamp 1621261055
transform 1 0 35328 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_359
timestamp 1621261055
transform 1 0 35616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_367
timestamp 1621261055
transform 1 0 36384 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_375
timestamp 1621261055
transform 1 0 37152 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_989
timestamp 1621261055
transform 1 0 38112 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_379
timestamp 1621261055
transform 1 0 37536 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_383
timestamp 1621261055
transform 1 0 37920 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_386
timestamp 1621261055
transform 1 0 38208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_394
timestamp 1621261055
transform 1 0 38976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_402
timestamp 1621261055
transform 1 0 39744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_383
timestamp 1621261055
transform 1 0 37920 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_391
timestamp 1621261055
transform 1 0 38688 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_399
timestamp 1621261055
transform 1 0 39456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1000
timestamp 1621261055
transform 1 0 40800 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_410
timestamp 1621261055
transform 1 0 40512 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_418
timestamp 1621261055
transform 1 0 41280 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_426
timestamp 1621261055
transform 1 0 42048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_407
timestamp 1621261055
transform 1 0 40224 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_411
timestamp 1621261055
transform 1 0 40608 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_414
timestamp 1621261055
transform 1 0 40896 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_422
timestamp 1621261055
transform 1 0 41664 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_430
timestamp 1621261055
transform 1 0 42432 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_438
timestamp 1621261055
transform 1 0 43200 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_438
timestamp 1621261055
transform 1 0 43200 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_434
timestamp 1621261055
transform 1 0 42816 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_990
timestamp 1621261055
transform 1 0 43392 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_446
timestamp 1621261055
transform 1 0 43968 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_449
timestamp 1621261055
transform 1 0 44256 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_441
timestamp 1621261055
transform 1 0 43488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_458
timestamp 1621261055
transform 1 0 45120 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_452
timestamp 1621261055
transform 1 0 44544 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_450
timestamp 1621261055
transform 1 0 44352 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_457
timestamp 1621261055
transform 1 0 45024 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_123
timestamp 1621261055
transform -1 0 44832 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _067_
timestamp 1621261055
transform -1 0 45120 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1001
timestamp 1621261055
transform 1 0 46080 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_465
timestamp 1621261055
transform 1 0 45792 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_473
timestamp 1621261055
transform 1 0 46560 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_481
timestamp 1621261055
transform 1 0 47328 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_466
timestamp 1621261055
transform 1 0 45888 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_469
timestamp 1621261055
transform 1 0 46176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_477
timestamp 1621261055
transform 1 0 46944 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_485
timestamp 1621261055
transform 1 0 47712 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_493
timestamp 1621261055
transform 1 0 48480 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_493
timestamp 1621261055
transform 1 0 48480 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_489
timestamp 1621261055
transform 1 0 48096 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_501
timestamp 1621261055
transform 1 0 49248 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_503
timestamp 1621261055
transform 1 0 49440 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_496
timestamp 1621261055
transform 1 0 48768 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_126
timestamp 1621261055
transform 1 0 48960 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_991
timestamp 1621261055
transform 1 0 48672 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _176_
timestamp 1621261055
transform 1 0 49152 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_509
timestamp 1621261055
transform 1 0 50016 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_511
timestamp 1621261055
transform 1 0 50208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1002
timestamp 1621261055
transform 1 0 51360 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_519
timestamp 1621261055
transform 1 0 50976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_527
timestamp 1621261055
transform 1 0 51744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_535
timestamp 1621261055
transform 1 0 52512 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_517
timestamp 1621261055
transform 1 0 50784 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_521
timestamp 1621261055
transform 1 0 51168 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_524
timestamp 1621261055
transform 1 0 51456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_532
timestamp 1621261055
transform 1 0 52224 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_540
timestamp 1621261055
transform 1 0 52992 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_548
timestamp 1621261055
transform 1 0 53760 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_549
timestamp 1621261055
transform 1 0 53856 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_547
timestamp 1621261055
transform 1 0 53664 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_543
timestamp 1621261055
transform 1 0 53280 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_556
timestamp 1621261055
transform 1 0 54528 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_551
timestamp 1621261055
transform 1 0 54048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_992
timestamp 1621261055
transform 1 0 53952 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_564
timestamp 1621261055
transform 1 0 55296 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_559
timestamp 1621261055
transform 1 0 54816 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_567
timestamp 1621261055
transform 1 0 55584 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_574
timestamp 1621261055
transform 1 0 56256 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_78_568
timestamp 1621261055
transform 1 0 55680 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_575
timestamp 1621261055
transform 1 0 56352 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_174
timestamp 1621261055
transform -1 0 55968 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _115_
timestamp 1621261055
transform -1 0 56256 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_579
timestamp 1621261055
transform 1 0 56736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_583
timestamp 1621261055
transform 1 0 57120 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1003
timestamp 1621261055
transform 1 0 56640 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_593
timestamp 1621261055
transform 1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_77_593
timestamp 1621261055
transform 1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_86
timestamp 1621261055
transform -1 0 57696 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_28
timestamp 1621261055
transform 1 0 57504 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output435
timestamp 1621261055
transform -1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output398
timestamp 1621261055
transform 1 0 57696 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_155
timestamp 1621261055
transform -1 0 58848 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_157
timestamp 1621261055
transform -1 0 58848 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_158
timestamp 1621261055
transform 1 0 1152 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output406
timestamp 1621261055
transform 1 0 1536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_36
timestamp 1621261055
transform 1 0 1920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_10
timestamp 1621261055
transform 1 0 2112 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_18
timestamp 1621261055
transform 1 0 2880 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_26
timestamp 1621261055
transform 1 0 3648 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output428
timestamp 1621261055
transform 1 0 4320 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_76
timestamp 1621261055
transform 1 0 4128 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_30
timestamp 1621261055
transform 1 0 4032 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_37
timestamp 1621261055
transform 1 0 4704 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_45
timestamp 1621261055
transform 1 0 5472 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_53
timestamp 1621261055
transform 1 0 6240 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1004
timestamp 1621261055
transform 1 0 6432 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output438
timestamp 1621261055
transform 1 0 7488 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_92
timestamp 1621261055
transform 1 0 7296 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_94
timestamp 1621261055
transform -1 0 9120 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_56
timestamp 1621261055
transform 1 0 6528 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_70
timestamp 1621261055
transform 1 0 7872 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_78
timestamp 1621261055
transform 1 0 8640 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_80
timestamp 1621261055
transform 1 0 8832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _183_
timestamp 1621261055
transform -1 0 10176 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output439
timestamp 1621261055
transform -1 0 9504 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_220
timestamp 1621261055
transform -1 0 9888 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_87
timestamp 1621261055
transform 1 0 9504 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_94
timestamp 1621261055
transform 1 0 10176 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_102
timestamp 1621261055
transform 1 0 10944 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _147_
timestamp 1621261055
transform 1 0 12576 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1005
timestamp 1621261055
transform 1 0 11712 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output442
timestamp 1621261055
transform 1 0 13824 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_207
timestamp 1621261055
transform 1 0 12384 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_111
timestamp 1621261055
transform 1 0 11808 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_115
timestamp 1621261055
transform 1 0 12192 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_122
timestamp 1621261055
transform 1 0 12864 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_130
timestamp 1621261055
transform 1 0 13632 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _010_
timestamp 1621261055
transform 1 0 14688 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _074_
timestamp 1621261055
transform 1 0 15360 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_139
timestamp 1621261055
transform 1 0 15168 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_136
timestamp 1621261055
transform 1 0 14208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_140
timestamp 1621261055
transform 1 0 14592 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_144
timestamp 1621261055
transform 1 0 14976 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_151
timestamp 1621261055
transform 1 0 15648 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_159
timestamp 1621261055
transform 1 0 16416 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1006
timestamp 1621261055
transform 1 0 16992 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_163
timestamp 1621261055
transform 1 0 16800 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_166
timestamp 1621261055
transform 1 0 17088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_174
timestamp 1621261055
transform 1 0 17856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_182
timestamp 1621261055
transform 1 0 18624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output409
timestamp 1621261055
transform 1 0 20160 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_190
timestamp 1621261055
transform 1 0 19392 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_202
timestamp 1621261055
transform 1 0 20544 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_210
timestamp 1621261055
transform 1 0 21312 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1007
timestamp 1621261055
transform 1 0 22272 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output411
timestamp 1621261055
transform -1 0 23712 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_40
timestamp 1621261055
transform -1 0 23328 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_218
timestamp 1621261055
transform 1 0 22080 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_221
timestamp 1621261055
transform 1 0 22368 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_235
timestamp 1621261055
transform 1 0 23712 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_243
timestamp 1621261055
transform 1 0 24480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _199_
timestamp 1621261055
transform -1 0 25920 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output412
timestamp 1621261055
transform -1 0 25248 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_42
timestamp 1621261055
transform -1 0 24864 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_229
timestamp 1621261055
transform -1 0 25632 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_251
timestamp 1621261055
transform 1 0 25248 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_258
timestamp 1621261055
transform 1 0 25920 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_266
timestamp 1621261055
transform 1 0 26688 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _161_
timestamp 1621261055
transform 1 0 28896 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1008
timestamp 1621261055
transform 1 0 27552 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_79_274
timestamp 1621261055
transform 1 0 27456 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_276
timestamp 1621261055
transform 1 0 27648 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_284
timestamp 1621261055
transform 1 0 28416 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_288
timestamp 1621261055
transform 1 0 28800 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_292
timestamp 1621261055
transform 1 0 29184 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_300
timestamp 1621261055
transform 1 0 29952 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_308
timestamp 1621261055
transform 1 0 30720 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_316
timestamp 1621261055
transform 1 0 31488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_324
timestamp 1621261055
transform 1 0 32256 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1009
timestamp 1621261055
transform 1 0 32832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_328
timestamp 1621261055
transform 1 0 32640 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_331
timestamp 1621261055
transform 1 0 32928 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_339
timestamp 1621261055
transform 1 0 33696 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_347
timestamp 1621261055
transform 1 0 34464 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_355
timestamp 1621261055
transform 1 0 35232 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_363
timestamp 1621261055
transform 1 0 36000 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_371
timestamp 1621261055
transform 1 0 36768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1010
timestamp 1621261055
transform 1 0 38112 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output422
timestamp 1621261055
transform -1 0 39456 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_62
timestamp 1621261055
transform -1 0 39072 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_379
timestamp 1621261055
transform 1 0 37536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_383
timestamp 1621261055
transform 1 0 37920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_386
timestamp 1621261055
transform 1 0 38208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_390
timestamp 1621261055
transform 1 0 38592 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_392
timestamp 1621261055
transform 1 0 38784 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_399
timestamp 1621261055
transform 1 0 39456 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_79_409
timestamp 1621261055
transform 1 0 40416 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_407
timestamp 1621261055
transform 1 0 40224 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_64
timestamp 1621261055
transform -1 0 40704 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output423
timestamp 1621261055
transform -1 0 41088 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_418
timestamp 1621261055
transform 1 0 41280 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_65
timestamp 1621261055
transform -1 0 41280 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_426
timestamp 1621261055
transform 1 0 42048 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_216
timestamp 1621261055
transform 1 0 42144 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _152_
timestamp 1621261055
transform 1 0 42336 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_79_432
timestamp 1621261055
transform 1 0 42624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1011
timestamp 1621261055
transform 1 0 43392 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_71
timestamp 1621261055
transform -1 0 45408 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_441
timestamp 1621261055
transform 1 0 43488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_449
timestamp 1621261055
transform 1 0 44256 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_457
timestamp 1621261055
transform 1 0 45024 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output426
timestamp 1621261055
transform -1 0 45792 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output427
timestamp 1621261055
transform -1 0 47328 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_73
timestamp 1621261055
transform -1 0 46944 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_74
timestamp 1621261055
transform -1 0 47520 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_465
timestamp 1621261055
transform 1 0 45792 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_473
timestamp 1621261055
transform 1 0 46560 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_483
timestamp 1621261055
transform 1 0 47520 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _020_
timestamp 1621261055
transform 1 0 48000 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1012
timestamp 1621261055
transform 1 0 48672 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_79_487
timestamp 1621261055
transform 1 0 47904 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_79_491
timestamp 1621261055
transform 1 0 48288 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_496
timestamp 1621261055
transform 1 0 48768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_504
timestamp 1621261055
transform 1 0 49536 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_512
timestamp 1621261055
transform 1 0 50304 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output431
timestamp 1621261055
transform -1 0 52128 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_80
timestamp 1621261055
transform -1 0 51744 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_520
timestamp 1621261055
transform 1 0 51072 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_524
timestamp 1621261055
transform 1 0 51456 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_531
timestamp 1621261055
transform 1 0 52128 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_539
timestamp 1621261055
transform 1 0 52896 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1013
timestamp 1621261055
transform 1 0 53952 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_135
timestamp 1621261055
transform -1 0 55776 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_547
timestamp 1621261055
transform 1 0 53664 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_549
timestamp 1621261055
transform 1 0 53856 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_551
timestamp 1621261055
transform 1 0 54048 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_559
timestamp 1621261055
transform 1 0 54816 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _070_
timestamp 1621261055
transform -1 0 56064 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output397
timestamp 1621261055
transform -1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output434
timestamp 1621261055
transform -1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_26
timestamp 1621261055
transform -1 0 57504 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_85
timestamp 1621261055
transform -1 0 56448 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_572
timestamp 1621261055
transform 1 0 56064 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_580
timestamp 1621261055
transform 1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_584
timestamp 1621261055
transform 1 0 57216 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_79_591
timestamp 1621261055
transform 1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_159
timestamp 1621261055
transform -1 0 58848 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_595
timestamp 1621261055
transform 1 0 58272 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_160
timestamp 1621261055
transform 1 0 1152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output368
timestamp 1621261055
transform 1 0 1536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output379
timestamp 1621261055
transform 1 0 2304 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output417
timestamp 1621261055
transform 1 0 3072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_52
timestamp 1621261055
transform 1 0 2880 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_8
timestamp 1621261055
transform 1 0 1920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_16
timestamp 1621261055
transform 1 0 2688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_24
timestamp 1621261055
transform 1 0 3456 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_29
timestamp 1621261055
transform 1 0 3936 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1014
timestamp 1621261055
transform 1 0 3840 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output390
timestamp 1621261055
transform 1 0 4320 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_41
timestamp 1621261055
transform 1 0 5088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_37
timestamp 1621261055
transform 1 0 4704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_43
timestamp 1621261055
transform 1 0 5280 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output399
timestamp 1621261055
transform 1 0 5376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_48
timestamp 1621261055
transform 1 0 5760 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_90
timestamp 1621261055
transform 1 0 5952 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output437
timestamp 1621261055
transform 1 0 6144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output400
timestamp 1621261055
transform 1 0 7008 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output401
timestamp 1621261055
transform -1 0 8736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_30
timestamp 1621261055
transform -1 0 8352 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_56
timestamp 1621261055
transform 1 0 6528 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_60
timestamp 1621261055
transform 1 0 6912 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_65
timestamp 1621261055
transform 1 0 7392 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_79
timestamp 1621261055
transform 1 0 8736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1015
timestamp 1621261055
transform 1 0 9120 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output402
timestamp 1621261055
transform 1 0 10176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output440
timestamp 1621261055
transform 1 0 10944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_32
timestamp 1621261055
transform 1 0 9984 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_84
timestamp 1621261055
transform 1 0 9216 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_98
timestamp 1621261055
transform 1 0 10560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_106
timestamp 1621261055
transform 1 0 11328 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output403
timestamp 1621261055
transform 1 0 11712 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output404
timestamp 1621261055
transform -1 0 13728 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output441
timestamp 1621261055
transform 1 0 12480 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_34
timestamp 1621261055
transform -1 0 13344 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_114
timestamp 1621261055
transform 1 0 12096 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_122
timestamp 1621261055
transform 1 0 12864 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_124
timestamp 1621261055
transform 1 0 13056 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_131
timestamp 1621261055
transform 1 0 13728 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_135
timestamp 1621261055
transform 1 0 14112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1016
timestamp 1621261055
transform 1 0 14400 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output405
timestamp 1621261055
transform 1 0 14880 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output443
timestamp 1621261055
transform -1 0 16032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_96
timestamp 1621261055
transform -1 0 15648 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_137
timestamp 1621261055
transform 1 0 14304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_139
timestamp 1621261055
transform 1 0 14496 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_147
timestamp 1621261055
transform 1 0 15264 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_155
timestamp 1621261055
transform 1 0 16032 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output370
timestamp 1621261055
transform 1 0 18048 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output407
timestamp 1621261055
transform 1 0 16992 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output408
timestamp 1621261055
transform 1 0 18816 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_163
timestamp 1621261055
transform 1 0 16800 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_169
timestamp 1621261055
transform 1 0 17376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_173
timestamp 1621261055
transform 1 0 17760 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_175
timestamp 1621261055
transform 1 0 17952 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_180
timestamp 1621261055
transform 1 0 18432 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_188
timestamp 1621261055
transform 1 0 19200 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_192
timestamp 1621261055
transform 1 0 19584 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1017
timestamp 1621261055
transform 1 0 19680 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_194
timestamp 1621261055
transform 1 0 19776 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output371
timestamp 1621261055
transform 1 0 20160 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_202
timestamp 1621261055
transform 1 0 20544 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_206
timestamp 1621261055
transform 1 0 20928 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_3
timestamp 1621261055
transform 1 0 21024 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_213
timestamp 1621261055
transform 1 0 21600 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output372
timestamp 1621261055
transform 1 0 21216 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_38
timestamp 1621261055
transform 1 0 21792 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output373
timestamp 1621261055
transform 1 0 22752 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output374
timestamp 1621261055
transform 1 0 24192 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output410
timestamp 1621261055
transform 1 0 21984 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_221
timestamp 1621261055
transform 1 0 22368 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_229
timestamp 1621261055
transform 1 0 23136 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_237
timestamp 1621261055
transform 1 0 23904 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_239
timestamp 1621261055
transform 1 0 24096 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1018
timestamp 1621261055
transform 1 0 24960 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output375
timestamp 1621261055
transform 1 0 25920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output413
timestamp 1621261055
transform -1 0 27072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_44
timestamp 1621261055
transform -1 0 26688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_244
timestamp 1621261055
transform 1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_249
timestamp 1621261055
transform 1 0 25056 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_80_257
timestamp 1621261055
transform 1 0 25824 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_262
timestamp 1621261055
transform 1 0 26304 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_270
timestamp 1621261055
transform 1 0 27072 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_272
timestamp 1621261055
transform 1 0 27264 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_5
timestamp 1621261055
transform -1 0 27552 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_279
timestamp 1621261055
transform 1 0 27936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output376
timestamp 1621261055
transform -1 0 27936 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_46
timestamp 1621261055
transform -1 0 28320 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output414
timestamp 1621261055
transform -1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_287
timestamp 1621261055
transform 1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_291
timestamp 1621261055
transform 1 0 29088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_48
timestamp 1621261055
transform -1 0 29472 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output415
timestamp 1621261055
transform -1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1019
timestamp 1621261055
transform 1 0 30240 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output378
timestamp 1621261055
transform 1 0 30720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output380
timestamp 1621261055
transform 1 0 32256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output416
timestamp 1621261055
transform 1 0 31488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_50
timestamp 1621261055
transform 1 0 31296 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_299
timestamp 1621261055
transform 1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_304
timestamp 1621261055
transform 1 0 30336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_312
timestamp 1621261055
transform 1 0 31104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_320
timestamp 1621261055
transform 1 0 31872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output381
timestamp 1621261055
transform 1 0 33792 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output418
timestamp 1621261055
transform -1 0 33408 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output419
timestamp 1621261055
transform -1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_7
timestamp 1621261055
transform 1 0 33600 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_54
timestamp 1621261055
transform -1 0 33024 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_56
timestamp 1621261055
transform -1 0 34560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_328
timestamp 1621261055
transform 1 0 32640 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_336
timestamp 1621261055
transform 1 0 33408 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_344
timestamp 1621261055
transform 1 0 34176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_352
timestamp 1621261055
transform 1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_359
timestamp 1621261055
transform 1 0 35616 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_356
timestamp 1621261055
transform 1 0 35328 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1020
timestamp 1621261055
transform 1 0 35520 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_9
timestamp 1621261055
transform -1 0 36000 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output382
timestamp 1621261055
transform -1 0 36384 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_367
timestamp 1621261055
transform 1 0 36384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_58
timestamp 1621261055
transform -1 0 36768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_375
timestamp 1621261055
transform 1 0 37152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output420
timestamp 1621261055
transform -1 0 37152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_60
timestamp 1621261055
transform 1 0 37344 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output384
timestamp 1621261055
transform -1 0 38976 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output385
timestamp 1621261055
transform 1 0 40032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output421
timestamp 1621261055
transform 1 0 37536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_13
timestamp 1621261055
transform -1 0 38592 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_15
timestamp 1621261055
transform 1 0 39840 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_383
timestamp 1621261055
transform 1 0 37920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_387
timestamp 1621261055
transform 1 0 38304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_394
timestamp 1621261055
transform 1 0 38976 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_80_402
timestamp 1621261055
transform 1 0 39744 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1021
timestamp 1621261055
transform 1 0 40800 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output386
timestamp 1621261055
transform 1 0 41760 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output424
timestamp 1621261055
transform -1 0 42912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_67
timestamp 1621261055
transform -1 0 42528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_409
timestamp 1621261055
transform 1 0 40416 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_414
timestamp 1621261055
transform 1 0 40896 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_80_422
timestamp 1621261055
transform 1 0 41664 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_427
timestamp 1621261055
transform 1 0 42144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_435
timestamp 1621261055
transform 1 0 42912 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_17
timestamp 1621261055
transform -1 0 43296 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output387
timestamp 1621261055
transform -1 0 43680 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_443
timestamp 1621261055
transform 1 0 43680 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_69
timestamp 1621261055
transform -1 0 44064 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_451
timestamp 1621261055
transform 1 0 44448 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output425
timestamp 1621261055
transform -1 0 44448 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_453
timestamp 1621261055
transform 1 0 44640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_19
timestamp 1621261055
transform -1 0 44928 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output388
timestamp 1621261055
transform -1 0 45312 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1022
timestamp 1621261055
transform 1 0 46080 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output389
timestamp 1621261055
transform 1 0 46560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_460
timestamp 1621261055
transform 1 0 45312 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_469
timestamp 1621261055
transform 1 0 46176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_477
timestamp 1621261055
transform 1 0 46944 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_485
timestamp 1621261055
transform 1 0 47712 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_80_487
timestamp 1621261055
transform 1 0 47904 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output391
timestamp 1621261055
transform 1 0 48000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_492
timestamp 1621261055
transform 1 0 48384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_78
timestamp 1621261055
transform -1 0 48768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_500
timestamp 1621261055
transform 1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output429
timestamp 1621261055
transform -1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_504
timestamp 1621261055
transform 1 0 49536 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output392
timestamp 1621261055
transform 1 0 49632 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_509
timestamp 1621261055
transform 1 0 50016 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output430
timestamp 1621261055
transform 1 0 50400 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1023
timestamp 1621261055
transform 1 0 51360 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output393
timestamp 1621261055
transform -1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output394
timestamp 1621261055
transform -1 0 53184 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_21
timestamp 1621261055
transform -1 0 51840 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_23
timestamp 1621261055
transform -1 0 52800 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_517
timestamp 1621261055
transform 1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_521
timestamp 1621261055
transform 1 0 51168 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_524
timestamp 1621261055
transform 1 0 51456 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_532
timestamp 1621261055
transform 1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output395
timestamp 1621261055
transform 1 0 54336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output432
timestamp 1621261055
transform -1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output433
timestamp 1621261055
transform -1 0 55488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_81
timestamp 1621261055
transform -1 0 53568 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_83
timestamp 1621261055
transform -1 0 55104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_84
timestamp 1621261055
transform -1 0 55680 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_542
timestamp 1621261055
transform 1 0 53184 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_550
timestamp 1621261055
transform 1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_558
timestamp 1621261055
transform 1 0 54720 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1024
timestamp 1621261055
transform 1 0 56640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input31
timestamp 1621261055
transform 1 0 57696 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output396
timestamp 1621261055
transform -1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_25
timestamp 1621261055
transform -1 0 55872 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_574
timestamp 1621261055
transform 1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_579
timestamp 1621261055
transform 1 0 56736 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_587
timestamp 1621261055
transform 1 0 57504 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_593
timestamp 1621261055
transform 1 0 58080 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_161
timestamp 1621261055
transform -1 0 58848 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_162
timestamp 1621261055
transform 1 0 1152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input12
timestamp 1621261055
transform 1 0 2400 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_9
timestamp 1621261055
transform 1 0 2016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_18
timestamp 1621261055
transform 1 0 2880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_26
timestamp 1621261055
transform 1 0 3648 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1025
timestamp 1621261055
transform 1 0 3840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input23
timestamp 1621261055
transform 1 0 5760 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input32
timestamp 1621261055
transform 1 0 4896 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_8  FILLER_81_29
timestamp 1621261055
transform 1 0 3936 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_37
timestamp 1621261055
transform 1 0 4704 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_44
timestamp 1621261055
transform 1 0 5376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_52
timestamp 1621261055
transform 1 0 6144 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1026
timestamp 1621261055
transform 1 0 6528 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input33
timestamp 1621261055
transform 1 0 7008 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input34
timestamp 1621261055
transform 1 0 8064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_57
timestamp 1621261055
transform 1 0 6624 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_66
timestamp 1621261055
transform 1 0 7488 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_70
timestamp 1621261055
transform 1 0 7872 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_76
timestamp 1621261055
transform 1 0 8448 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1027
timestamp 1621261055
transform 1 0 9216 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  input35
timestamp 1621261055
transform 1 0 9696 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input36
timestamp 1621261055
transform 1 0 11040 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_85
timestamp 1621261055
transform 1 0 9312 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_93
timestamp 1621261055
transform 1 0 10080 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_101
timestamp 1621261055
transform 1 0 10848 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_108
timestamp 1621261055
transform 1 0 11520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1028
timestamp 1621261055
transform 1 0 11904 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input37
timestamp 1621261055
transform 1 0 12768 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_2  output369
timestamp 1621261055
transform -1 0 14208 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_1
timestamp 1621261055
transform -1 0 13824 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_113
timestamp 1621261055
transform 1 0 12000 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_126
timestamp 1621261055
transform 1 0 13248 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1029
timestamp 1621261055
transform 1 0 14592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input2
timestamp 1621261055
transform 1 0 15936 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input38
timestamp 1621261055
transform 1 0 15072 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_136
timestamp 1621261055
transform 1 0 14208 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_141
timestamp 1621261055
transform 1 0 14688 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_149
timestamp 1621261055
transform 1 0 15456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_153
timestamp 1621261055
transform 1 0 15840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_159
timestamp 1621261055
transform 1 0 16416 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1030
timestamp 1621261055
transform 1 0 17280 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input3
timestamp 1621261055
transform 1 0 17760 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input4
timestamp 1621261055
transform 1 0 19104 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_1  FILLER_81_167
timestamp 1621261055
transform 1 0 17184 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_169
timestamp 1621261055
transform 1 0 17376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_178
timestamp 1621261055
transform 1 0 18240 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_186
timestamp 1621261055
transform 1 0 19008 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1031
timestamp 1621261055
transform 1 0 19968 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input5
timestamp 1621261055
transform 1 0 20640 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input6
timestamp 1621261055
transform 1 0 21888 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_192
timestamp 1621261055
transform 1 0 19584 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_197
timestamp 1621261055
transform 1 0 20064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_201
timestamp 1621261055
transform 1 0 20448 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_208
timestamp 1621261055
transform 1 0 21120 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1032
timestamp 1621261055
transform 1 0 22656 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input7
timestamp 1621261055
transform 1 0 23808 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_220
timestamp 1621261055
transform 1 0 22272 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_225
timestamp 1621261055
transform 1 0 22752 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_233
timestamp 1621261055
transform 1 0 23520 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_235
timestamp 1621261055
transform 1 0 23712 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_241
timestamp 1621261055
transform 1 0 24288 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1033
timestamp 1621261055
transform 1 0 25344 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input8
timestamp 1621261055
transform 1 0 25824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input9
timestamp 1621261055
transform 1 0 26976 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_249
timestamp 1621261055
transform 1 0 25056 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_251
timestamp 1621261055
transform 1 0 25248 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_253
timestamp 1621261055
transform 1 0 25440 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_261
timestamp 1621261055
transform 1 0 26208 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1034
timestamp 1621261055
transform 1 0 28032 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input10
timestamp 1621261055
transform 1 0 28608 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_274
timestamp 1621261055
transform 1 0 27456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_278
timestamp 1621261055
transform 1 0 27840 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_281
timestamp 1621261055
transform 1 0 28128 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_285
timestamp 1621261055
transform 1 0 28512 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_290
timestamp 1621261055
transform 1 0 28992 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1035
timestamp 1621261055
transform 1 0 30720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input11
timestamp 1621261055
transform 1 0 29856 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input13
timestamp 1621261055
transform 1 0 31680 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_298
timestamp 1621261055
transform 1 0 29760 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_304
timestamp 1621261055
transform 1 0 30336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_309
timestamp 1621261055
transform 1 0 30816 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_317
timestamp 1621261055
transform 1 0 31584 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_322
timestamp 1621261055
transform 1 0 32064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1036
timestamp 1621261055
transform 1 0 33408 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input14
timestamp 1621261055
transform 1 0 33888 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input15
timestamp 1621261055
transform 1 0 34848 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output377
timestamp 1621261055
transform 1 0 32448 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_330
timestamp 1621261055
transform 1 0 32832 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_334
timestamp 1621261055
transform 1 0 33216 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_337
timestamp 1621261055
transform 1 0 33504 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_346
timestamp 1621261055
transform 1 0 34368 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_350
timestamp 1621261055
transform 1 0 34752 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1037
timestamp 1621261055
transform 1 0 36096 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input16 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 36576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_8  FILLER_81_355
timestamp 1621261055
transform 1 0 35232 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_363
timestamp 1621261055
transform 1 0 36000 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_365
timestamp 1621261055
transform 1 0 36192 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_375
timestamp 1621261055
transform 1 0 37152 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1038
timestamp 1621261055
transform 1 0 38784 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input17
timestamp 1621261055
transform 1 0 38016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_4  input18
timestamp 1621261055
transform 1 0 39648 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_1  FILLER_81_383
timestamp 1621261055
transform 1 0 37920 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_388
timestamp 1621261055
transform 1 0 38400 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_393
timestamp 1621261055
transform 1 0 38880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1039
timestamp 1621261055
transform 1 0 41472 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input19
timestamp 1621261055
transform 1 0 41952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output383
timestamp 1621261055
transform -1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_11
timestamp 1621261055
transform -1 0 40608 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_407
timestamp 1621261055
transform 1 0 40224 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_415
timestamp 1621261055
transform 1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_419
timestamp 1621261055
transform 1 0 41376 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_421
timestamp 1621261055
transform 1 0 41568 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_429
timestamp 1621261055
transform 1 0 42336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1040
timestamp 1621261055
transform 1 0 44160 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input20
timestamp 1621261055
transform 1 0 42816 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input21
timestamp 1621261055
transform 1 0 44640 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_433
timestamp 1621261055
transform 1 0 42720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_440
timestamp 1621261055
transform 1 0 43392 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_449
timestamp 1621261055
transform 1 0 44256 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_457
timestamp 1621261055
transform 1 0 45024 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1041
timestamp 1621261055
transform 1 0 46848 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input22
timestamp 1621261055
transform 1 0 45888 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input24
timestamp 1621261055
transform 1 0 47520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_465
timestamp 1621261055
transform 1 0 45792 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_472
timestamp 1621261055
transform 1 0 46464 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_477
timestamp 1621261055
transform 1 0 46944 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_481
timestamp 1621261055
transform 1 0 47328 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1042
timestamp 1621261055
transform 1 0 49536 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input25
timestamp 1621261055
transform 1 0 48576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_487
timestamp 1621261055
transform 1 0 47904 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_491
timestamp 1621261055
transform 1 0 48288 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_493
timestamp 1621261055
transform 1 0 48480 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_500
timestamp 1621261055
transform 1 0 49152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_505
timestamp 1621261055
transform 1 0 49632 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_513
timestamp 1621261055
transform 1 0 50400 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1043
timestamp 1621261055
transform 1 0 52224 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input26
timestamp 1621261055
transform 1 0 50688 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_4  input27
timestamp 1621261055
transform 1 0 52704 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_1  FILLER_81_515
timestamp 1621261055
transform 1 0 50592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_522
timestamp 1621261055
transform 1 0 51264 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_530
timestamp 1621261055
transform 1 0 52032 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_533
timestamp 1621261055
transform 1 0 52320 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1044
timestamp 1621261055
transform 1 0 54912 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input28
timestamp 1621261055
transform 1 0 53856 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_4  input29
timestamp 1621261055
transform 1 0 55392 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_543
timestamp 1621261055
transform 1 0 53280 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_547
timestamp 1621261055
transform 1 0 53664 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_553
timestamp 1621261055
transform 1 0 54240 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_557
timestamp 1621261055
transform 1 0 54624 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_559
timestamp 1621261055
transform 1 0 54816 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_561
timestamp 1621261055
transform 1 0 55008 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1045
timestamp 1621261055
transform 1 0 57600 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input30
timestamp 1621261055
transform 1 0 56640 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_571
timestamp 1621261055
transform 1 0 55968 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_575
timestamp 1621261055
transform 1 0 56352 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_577
timestamp 1621261055
transform 1 0 56544 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_584
timestamp 1621261055
transform 1 0 57216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_589
timestamp 1621261055
transform 1 0 57696 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_163
timestamp 1621261055
transform -1 0 58848 0 1 56610
box -38 -49 422 715
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 114 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 115 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 116 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 117 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 118 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 119 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 120 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 121 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 122 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 123 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 124 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 125 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 126 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 127 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 128 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 129 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 130 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 131 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 132 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 133 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 134 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 135 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 136 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 137 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 138 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 139 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 140 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 141 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 142 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 143 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 144 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 145 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 146 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 147 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 148 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 149 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 150 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 151 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 152 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 153 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 154 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 155 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 156 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 157 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 158 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 159 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 160 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 161 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 162 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 163 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 164 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 165 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 166 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 167 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 168 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 169 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 170 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 171 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 172 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 173 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 174 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 175 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 176 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 177 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 178 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 179 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 180 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 181 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 182 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 183 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 184 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 185 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 186 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 187 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 188 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 189 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 190 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 191 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 192 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 193 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 194 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 195 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 196 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 197 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 198 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 199 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 200 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 201 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 202 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 203 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 204 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 205 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 206 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 207 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 208 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 209 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 210 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 211 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 212 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 213 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 214 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 215 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 216 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 217 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 218 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 219 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 220 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 221 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 222 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 223 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 224 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 225 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 226 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 227 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 228 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 229 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 230 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 231 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 232 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 233 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 234 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 235 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 236 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 237 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 238 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 239 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 240 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 241 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 242 nsew signal tristate
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 243 nsew signal tristate
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 244 nsew signal tristate
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 245 nsew signal tristate
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 246 nsew signal tristate
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 247 nsew signal tristate
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 248 nsew signal tristate
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 249 nsew signal tristate
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 250 nsew signal tristate
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 251 nsew signal tristate
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 252 nsew signal tristate
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 253 nsew signal tristate
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 254 nsew signal tristate
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 255 nsew signal tristate
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 256 nsew signal tristate
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 257 nsew signal tristate
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 258 nsew signal tristate
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 259 nsew signal tristate
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 260 nsew signal tristate
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 261 nsew signal tristate
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 262 nsew signal tristate
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 263 nsew signal tristate
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 264 nsew signal tristate
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 265 nsew signal tristate
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 266 nsew signal tristate
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 267 nsew signal tristate
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 268 nsew signal tristate
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 269 nsew signal tristate
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 270 nsew signal tristate
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 271 nsew signal tristate
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 272 nsew signal tristate
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 273 nsew signal tristate
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 274 nsew signal tristate
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 275 nsew signal tristate
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 276 nsew signal tristate
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 277 nsew signal tristate
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 278 nsew signal tristate
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 279 nsew signal tristate
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 280 nsew signal tristate
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 281 nsew signal tristate
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 282 nsew signal tristate
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 283 nsew signal tristate
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 284 nsew signal tristate
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 285 nsew signal tristate
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 286 nsew signal tristate
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 287 nsew signal tristate
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 288 nsew signal tristate
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 289 nsew signal tristate
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 290 nsew signal tristate
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 291 nsew signal tristate
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 292 nsew signal tristate
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 293 nsew signal tristate
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 294 nsew signal tristate
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 295 nsew signal tristate
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 296 nsew signal tristate
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 297 nsew signal tristate
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 298 nsew signal tristate
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 299 nsew signal tristate
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 300 nsew signal tristate
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 301 nsew signal tristate
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 302 nsew signal tristate
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 303 nsew signal tristate
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 304 nsew signal tristate
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 305 nsew signal tristate
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 306 nsew signal tristate
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 307 nsew signal tristate
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 308 nsew signal tristate
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 309 nsew signal tristate
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 310 nsew signal tristate
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 311 nsew signal tristate
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 312 nsew signal tristate
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 313 nsew signal tristate
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 314 nsew signal tristate
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 315 nsew signal tristate
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 316 nsew signal tristate
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 317 nsew signal tristate
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 318 nsew signal tristate
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 319 nsew signal tristate
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 320 nsew signal tristate
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 321 nsew signal tristate
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 322 nsew signal tristate
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 323 nsew signal tristate
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 324 nsew signal tristate
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 325 nsew signal tristate
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 326 nsew signal tristate
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 327 nsew signal tristate
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 328 nsew signal tristate
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 329 nsew signal tristate
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 330 nsew signal tristate
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 331 nsew signal tristate
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 332 nsew signal tristate
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 333 nsew signal tristate
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 334 nsew signal tristate
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 335 nsew signal tristate
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 336 nsew signal tristate
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 337 nsew signal tristate
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 338 nsew signal tristate
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 339 nsew signal tristate
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 340 nsew signal tristate
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 341 nsew signal tristate
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 342 nsew signal tristate
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 343 nsew signal tristate
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 344 nsew signal tristate
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 345 nsew signal tristate
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 346 nsew signal tristate
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 347 nsew signal tristate
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 348 nsew signal tristate
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 349 nsew signal tristate
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 350 nsew signal tristate
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 351 nsew signal tristate
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 352 nsew signal tristate
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 353 nsew signal tristate
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 354 nsew signal tristate
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 355 nsew signal tristate
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 356 nsew signal tristate
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 357 nsew signal tristate
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 358 nsew signal tristate
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 359 nsew signal tristate
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 360 nsew signal tristate
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 361 nsew signal tristate
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 362 nsew signal tristate
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 363 nsew signal tristate
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 364 nsew signal tristate
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 365 nsew signal tristate
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 366 nsew signal tristate
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 367 nsew signal tristate
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 368 nsew signal tristate
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 369 nsew signal tristate
rlabel metal2 s 13172 0 13228 800 6 la_oen[0]
port 370 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oen[100]
port 371 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oen[101]
port 372 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oen[102]
port 373 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oen[103]
port 374 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oen[104]
port 375 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oen[105]
port 376 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oen[106]
port 377 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oen[107]
port 378 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oen[108]
port 379 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oen[109]
port 380 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oen[10]
port 381 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oen[110]
port 382 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oen[111]
port 383 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oen[112]
port 384 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oen[113]
port 385 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oen[114]
port 386 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oen[115]
port 387 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oen[116]
port 388 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oen[117]
port 389 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oen[118]
port 390 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oen[119]
port 391 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oen[120]
port 393 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oen[121]
port 394 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oen[122]
port 395 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oen[123]
port 396 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oen[124]
port 397 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oen[125]
port 398 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oen[126]
port 399 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oen[127]
port 400 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oen[12]
port 401 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oen[13]
port 402 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oen[14]
port 403 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oen[15]
port 404 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oen[16]
port 405 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oen[18]
port 407 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oen[19]
port 408 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oen[1]
port 409 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oen[20]
port 410 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oen[21]
port 411 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oen[22]
port 412 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oen[24]
port 414 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oen[25]
port 415 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oen[26]
port 416 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oen[27]
port 417 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oen[28]
port 418 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oen[2]
port 420 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oen[30]
port 421 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oen[31]
port 422 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oen[32]
port 423 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oen[33]
port 424 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oen[34]
port 425 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oen[36]
port 427 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oen[37]
port 428 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oen[38]
port 429 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oen[39]
port 430 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oen[3]
port 431 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oen[40]
port 432 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oen[42]
port 434 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oen[43]
port 435 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oen[44]
port 436 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oen[45]
port 437 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oen[46]
port 438 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oen[48]
port 440 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oen[49]
port 441 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oen[4]
port 442 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oen[50]
port 443 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oen[51]
port 444 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oen[52]
port 445 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oen[54]
port 447 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oen[55]
port 448 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oen[56]
port 449 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oen[57]
port 450 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oen[58]
port 451 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oen[60]
port 454 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oen[61]
port 455 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oen[62]
port 456 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oen[63]
port 457 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oen[64]
port 458 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oen[66]
port 460 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oen[67]
port 461 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oen[68]
port 462 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oen[69]
port 463 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oen[6]
port 464 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oen[70]
port 465 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oen[72]
port 467 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oen[73]
port 468 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oen[74]
port 469 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oen[75]
port 470 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oen[76]
port 471 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oen[78]
port 473 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oen[79]
port 474 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oen[7]
port 475 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oen[80]
port 476 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oen[81]
port 477 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oen[82]
port 478 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oen[84]
port 480 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oen[85]
port 481 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oen[86]
port 482 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oen[87]
port 483 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oen[88]
port 484 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oen[89]
port 485 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oen[8]
port 486 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oen[90]
port 487 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oen[91]
port 488 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oen[92]
port 489 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oen[93]
port 490 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oen[94]
port 491 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oen[95]
port 492 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oen[96]
port 493 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oen[97]
port 494 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oen[98]
port 495 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oen[99]
port 496 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oen[9]
port 497 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 498 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 499 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 500 nsew signal tristate
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 501 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 502 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 503 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 504 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 505 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 506 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 507 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 508 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 509 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 510 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 511 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 512 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 513 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 514 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 515 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 516 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 517 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 518 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 519 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 520 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 521 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 522 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 523 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 524 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 525 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 526 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 527 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 528 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 529 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 530 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 531 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 532 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 533 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 534 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 535 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 536 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 537 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 538 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 539 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 540 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 541 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 542 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 543 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 544 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 545 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 546 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 547 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 548 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 549 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 550 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 551 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 552 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 553 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 554 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 555 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 556 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 557 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 558 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 559 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 560 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 561 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 562 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 563 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 564 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 565 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 566 nsew signal tristate
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 567 nsew signal tristate
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 568 nsew signal tristate
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 569 nsew signal tristate
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 570 nsew signal tristate
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 571 nsew signal tristate
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 572 nsew signal tristate
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 573 nsew signal tristate
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 574 nsew signal tristate
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 575 nsew signal tristate
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 576 nsew signal tristate
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 577 nsew signal tristate
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 578 nsew signal tristate
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 579 nsew signal tristate
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 580 nsew signal tristate
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 581 nsew signal tristate
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 582 nsew signal tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew signal tristate
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 584 nsew signal tristate
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 585 nsew signal tristate
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 586 nsew signal tristate
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 587 nsew signal tristate
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 588 nsew signal tristate
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 589 nsew signal tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew signal tristate
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 591 nsew signal tristate
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 592 nsew signal tristate
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 593 nsew signal tristate
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 594 nsew signal tristate
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 595 nsew signal tristate
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 596 nsew signal tristate
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 597 nsew signal tristate
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 598 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 599 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 600 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 601 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 602 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 603 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 604 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 606 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 607 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 608 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 609 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 610 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 611 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 612 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 613 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 614 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 615 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 616 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 618 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 619 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
