* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_ls__decap_8 abstract view
.subckt sky130_fd_sc_ls__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__fill_1 abstract view
.subckt sky130_fd_sc_ls__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__fill_diode_2 abstract view
.subckt sky130_fd_sc_ls__fill_diode_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__decap_4 abstract view
.subckt sky130_fd_sc_ls__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__diode_2 abstract view
.subckt sky130_fd_sc_ls__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__clkbuf_2 abstract view
.subckt sky130_fd_sc_ls__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_ls__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__conb_1 abstract view
.subckt sky130_fd_sc_ls__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__clkbuf_1 abstract view
.subckt sky130_fd_sc_ls__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 vdd gnd Y B A C
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 vdd gnd Y A
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 vdd gnd Y A
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 vdd gnd Y A
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__buf_2 abstract view
.subckt sky130_fd_sc_ls__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 vdd gnd Y A
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 vdd gnd Y A
.ends

* Black-box entry subcircuit for INV abstract view
.subckt INV vdd gnd Y A
.ends

* Black-box entry subcircuit for sky130_fd_sc_ls__clkbuf_4 abstract view
.subckt sky130_fd_sc_ls__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 vdd gnd Y A
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 vdd gnd Y B C A D
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 vdd gnd Y A
.ends

* Black-box entry subcircuit for AND2X1 abstract view
.subckt AND2X1 vdd gnd Y A B
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 vdd gnd Y B A
.ends

* Black-box entry subcircuit for HAX1 abstract view
.subckt HAX1 vdd gnd YS YC B A
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i vccd1 vssd1
+ vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 vssa2_uq0 vssa1_uq0 vssd2_uq0 vdda2_uq0 vdda1_uq0
+ vccd2_uq0
XFILLER_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_213 _208_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_202 _068_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_224 _218_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput401 _221_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_ls__clkbuf_2
Xoutput434 _056_/LO vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_ls__clkbuf_2
Xoutput423 _051_/LO vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_ls__clkbuf_2
Xoutput412 _046_/LO vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_ls__clkbuf_2
Xoutput456 _169_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_ls__clkbuf_2
Xoutput478 _074_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_ls__clkbuf_2
Xoutput445 _159_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_ls__clkbuf_2
Xoutput467 _179_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput489 _084_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_927 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_916 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_905 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_702 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_735 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_200_ vssd1 vssd1 vccd1 vccd1 _200_/HI _200_/LO sky130_fd_sc_ls__conb_1
XFILLER_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_131_ vssd1 vssd1 vccd1 vccd1 _131_/HI _131_/LO sky130_fd_sc_ls__conb_1
XPHY_779 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_062_ vssd1 vssd1 vccd1 vccd1 _062_/HI _062_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_510 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_598 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_114_ vssd1 vssd1 vccd1 vccd1 _114_/HI _114_/LO sky130_fd_sc_ls__conb_1
X_045_ vssd1 vssd1 vccd1 vccd1 _045_/HI _045_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput301 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input301/X sky130_fd_sc_ls__clkbuf_1
Xinput312 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 input312/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput345 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 input345/X sky130_fd_sc_ls__clkbuf_1
Xinput334 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input334/X sky130_fd_sc_ls__clkbuf_1
Xinput323 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 input323/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput367 wbs_we_i vssd1 vssd1 vccd1 vccd1 input367/X sky130_fd_sc_ls__clkbuf_1
Xinput356 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input356/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_340 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_362 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_5 _020_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_028_ vssd1 vssd1 vccd1 vccd1 _028_/HI _028_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput120 la_data_in[58] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput131 la_data_in[68] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_ls__clkbuf_1
Xinput142 la_data_in[78] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_ls__clkbuf_1
Xinput153 la_data_in[88] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_ls__clkbuf_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput186 la_oen[117] vssd1 vssd1 vccd1 vccd1 input186/X sky130_fd_sc_ls__clkbuf_1
Xinput175 la_oen[107] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_ls__clkbuf_1
Xinput164 la_data_in[98] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput197 la_oen[127] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_170 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_192 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_181 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_225 _191_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_203 _188_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_214 _208_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput402 _016_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_ls__clkbuf_2
Xoutput424 INV/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_ls__clkbuf_2
Xoutput413 BUFX2/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_ls__clkbuf_2
Xoutput435 _057_/LO vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_ls__clkbuf_2
Xoutput446 _160_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_ls__clkbuf_2
Xoutput457 _170_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_ls__clkbuf_2
Xoutput468 _180_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_ls__clkbuf_2
Xoutput479 _075_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_ls__clkbuf_2
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_917 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_906 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_939 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_703 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_725 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_747 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_130_ vssd1 vssd1 vccd1 vccd1 _130_/HI _130_/LO sky130_fd_sc_ls__conb_1
XFILLER_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_061_ vssd1 vssd1 vccd1 vccd1 _061_/HI _061_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_500 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_511 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_533 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_555 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_113_ vssd1 vssd1 vccd1 vccd1 _113_/HI _113_/LO sky130_fd_sc_ls__conb_1
X_044_ vssd1 vssd1 vccd1 vccd1 _044_/HI _044_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput302 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input302/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput313 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 input313/X sky130_fd_sc_ls__clkbuf_1
Xinput324 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 input324/X sky130_fd_sc_ls__clkbuf_1
Xinput335 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 input335/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput346 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 input346/X sky130_fd_sc_ls__clkbuf_1
Xinput357 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input357/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_330 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_352 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_363 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_396 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_6 _000_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
X_027_ vssd1 vssd1 vccd1 vccd1 _027_/HI _027_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput110 la_data_in[49] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput143 la_data_in[79] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_ls__clkbuf_1
Xinput121 la_data_in[59] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput132 la_data_in[69] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_ls__clkbuf_1
Xinput154 la_data_in[89] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_ls__clkbuf_1
Xinput187 la_oen[118] vssd1 vssd1 vccd1 vccd1 input187/X sky130_fd_sc_ls__clkbuf_1
Xinput176 la_oen[108] vssd1 vssd1 vccd1 vccd1 input176/X sky130_fd_sc_ls__clkbuf_1
Xinput165 la_data_in[99] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput198 la_oen[12] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_ls__clkbuf_1
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_171 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_193 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_182 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_204 _188_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_215 _212_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_226 _191_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput425 _052_/LO vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_ls__clkbuf_2
Xoutput414 _047_/LO vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_ls__clkbuf_2
Xoutput403 _017_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_ls__clkbuf_2
Xoutput436 _058_/LO vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_ls__clkbuf_2
Xoutput447 _161_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_ls__clkbuf_2
Xoutput469 _181_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_ls__clkbuf_2
Xoutput458 _171_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_918 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_907 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_929 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_704 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_737 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_060_ vssd1 vssd1 vccd1 vccd1 _060_/HI _060_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_189_ vssd1 vssd1 vccd1 vccd1 _189_/HI _189_/LO sky130_fd_sc_ls__conb_1
XFILLER_43_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_501 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_512 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_589 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_112_ vssd1 vssd1 vccd1 vccd1 _112_/HI _112_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_043_ vssd1 vssd1 vccd1 vccd1 _043_/HI _043_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput303 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input303/X sky130_fd_sc_ls__clkbuf_1
Xinput336 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 input336/X sky130_fd_sc_ls__clkbuf_1
Xinput325 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 input325/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput314 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 input314/X sky130_fd_sc_ls__clkbuf_1
Xinput347 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 input347/X sky130_fd_sc_ls__clkbuf_1
Xinput358 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input358/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_320 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_342 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_353 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_397 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_7 _000_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_026_ vssd1 vssd1 vccd1 vccd1 _026_/HI _026_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput111 la_data_in[4] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_ls__clkbuf_1
Xinput100 la_data_in[3] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_ls__clkbuf_1
Xinput133 la_data_in[6] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_ls__clkbuf_1
Xinput122 la_data_in[5] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput144 la_data_in[7] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput177 la_oen[109] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_ls__clkbuf_1
Xinput155 la_data_in[8] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_ls__clkbuf_1
Xinput166 la_data_in[9] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput188 la_oen[119] vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_ls__clkbuf_1
Xinput199 la_oen[13] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_ls__clkbuf_1
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_172 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_194 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_183 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_009_ vssd1 vssd1 vccd1 vccd1 _009_/HI _009_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_205 _199_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_216 _212_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput415 BUFX4/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_ls__clkbuf_2
Xoutput404 _018_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_ls__clkbuf_2
Xoutput426 INVX1/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_ls__clkbuf_2
Xoutput437 _037_/LO vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_ls__clkbuf_2
Xoutput448 _162_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_ls__clkbuf_2
Xoutput459 _172_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_ls__clkbuf_2
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_908 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_705 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_738 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_188_ vssd1 vssd1 vccd1 vccd1 _188_/HI _188_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_502 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_546 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_111_ vssd1 vssd1 vccd1 vccd1 _111_/HI _111_/LO sky130_fd_sc_ls__conb_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_042_ vssd1 vssd1 vccd1 vccd1 _042_/HI _042_/LO sky130_fd_sc_ls__conb_1
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput304 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 input304/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput326 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 input326/X sky130_fd_sc_ls__clkbuf_1
Xinput315 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 input315/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput348 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 input348/X sky130_fd_sc_ls__clkbuf_1
Xinput359 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input359/X sky130_fd_sc_ls__clkbuf_1
Xinput337 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 input337/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_310 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_321 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_343 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_354 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_387 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_8 _001_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_025_ vssd1 vssd1 vccd1 vccd1 _025_/HI _025_/LO sky130_fd_sc_ls__conb_1
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput101 la_data_in[40] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_ls__clkbuf_1
XFILLER_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput145 la_data_in[80] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_ls__clkbuf_1
Xinput112 la_data_in[50] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_ls__clkbuf_1
Xinput123 la_data_in[60] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_ls__clkbuf_1
Xinput134 la_data_in[70] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_ls__clkbuf_1
XFILLER_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput167 la_oen[0] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_ls__clkbuf_1
Xinput156 la_data_in[90] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_ls__clkbuf_1
Xinput178 la_oen[10] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_ls__clkbuf_1
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput189 la_oen[11] vssd1 vssd1 vccd1 vccd1 input189/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_173 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_184 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_195 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_008_ vssd1 vssd1 vccd1 vccd1 _008_/HI _008_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_206 _199_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_217 _214_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput416 _048_/LO vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_ls__clkbuf_2
Xoutput405 _222_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_ls__clkbuf_2
Xoutput427 _053_/LO vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_ls__clkbuf_2
Xoutput438 _038_/LO vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_ls__clkbuf_2
Xoutput449 _163_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_ls__clkbuf_2
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_909 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_706 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_187_ vssd1 vssd1 vccd1 vccd1 _187_/HI _187_/LO sky130_fd_sc_ls__conb_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_503 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_536 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_110_ vssd1 vssd1 vccd1 vccd1 _110_/HI _110_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_041_ vssd1 vssd1 vccd1 vccd1 _041_/HI _041_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput327 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 input327/X sky130_fd_sc_ls__clkbuf_1
Xinput305 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 input305/X sky130_fd_sc_ls__clkbuf_1
Xinput316 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 input316/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput349 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 input349/X sky130_fd_sc_ls__clkbuf_1
Xinput338 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 input338/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_300 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_311 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_388 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_399 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_9 _001_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
X_024_ vssd1 vssd1 vccd1 vccd1 _024_/HI _024_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput102 la_data_in[41] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_ls__clkbuf_1
Xinput135 la_data_in[71] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_ls__clkbuf_1
Xinput113 la_data_in[51] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_ls__clkbuf_1
Xinput124 la_data_in[61] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_ls__clkbuf_1
Xinput168 la_oen[100] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput146 la_data_in[81] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_ls__clkbuf_1
Xinput157 la_data_in[91] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput179 la_oen[110] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_185 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_174 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_196 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_007_ vssd1 vssd1 vccd1 vccd1 _007_/HI _007_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_207 _201_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_218 _214_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput417 _036_/LO vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_ls__clkbuf_2
Xoutput406 _035_/LO vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput439 AND2X2/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_ls__clkbuf_2
Xoutput428 AND2X1/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_ls__clkbuf_2
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XAOI21X1 vccd1 vssd1 AOI21X1/Y input36/X input37/X input35/X AOI21X1
XFILLER_10_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_707 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_729 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_186_ vssd1 vssd1 vccd1 vccd1 _186_/HI _186_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_504 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_537 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_040_ vssd1 vssd1 vccd1 vccd1 _040_/HI _040_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_169_ vssd1 vssd1 vccd1 vccd1 _169_/HI _169_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput306 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 input306/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput317 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input317/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput339 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 input339/X sky130_fd_sc_ls__clkbuf_1
Xinput328 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 input328/X sky130_fd_sc_ls__clkbuf_1
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_301 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_312 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_334 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_378 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_023_ vssd1 vssd1 vccd1 vccd1 _023_/HI _023_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_890 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput103 la_data_in[42] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_ls__clkbuf_1
Xinput114 la_data_in[52] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_ls__clkbuf_1
Xinput125 la_data_in[62] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_ls__clkbuf_1
Xinput136 la_data_in[72] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput169 la_oen[101] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_ls__clkbuf_1
Xinput158 la_data_in[92] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_ls__clkbuf_1
Xinput147 la_data_in[82] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_ls__clkbuf_1
XFILLER_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_164 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_175 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_186 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_197 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_006_ vssd1 vssd1 vccd1 vccd1 _006_/HI _006_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_219 _215_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_208 _201_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput407 _042_/LO vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_ls__clkbuf_2
Xoutput429 INVX2/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_ls__clkbuf_2
Xoutput418 CLKBUF1/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_ls__clkbuf_2
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_71_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_708 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_719 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_185_ vssd1 vssd1 vccd1 vccd1 _185_/HI _185_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_505 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_527 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_538 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput590 _213_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_168_ vssd1 vssd1 vccd1 vccd1 _168_/HI _168_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_099_ vssd1 vssd1 vccd1 vccd1 _099_/HI _099_/LO sky130_fd_sc_ls__conb_1
XFILLER_34_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput318 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input318/X sky130_fd_sc_ls__clkbuf_1
Xinput307 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 input307/X sky130_fd_sc_ls__clkbuf_1
Xinput329 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input329/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_302 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_335 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_368 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_379 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_022_ vssd1 vssd1 vccd1 vccd1 _022_/HI _022_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_880 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_891 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput104 la_data_in[43] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_ls__clkbuf_1
Xinput115 la_data_in[53] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_ls__clkbuf_1
Xinput126 la_data_in[63] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_ls__clkbuf_1
XFILLER_56_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput148 la_data_in[83] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_ls__clkbuf_1
Xinput137 la_data_in[73] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_ls__clkbuf_1
Xinput159 la_data_in[93] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_165 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_176 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_187 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_198 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_005_ vssd1 vssd1 vccd1 vccd1 _005_/HI _005_/LO sky130_fd_sc_ls__conb_1
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_209 _206_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput408 _043_/LO vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_ls__clkbuf_2
Xoutput419 _049_/LO vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_ls__clkbuf_2
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_709 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XINVX1 vccd1 vssd1 INVX1/Y INVX1/A INVX1
XFILLER_73_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_184_ vssd1 vssd1 vccd1 vccd1 _184_/HI _184_/LO sky130_fd_sc_ls__conb_1
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_506 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_528 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput580 _204_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_ls__clkbuf_2
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput591 _214_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_167_ vssd1 vssd1 vccd1 vccd1 _167_/HI _167_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_098_ vssd1 vssd1 vccd1 vccd1 _098_/HI _098_/LO sky130_fd_sc_ls__conb_1
XFILLER_27_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput308 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 input308/X sky130_fd_sc_ls__clkbuf_1
Xinput319 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 input319/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_303 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_336 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_021_ vssd1 vssd1 vccd1 vccd1 _021_/HI _021_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_881 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_892 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_219_ vssd1 vssd1 vccd1 vccd1 _219_/HI _219_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput116 la_data_in[54] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_ls__clkbuf_1
Xinput105 la_data_in[44] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput127 la_data_in[64] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_ls__clkbuf_1
Xinput138 la_data_in[74] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_ls__clkbuf_1
Xinput149 la_data_in[84] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_ls__clkbuf_1
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_166 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_199 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_188 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_177 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_004_ vssd1 vssd1 vccd1 vccd1 _004_/HI _004_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput409 _044_/LO vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_ls__clkbuf_2
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XINVX2 vccd1 vssd1 INVX2/Y INVX2/A INVX2
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_183_ vssd1 vssd1 vccd1 vccd1 _183_/HI _183_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_507 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_518 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_529 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput570 _158_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_ls__clkbuf_2
Xoutput581 _205_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_ls__clkbuf_2
Xoutput592 _215_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_ls__clkbuf_2
XFILLER_75_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_166_ vssd1 vssd1 vccd1 vccd1 _166_/HI _166_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_097_ vssd1 vssd1 vccd1 vccd1 _097_/HI _097_/LO sky130_fd_sc_ls__conb_1
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_190 _143_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput309 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 input309/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_304 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_326 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_359 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_020_ vssd1 vssd1 vccd1 vccd1 _020_/HI _020_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_871 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_893 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_218_ vssd1 vssd1 vccd1 vccd1 _218_/HI _218_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_149_ vssd1 vssd1 vccd1 vccd1 _149_/HI _149_/LO sky130_fd_sc_ls__conb_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput106 la_data_in[45] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_ls__clkbuf_1
Xinput117 la_data_in[55] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_ls__clkbuf_1
Xinput128 la_data_in[65] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_ls__clkbuf_1
Xinput139 la_data_in[75] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_167 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_189 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_178 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_90 _037_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
X_003_ vssd1 vssd1 vccd1 vccd1 _003_/HI _003_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_690 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_182_ vssd1 vssd1 vccd1 vccd1 _182_/HI _182_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_508 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_519 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput571 _068_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_ls__clkbuf_2
Xoutput560 _067_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput593 _216_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_ls__clkbuf_2
Xoutput582 _206_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_165_ vssd1 vssd1 vccd1 vccd1 _165_/HI _165_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_096_ vssd1 vssd1 vccd1 vccd1 _096_/HI _096_/LO sky130_fd_sc_ls__conb_1
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_191 _147_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_180 _137_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_305 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_316 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput390 _220_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_ls__clkbuf_2
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_872 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_850 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_894 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_217_ vssd1 vssd1 vccd1 vccd1 _217_/HI _217_/LO sky130_fd_sc_ls__conb_1
X_148_ vssd1 vssd1 vccd1 vccd1 _148_/HI _148_/LO sky130_fd_sc_ls__conb_1
X_079_ vssd1 vssd1 vccd1 vccd1 _079_/HI _079_/LO sky130_fd_sc_ls__conb_1
XFILLER_32_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput107 la_data_in[46] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_ls__clkbuf_1
Xinput118 la_data_in[56] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_ls__clkbuf_1
Xinput129 la_data_in[66] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_168 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_179 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_002_ vssd1 vssd1 vccd1 vccd1 _002_/HI _002_/LO sky130_fd_sc_ls__conb_1
XANTENNA_91 AND2X2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_80 INVX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_680 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_691 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput290 la_oen[96] vssd1 vssd1 vccd1 vccd1 input290/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XINVX4 vccd1 vssd1 INVX4/Y INVX4/A INVX4
XFILLER_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_181_ vssd1 vssd1 vccd1 vccd1 _181_/HI _181_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_509 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput550 _139_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_ls__clkbuf_2
Xoutput572 _187_/LO vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_ls__clkbuf_2
Xoutput561 _149_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_ls__clkbuf_2
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput594 _217_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_ls__clkbuf_2
Xoutput583 _207_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_ls__clkbuf_2
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_164_ vssd1 vssd1 vccd1 vccd1 _164_/HI _164_/LO sky130_fd_sc_ls__conb_1
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_095_ vssd1 vssd1 vccd1 vccd1 _095_/HI _095_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_170 _124_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_192 _147_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_181 _137_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_306 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_317 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_339 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput380 _024_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_ls__clkbuf_2
Xoutput391 _029_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_ls__clkbuf_2
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_862 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_851 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_216_ vssd1 vssd1 vccd1 vccd1 _216_/HI _216_/LO sky130_fd_sc_ls__conb_1
X_147_ vssd1 vssd1 vccd1 vccd1 _147_/HI _147_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_078_ vssd1 vssd1 vccd1 vccd1 _078_/HI _078_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput108 la_data_in[47] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_ls__clkbuf_1
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput119 la_data_in[57] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_ls__clkbuf_1
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_169 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_81 INVX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_70 INV/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_92 AND2X2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
X_001_ vssd1 vssd1 vccd1 vccd1 _001_/HI _001_/LO sky130_fd_sc_ls__conb_1
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_670 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_681 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput90 la_data_in[30] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_ls__clkbuf_1
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput280 la_oen[87] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput291 la_oen[97] vssd1 vssd1 vccd1 vccd1 input291/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_180_ vssd1 vssd1 vccd1 vccd1 _180_/HI _180_/LO sky130_fd_sc_ls__conb_1
XFILLER_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput562 _150_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_ls__clkbuf_2
Xoutput551 _140_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_ls__clkbuf_2
Xoutput540 _130_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_ls__clkbuf_2
Xoutput595 _190_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_ls__clkbuf_2
Xoutput573 _188_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_ls__clkbuf_2
Xoutput584 _189_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_163_ vssd1 vssd1 vccd1 vccd1 _163_/HI _163_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_094_ vssd1 vssd1 vccd1 vccd1 _094_/HI _094_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_160 _107_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_171 _125_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_193 _148_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_182 _138_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_307 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_318 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_329 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput370 _020_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_ls__clkbuf_2
Xoutput392 _010_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_ls__clkbuf_2
Xoutput381 _005_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_863 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_830 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_896 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_215_ vssd1 vssd1 vccd1 vccd1 _215_/HI _215_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_146_ vssd1 vssd1 vccd1 vccd1 _146_/HI _146_/LO sky130_fd_sc_ls__conb_1
X_077_ vssd1 vssd1 vccd1 vccd1 _077_/HI _077_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput109 la_data_in[48] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_ls__clkbuf_1
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_71 INV/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_60 _050_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_93 _039_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
X_000_ vssd1 vssd1 vccd1 vccd1 _000_/HI _000_/LO sky130_fd_sc_ls__conb_1
XANTENNA_82 INVX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_660 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_129_ vssd1 vssd1 vccd1 vccd1 _129_/HI _129_/LO sky130_fd_sc_ls__conb_1
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput80 la_data_in[21] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_ls__clkbuf_1
Xinput91 la_data_in[31] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_ls__clkbuf_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_490 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput281 la_oen[88] vssd1 vssd1 vccd1 vccd1 input281/X sky130_fd_sc_ls__clkbuf_1
Xinput270 la_oen[78] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_ls__clkbuf_1
Xinput292 la_oen[98] vssd1 vssd1 vccd1 vccd1 input292/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput541 _131_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_ls__clkbuf_2
Xoutput530 _121_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_ls__clkbuf_2
Xoutput563 _151_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_ls__clkbuf_2
Xoutput552 _141_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput596 _218_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_ls__clkbuf_2
Xoutput585 _208_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_ls__clkbuf_2
Xoutput574 _198_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_ls__clkbuf_2
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_162_ vssd1 vssd1 vccd1 vccd1 _162_/HI _162_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_093_ vssd1 vssd1 vccd1 vccd1 _093_/HI _093_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_150 _096_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_161 _110_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_194 _148_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_172 _125_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_183 _138_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_ls__buf_2
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_308 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_319 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput371 _000_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_ls__clkbuf_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput393 _030_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_ls__clkbuf_2
Xoutput382 _006_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_820 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_853 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_214_ vssd1 vssd1 vccd1 vccd1 _214_/HI _214_/LO sky130_fd_sc_ls__conb_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_145_ vssd1 vssd1 vccd1 vccd1 _145_/HI _145_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_076_ vssd1 vssd1 vccd1 vccd1 _076_/HI _076_/LO sky130_fd_sc_ls__conb_1
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_50 _046_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_83 INVX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_61 HAX1/YS vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_72 _052_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_94 _039_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_650 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_672 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_128_ vssd1 vssd1 vccd1 vccd1 _128_/HI _128_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_059_ vssd1 vssd1 vccd1 vccd1 _059_/HI _059_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput81 la_data_in[22] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_ls__clkbuf_1
Xinput70 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_ls__clkbuf_1
Xinput92 la_data_in[32] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_ls__clkbuf_1
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_480 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_78_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_491 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput271 la_oen[79] vssd1 vssd1 vccd1 vccd1 input271/X sky130_fd_sc_ls__clkbuf_1
Xinput260 la_oen[69] vssd1 vssd1 vccd1 vccd1 input260/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput293 la_oen[99] vssd1 vssd1 vccd1 vccd1 input293/X sky130_fd_sc_ls__clkbuf_1
Xinput282 la_oen[89] vssd1 vssd1 vccd1 vccd1 input282/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput520 _112_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_ls__clkbuf_2
Xoutput553 _142_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_ls__clkbuf_2
Xoutput542 _132_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_ls__clkbuf_2
Xoutput531 _122_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_ls__clkbuf_2
Xoutput564 _152_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_ls__clkbuf_2
Xoutput586 _209_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_ls__clkbuf_2
Xoutput575 _199_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput597 _219_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_ls__clkbuf_2
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_161_ vssd1 vssd1 vccd1 vccd1 _161_/HI _161_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_092_ vssd1 vssd1 vccd1 vccd1 _092_/HI _092_/LO sky130_fd_sc_ls__conb_1
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_140 _082_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_151 _098_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_184 _139_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_173 _126_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_162 _112_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_195 _151_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_ls__buf_2
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_309 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput383 _025_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_ls__clkbuf_2
Xoutput394 _011_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_ls__clkbuf_2
Xoutput372 _001_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_ls__clkbuf_2
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_810 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_854 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_887 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_213_ vssd1 vssd1 vccd1 vccd1 _213_/HI _213_/LO sky130_fd_sc_ls__conb_1
XPHY_898 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_144_ vssd1 vssd1 vccd1 vccd1 _144_/HI _144_/LO sky130_fd_sc_ls__conb_1
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_075_ vssd1 vssd1 vccd1 vccd1 _075_/HI _075_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_40 _035_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_73 _052_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_62 HAX1/YS vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_84 INVX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_51 BUFX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_95 _041_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_640 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_673 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_127_ vssd1 vssd1 vccd1 vccd1 _127_/HI _127_/LO sky130_fd_sc_ls__conb_1
X_058_ vssd1 vssd1 vccd1 vccd1 _058_/HI _058_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput60 la_data_in[119] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_ls__clkbuf_1
Xinput71 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_ls__clkbuf_1
Xinput82 la_data_in[23] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_ls__clkbuf_1
Xinput93 la_data_in[33] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_ls__clkbuf_1
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_470 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_45_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput272 la_oen[7] vssd1 vssd1 vccd1 vccd1 input272/X sky130_fd_sc_ls__clkbuf_1
Xinput250 la_oen[5] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_ls__clkbuf_1
Xinput261 la_oen[6] vssd1 vssd1 vccd1 vccd1 input261/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput294 la_oen[9] vssd1 vssd1 vccd1 vccd1 input294/X sky130_fd_sc_ls__clkbuf_1
Xinput283 la_oen[8] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XINVX8 vccd1 vssd1 INVX8/Y INVX8/A INVX8
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_70_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput510 _103_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_ls__clkbuf_2
Xoutput554 _143_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_ls__clkbuf_2
Xoutput543 _133_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_ls__clkbuf_2
Xoutput532 _123_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_ls__clkbuf_2
Xoutput521 _113_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_ls__clkbuf_2
Xoutput587 _210_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_ls__clkbuf_2
Xoutput565 _153_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_ls__clkbuf_2
Xoutput576 _200_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput598 _191_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_ls__clkbuf_2
XFILLER_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_160_ vssd1 vssd1 vccd1 vccd1 _160_/HI _160_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_091_ vssd1 vssd1 vccd1 vccd1 _091_/HI _091_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_141 _083_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_152 _098_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_130 _183_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_163 _114_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_185 _139_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_174 _126_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_196 _151_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_ls__buf_2
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput395 _031_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_ls__clkbuf_2
Xoutput384 _026_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_ls__clkbuf_2
Xoutput373 _021_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_811 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_800 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_822 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_212_ vssd1 vssd1 vccd1 vccd1 _212_/HI _212_/LO sky130_fd_sc_ls__conb_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_143_ vssd1 vssd1 vccd1 vccd1 _143_/HI _143_/LO sky130_fd_sc_ls__conb_1
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_074_ vssd1 vssd1 vccd1 vccd1 _074_/HI _074_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_41 _042_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_30 _010_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_74 _052_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_63 HAX1/YS vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_52 BUFX2/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_96 _041_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_85 _055_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_630 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_663 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_696 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_126_ vssd1 vssd1 vccd1 vccd1 _126_/HI _126_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_057_ vssd1 vssd1 vccd1 vccd1 _057_/HI _057_/LO sky130_fd_sc_ls__conb_1
XFILLER_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput50 la_data_in[10] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_ls__clkbuf_1
Xinput61 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_ls__clkbuf_1
Xinput72 la_data_in[14] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_ls__clkbuf_1
Xinput94 la_data_in[34] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_ls__clkbuf_1
Xinput83 la_data_in[24] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_460 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_482 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_109_ vssd1 vssd1 vccd1 vccd1 _109_/HI _109_/LO sky130_fd_sc_ls__conb_1
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput262 la_oen[70] vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_ls__clkbuf_1
Xinput251 la_oen[60] vssd1 vssd1 vccd1 vccd1 input251/X sky130_fd_sc_ls__clkbuf_1
Xinput240 la_oen[50] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput284 la_oen[90] vssd1 vssd1 vccd1 vccd1 input284/X sky130_fd_sc_ls__clkbuf_1
Xinput273 la_oen[80] vssd1 vssd1 vccd1 vccd1 input273/X sky130_fd_sc_ls__clkbuf_1
Xinput295 wb_clk_i vssd1 vssd1 vccd1 vccd1 input295/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_290 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput511 _104_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_ls__clkbuf_2
Xoutput500 _094_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_ls__clkbuf_2
Xoutput533 _124_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_ls__clkbuf_2
Xoutput544 _134_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_ls__clkbuf_2
Xoutput522 _114_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_ls__clkbuf_2
Xoutput566 _154_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_ls__clkbuf_2
Xoutput555 _144_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput577 _201_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_ls__clkbuf_2
Xoutput588 _211_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_ls__clkbuf_2
Xoutput599 _192_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_ls__clkbuf_2
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_090_ vssd1 vssd1 vccd1 vccd1 _090_/HI _090_/LO sky130_fd_sc_ls__conb_1
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_131 _186_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_142 _083_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_120 _174_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_175 _131_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_153 _062_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_164 _114_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_186 _140_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_197 _153_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_ls__buf_2
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput396 _032_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_ls__clkbuf_2
Xoutput385 _007_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_ls__clkbuf_2
Xoutput374 _002_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_ls__clkbuf_2
XFILLER_19_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_801 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_845 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_812 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_878 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_856 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_211_ vssd1 vssd1 vccd1 vccd1 _211_/HI _211_/LO sky130_fd_sc_ls__conb_1
XPHY_889 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_142_ vssd1 vssd1 vccd1 vccd1 _142_/HI _142_/LO sky130_fd_sc_ls__conb_1
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_11_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_073_ vssd1 vssd1 vccd1 vccd1 _073_/HI _073_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_31 _010_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_20 _025_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_42 _042_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_53 BUFX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_64 HAX1/YC vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_75 INVX1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_86 _055_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_97 AOI21X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_79_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_620 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_631 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_642 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_664 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_697 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_125_ vssd1 vssd1 vccd1 vccd1 _125_/HI _125_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_056_ vssd1 vssd1 vccd1 vccd1 _056_/HI _056_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput40 la_data_in[100] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_ls__clkbuf_1
Xinput62 la_data_in[120] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_ls__clkbuf_1
Xinput73 la_data_in[15] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_ls__clkbuf_1
Xinput51 la_data_in[110] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_ls__clkbuf_1
Xinput84 la_data_in[25] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_ls__clkbuf_1
Xinput95 la_data_in[35] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_ls__clkbuf_1
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_450 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_108_ vssd1 vssd1 vccd1 vccd1 _108_/HI _108_/LO sky130_fd_sc_ls__conb_1
X_039_ vssd1 vssd1 vccd1 vccd1 _039_/HI _039_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput263 la_oen[71] vssd1 vssd1 vccd1 vccd1 input263/X sky130_fd_sc_ls__clkbuf_1
Xinput252 la_oen[61] vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_ls__clkbuf_1
Xinput241 la_oen[51] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_ls__clkbuf_1
Xinput230 la_oen[41] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput285 la_oen[91] vssd1 vssd1 vccd1 vccd1 input285/X sky130_fd_sc_ls__clkbuf_1
Xinput274 la_oen[81] vssd1 vssd1 vccd1 vccd1 input274/X sky130_fd_sc_ls__clkbuf_1
Xinput296 wb_rst_i vssd1 vssd1 vccd1 vccd1 input296/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_280 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_291 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_76_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_72_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput501 _095_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_ls__clkbuf_2
Xoutput523 _115_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_ls__clkbuf_2
Xoutput545 _135_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_ls__clkbuf_2
Xoutput534 _125_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_ls__clkbuf_2
Xoutput512 _105_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_ls__clkbuf_2
Xoutput567 _155_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_ls__clkbuf_2
Xoutput556 _145_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_ls__clkbuf_2
Xoutput578 _202_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput589 _212_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_143 _085_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_121 _175_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_110 _167_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_132 _186_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_165 _121_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_176 _131_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_154 _062_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_198 _153_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_187 _140_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_ls__buf_2
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XBUFX2 vccd1 vssd1 BUFX2/Y BUFX2/A BUFX2
Xoutput386 _027_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_ls__clkbuf_2
Xoutput375 _022_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_ls__clkbuf_2
Xoutput397 _033_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_802 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_835 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_813 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_879 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_210_ vssd1 vssd1 vccd1 vccd1 _210_/HI _210_/LO sky130_fd_sc_ls__conb_1
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_141_ vssd1 vssd1 vccd1 vccd1 _141_/HI _141_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_072_ vssd1 vssd1 vccd1 vccd1 _072_/HI _072_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_21 _025_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_32 _034_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_10 _021_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_54 BUFX4/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_65 HAX1/YC vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_43 _044_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_98 AOI21X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_76 INVX1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_87 INVX8/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_75_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_610 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_621 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_654 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_687 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_698 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_124_ vssd1 vssd1 vccd1 vccd1 _124_/HI _124_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_055_ vssd1 vssd1 vccd1 vccd1 _055_/HI _055_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput30 io_in[36] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_ls__clkbuf_1
Xinput63 la_data_in[121] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_ls__clkbuf_1
Xinput41 la_data_in[101] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_ls__clkbuf_1
Xinput52 la_data_in[111] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_ls__clkbuf_1
Xinput96 la_data_in[36] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_ls__clkbuf_1
Xinput74 la_data_in[16] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_ls__clkbuf_1
Xinput85 la_data_in[26] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_ls__clkbuf_1
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_440 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_107_ vssd1 vssd1 vccd1 vccd1 _107_/HI _107_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_038_ vssd1 vssd1 vccd1 vccd1 _038_/HI _038_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput220 la_oen[32] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput253 la_oen[62] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_ls__clkbuf_1
Xinput242 la_oen[52] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_ls__clkbuf_1
Xinput231 la_oen[42] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput286 la_oen[92] vssd1 vssd1 vccd1 vccd1 input286/X sky130_fd_sc_ls__clkbuf_1
Xinput275 la_oen[82] vssd1 vssd1 vccd1 vccd1 input275/X sky130_fd_sc_ls__clkbuf_1
Xinput264 la_oen[72] vssd1 vssd1 vccd1 vccd1 input264/X sky130_fd_sc_ls__clkbuf_1
Xinput297 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input297/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_270 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_281 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_292 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput502 _096_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_ls__clkbuf_2
Xoutput535 _126_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_ls__clkbuf_2
Xoutput524 _116_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_ls__clkbuf_2
Xoutput513 _106_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_ls__clkbuf_2
Xoutput568 _156_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_ls__clkbuf_2
Xoutput557 _146_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_ls__clkbuf_2
Xoutput546 _136_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput579 _203_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_ls__clkbuf_2
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_100 _159_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_133 _075_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_111 _168_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_122 _175_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_166 _121_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_144 _085_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_155 _101_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_188 _141_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_199 _155_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_177 _134_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_ls__clkbuf_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput387 _008_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_ls__clkbuf_2
Xoutput376 _003_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_ls__clkbuf_2
Xoutput398 _034_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_836 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_803 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_847 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_140_ vssd1 vssd1 vccd1 vccd1 _140_/HI _140_/LO sky130_fd_sc_ls__conb_1
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_51_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_071_ vssd1 vssd1 vccd1 vccd1 _071_/HI _071_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_22 _025_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_11 _021_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_66 HAX1/YC vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_44 _044_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_33 _014_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_55 _036_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_88 INVX8/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_77 INVX1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XINV vccd1 vssd1 INV/Y INV/A INV
XFILLER_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_99 _159_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_600 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_622 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_655 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_123_ vssd1 vssd1 vccd1 vccd1 _123_/HI _123_/LO sky130_fd_sc_ls__conb_1
X_054_ vssd1 vssd1 vccd1 vccd1 _054_/HI _054_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput20 io_in[27] vssd1 vssd1 vccd1 vccd1 INVX1/A sky130_fd_sc_ls__clkbuf_4
Xinput31 io_in[37] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_ls__clkbuf_1
Xinput64 la_data_in[122] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_ls__clkbuf_1
Xinput53 la_data_in[112] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_ls__clkbuf_1
Xinput42 la_data_in[102] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_ls__clkbuf_1
Xinput97 la_data_in[37] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_ls__clkbuf_1
Xinput75 la_data_in[17] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_ls__clkbuf_1
Xinput86 la_data_in[27] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_ls__clkbuf_1
XFILLER_6_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_16_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_430 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1040 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_496 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_106_ vssd1 vssd1 vccd1 vccd1 _106_/HI _106_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_037_ vssd1 vssd1 vccd1 vccd1 _037_/HI _037_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput210 la_oen[23] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput254 la_oen[63] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_ls__clkbuf_1
Xinput221 la_oen[33] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_ls__clkbuf_1
Xinput243 la_oen[53] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_ls__clkbuf_1
Xinput232 la_oen[43] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput287 la_oen[93] vssd1 vssd1 vccd1 vccd1 input287/X sky130_fd_sc_ls__clkbuf_1
Xinput276 la_oen[83] vssd1 vssd1 vccd1 vccd1 input276/X sky130_fd_sc_ls__clkbuf_1
Xinput265 la_oen[73] vssd1 vssd1 vccd1 vccd1 input265/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput298 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input298/X sky130_fd_sc_ls__clkbuf_1
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_260 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_271 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_293 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput536 _127_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_ls__clkbuf_2
Xoutput525 _117_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_ls__clkbuf_2
Xoutput514 _107_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_ls__clkbuf_2
Xoutput503 _097_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_ls__clkbuf_2
Xoutput569 _157_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_ls__clkbuf_2
Xoutput558 _147_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_ls__clkbuf_2
Xoutput547 _137_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_112 _168_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_101 _159_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_134 _075_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_123 _177_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_167 _122_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_145 _087_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_156 _101_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_189 _141_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_178 _134_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 BUFX2/A sky130_fd_sc_ls__buf_2
XFILLER_64_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XBUFX4 vccd1 vssd1 BUFX4/Y BUFX4/A BUFX4
Xoutput377 _023_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_ls__clkbuf_2
Xoutput388 _028_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_ls__clkbuf_2
Xoutput399 _014_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_ls__clkbuf_2
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_804 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_070_ vssd1 vssd1 vccd1 vccd1 _070_/HI _070_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_199_ vssd1 vssd1 vccd1 vccd1 _199_/HI _199_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_23 _026_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_12 _022_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_34 _014_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_56 _036_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_45 _045_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_78 AND2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_89 _037_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_67 _051_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_601 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_612 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_645 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_689 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_122_ vssd1 vssd1 vccd1 vccd1 _122_/HI _122_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_053_ vssd1 vssd1 vccd1 vccd1 _053_/HI _053_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_3_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_78_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput21 io_in[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_ls__clkbuf_1
Xinput10 io_in[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_ls__clkbuf_1
Xinput32 io_in[3] vssd1 vssd1 vccd1 vccd1 AND2X2/B sky130_fd_sc_ls__buf_2
Xinput43 la_data_in[103] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_ls__clkbuf_1
Xinput54 la_data_in[113] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_ls__clkbuf_1
Xinput65 la_data_in[123] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_ls__clkbuf_1
Xinput87 la_data_in[28] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_ls__clkbuf_1
Xinput76 la_data_in[18] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_ls__clkbuf_1
Xinput98 la_data_in[38] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_ls__clkbuf_1
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_420 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1041 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_497 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_105_ vssd1 vssd1 vccd1 vccd1 _105_/HI _105_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_036_ vssd1 vssd1 vccd1 vccd1 _036_/HI _036_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput200 la_oen[14] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_ls__clkbuf_1
Xinput211 la_oen[24] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput222 la_oen[34] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_ls__clkbuf_1
Xinput244 la_oen[54] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_ls__clkbuf_1
Xinput233 la_oen[44] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput288 la_oen[94] vssd1 vssd1 vccd1 vccd1 input288/X sky130_fd_sc_ls__clkbuf_1
Xinput266 la_oen[74] vssd1 vssd1 vccd1 vccd1 input266/X sky130_fd_sc_ls__clkbuf_1
Xinput255 la_oen[64] vssd1 vssd1 vccd1 vccd1 input255/X sky130_fd_sc_ls__clkbuf_1
Xinput277 la_oen[84] vssd1 vssd1 vccd1 vccd1 input277/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput299 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input299/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_261 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_250 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_272 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_294 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_019_ vssd1 vssd1 vccd1 vccd1 _019_/HI _019_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput526 _118_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_ls__clkbuf_2
Xoutput515 _108_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_ls__clkbuf_2
Xoutput504 _098_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_ls__clkbuf_2
Xoutput559 _148_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_ls__clkbuf_2
Xoutput537 _128_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_ls__clkbuf_2
Xoutput548 _138_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_102 _160_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_124 _178_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_113 _069_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_157 _106_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_135 _077_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_146 _087_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_179 _137_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_168 _122_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput8 io_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput378 _004_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_ls__clkbuf_2
Xoutput389 _009_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_827 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_805 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_849 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_198_ vssd1 vssd1 vccd1 vccd1 _198_/HI _198_/LO sky130_fd_sc_ls__conb_1
XFILLER_41_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_13 _022_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_46 _045_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_57 CLKBUF1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_35 _015_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_24 _027_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_68 _051_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_79 AND2X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_21_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_602 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_613 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_646 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_121_ vssd1 vssd1 vccd1 vccd1 _121_/HI _121_/LO sky130_fd_sc_ls__conb_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_052_ vssd1 vssd1 vccd1 vccd1 _052_/HI _052_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput22 io_in[29] vssd1 vssd1 vccd1 vccd1 INVX2/A sky130_fd_sc_ls__clkbuf_4
Xinput11 io_in[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_ls__buf_2
Xinput33 io_in[4] vssd1 vssd1 vccd1 vccd1 AND2X2/A sky130_fd_sc_ls__buf_2
Xinput44 la_data_in[104] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_ls__clkbuf_1
Xinput55 la_data_in[114] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_ls__clkbuf_1
Xinput66 la_data_in[124] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_ls__clkbuf_1
Xinput77 la_data_in[19] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_ls__clkbuf_1
Xinput88 la_data_in[29] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_ls__clkbuf_1
Xinput99 la_data_in[39] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_ls__clkbuf_1
XFILLER_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_410 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_421 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1031 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_104_ vssd1 vssd1 vccd1 vccd1 _104_/HI _104_/LO sky130_fd_sc_ls__conb_1
X_035_ vssd1 vssd1 vccd1 vccd1 _035_/HI _035_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput201 la_oen[15] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_ls__clkbuf_1
Xinput234 la_oen[45] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_ls__clkbuf_1
Xinput223 la_oen[35] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_ls__clkbuf_1
Xinput245 la_oen[55] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_ls__clkbuf_1
Xinput212 la_oen[25] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput278 la_oen[85] vssd1 vssd1 vccd1 vccd1 input278/X sky130_fd_sc_ls__clkbuf_1
Xinput267 la_oen[75] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_ls__clkbuf_1
Xinput256 la_oen[65] vssd1 vssd1 vccd1 vccd1 input256/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput289 la_oen[95] vssd1 vssd1 vccd1 vccd1 input289/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_251 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_262 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_284 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_295 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_018_ vssd1 vssd1 vccd1 vccd1 _018_/HI _018_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput516 _063_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_ls__clkbuf_2
Xoutput527 _064_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_ls__clkbuf_2
Xoutput505 _062_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_ls__clkbuf_2
Xoutput549 _066_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_ls__clkbuf_2
Xoutput538 _065_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_125 _070_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_103 _160_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_114 _069_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_147 _094_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_136 _077_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_158 _106_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_169 _124_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput9 io_in[17] vssd1 vssd1 vccd1 vccd1 BUFX4/A sky130_fd_sc_ls__buf_2
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput368 _012_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_ls__clkbuf_2
Xoutput379 _013_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_817 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_197_ vssd1 vssd1 vccd1 vccd1 _197_/HI _197_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_14 _023_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_25 _027_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_36 _015_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_47 AOI22X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_58 CLKBUF1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_69 INV/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_603 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_636 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_120_ vssd1 vssd1 vccd1 vccd1 _120_/HI _120_/LO sky130_fd_sc_ls__conb_1
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_051_ vssd1 vssd1 vccd1 vccd1 _051_/HI _051_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput12 io_in[1] vssd1 vssd1 vccd1 vccd1 AND2X1/A sky130_fd_sc_ls__buf_2
Xinput34 io_in[5] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_ls__clkbuf_1
Xinput23 io_in[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_ls__clkbuf_1
Xinput45 la_data_in[105] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_ls__clkbuf_1
Xinput67 la_data_in[125] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_ls__clkbuf_1
Xinput78 la_data_in[1] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_ls__clkbuf_1
Xinput89 la_data_in[2] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_ls__clkbuf_1
Xinput56 la_data_in[115] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_ls__clkbuf_1
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_400 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1010 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_455 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_488 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_103_ vssd1 vssd1 vccd1 vccd1 _103_/HI _103_/LO sky130_fd_sc_ls__conb_1
X_034_ vssd1 vssd1 vccd1 vccd1 _034_/HI _034_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput202 la_oen[16] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput235 la_oen[46] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_ls__clkbuf_1
Xinput213 la_oen[26] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_ls__clkbuf_1
Xinput224 la_oen[36] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput257 la_oen[66] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_ls__clkbuf_1
Xinput246 la_oen[56] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_ls__clkbuf_1
Xinput279 la_oen[86] vssd1 vssd1 vccd1 vccd1 input279/X sky130_fd_sc_ls__clkbuf_1
Xinput268 la_oen[76] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_252 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_296 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_017_ vssd1 vssd1 vccd1 vccd1 _017_/HI _017_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput517 _109_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_ls__clkbuf_2
Xoutput506 _099_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput539 _129_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_ls__clkbuf_2
Xoutput528 _119_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XAOI22X1 vccd1 vssd1 AOI22X1/Y input4/X input3/X input5/X input2/X AOI22X1
XFILLER_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_104 _161_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_115 _170_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_137 _079_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_148 _094_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_126 _070_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_159 _107_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput369 _019_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_ls__clkbuf_2
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_818 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_829 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_196_ vssd1 vssd1 vccd1 vccd1 _196_/HI _196_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_15 _023_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_48 AOI22X1/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_37 _017_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_26 _008_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_59 _050_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_604 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_637 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_050_ vssd1 vssd1 vccd1 vccd1 _050_/HI _050_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput13 io_in[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_ls__clkbuf_1
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput24 io_in[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_ls__clkbuf_1
Xinput35 io_in[6] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_ls__clkbuf_2
Xinput46 la_data_in[106] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_ls__clkbuf_1
Xinput68 la_data_in[126] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_ls__clkbuf_1
Xinput57 la_data_in[116] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_ls__clkbuf_1
Xinput79 la_data_in[20] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_ls__clkbuf_1
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_179_ vssd1 vssd1 vccd1 vccd1 _179_/HI _179_/LO sky130_fd_sc_ls__conb_1
XFILLER_42_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_401 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_412 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_1022 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_445 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_478 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_102_ vssd1 vssd1 vccd1 vccd1 _102_/HI _102_/LO sky130_fd_sc_ls__conb_1
X_033_ vssd1 vssd1 vccd1 vccd1 _033_/HI _033_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_990 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput225 la_oen[37] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_ls__clkbuf_1
Xinput236 la_oen[47] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_ls__clkbuf_1
Xinput214 la_oen[27] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_ls__clkbuf_1
Xinput203 la_oen[17] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_ls__clkbuf_1
Xinput269 la_oen[77] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_ls__clkbuf_1
Xinput258 la_oen[67] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_ls__clkbuf_1
Xinput247 la_oen[57] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_242 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_264 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_297 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_016_ vssd1 vssd1 vccd1 vccd1 _016_/HI _016_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput507 _100_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_ls__clkbuf_2
Xoutput518 _110_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_ls__clkbuf_2
Xoutput529 _120_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_105 _161_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_116 _172_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_149 _096_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_138 _079_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_127 _180_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_808 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_819 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_195_ vssd1 vssd1 vccd1 vccd1 _195_/HI _195_/LO sky130_fd_sc_ls__conb_1
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_27 _008_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_38 _017_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_16 _024_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_49 _046_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_605 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput25 io_in[31] vssd1 vssd1 vccd1 vccd1 INVX4/A sky130_fd_sc_ls__clkbuf_4
Xinput14 io_in[21] vssd1 vssd1 vccd1 vccd1 HAX1/B sky130_fd_sc_ls__buf_2
Xinput36 io_in[7] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_ls__buf_2
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput69 la_data_in[127] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_ls__clkbuf_1
Xinput47 la_data_in[107] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_ls__clkbuf_1
Xinput58 la_data_in[117] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_ls__clkbuf_1
X_178_ vssd1 vssd1 vccd1 vccd1 _178_/HI _178_/LO sky130_fd_sc_ls__conb_1
XFILLER_35_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_402 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_424 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_446 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_479 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_101_ vssd1 vssd1 vccd1 vccd1 _101_/HI _101_/LO sky130_fd_sc_ls__conb_1
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_032_ vssd1 vssd1 vccd1 vccd1 _032_/HI _032_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_980 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_991 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput226 la_oen[38] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_ls__clkbuf_1
Xinput215 la_oen[28] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_ls__clkbuf_1
Xinput204 la_oen[18] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput259 la_oen[68] vssd1 vssd1 vccd1 vccd1 input259/X sky130_fd_sc_ls__clkbuf_1
Xinput237 la_oen[48] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_ls__clkbuf_1
Xinput248 la_oen[58] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_210 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_243 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_265 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_276 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_287 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_298 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_015_ vssd1 vssd1 vccd1 vccd1 _015_/HI _015_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput508 _101_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_ls__clkbuf_2
Xoutput519 _111_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_106 _162_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_139 _082_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_128 _183_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_117 _173_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_809 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_194_ vssd1 vssd1 vccd1 vccd1 _194_/HI _194_/LO sky130_fd_sc_ls__conb_1
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_17 _024_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_39 _035_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_28 _220_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_606 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_628 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput26 io_in[32] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_ls__clkbuf_1
Xinput15 io_in[22] vssd1 vssd1 vccd1 vccd1 HAX1/A sky130_fd_sc_ls__buf_2
Xinput37 io_in[8] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_ls__buf_2
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput48 la_data_in[108] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_ls__clkbuf_1
Xinput59 la_data_in[118] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_ls__clkbuf_1
X_177_ vssd1 vssd1 vccd1 vccd1 _177_/HI _177_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_403 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1002 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_436 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_469 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_100_ vssd1 vssd1 vccd1 vccd1 _100_/HI _100_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_031_ vssd1 vssd1 vccd1 vccd1 _031_/HI _031_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_981 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput227 la_oen[39] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_ls__clkbuf_1
Xinput216 la_oen[29] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_ls__clkbuf_1
Xinput205 la_oen[19] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput238 la_oen[49] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_ls__clkbuf_1
Xinput249 la_oen[59] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_ls__clkbuf_1
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_200 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_233 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_266 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_288 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_299 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_014_ vssd1 vssd1 vccd1 vccd1 _014_/HI _014_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput509 _102_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_ls__clkbuf_2
XFILLER_5_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_107 _162_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_118 _173_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_129 _183_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_193_ vssd1 vssd1 vccd1 vccd1 _193_/HI _193_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_29 _220_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_18 _005_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_607 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_618 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput27 io_in[33] vssd1 vssd1 vccd1 vccd1 INVX8/A sky130_fd_sc_ls__clkbuf_4
Xinput16 io_in[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_ls__clkbuf_1
Xinput38 io_in[9] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_ls__clkbuf_1
Xinput49 la_data_in[109] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_ls__clkbuf_1
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_176_ vssd1 vssd1 vccd1 vccd1 _176_/HI _176_/LO sky130_fd_sc_ls__conb_1
XFILLER_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_404 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1003 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1036 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_030_ vssd1 vssd1 vccd1 vccd1 _030_/HI _030_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_971 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_159_ vssd1 vssd1 vccd1 vccd1 _159_/HI _159_/LO sky130_fd_sc_ls__conb_1
XFILLER_40_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput217 la_oen[2] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_ls__clkbuf_1
Xinput206 la_oen[1] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_ls__clkbuf_1
Xinput239 la_oen[4] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_ls__clkbuf_1
Xinput228 la_oen[3] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_201 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_278 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_289 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_013_ vssd1 vssd1 vccd1 vccd1 _013_/HI _013_/LO sky130_fd_sc_ls__conb_1
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_790 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_119 _174_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_108 _164_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_192_ vssd1 vssd1 vccd1 vccd1 _192_/HI _192_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_19 _005_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_70_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_608 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_619 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput28 io_in[34] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_ls__clkbuf_1
Xinput17 io_in[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_ls__clkbuf_1
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_175_ vssd1 vssd1 vccd1 vccd1 _175_/HI _175_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput39 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_ls__clkbuf_1
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XCLKBUF1 vccd1 vssd1 CLKBUF1/Y input11/X CLKBUF1
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_405 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1004 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_1037 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput490 _085_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_ls__clkbuf_2
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_972 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_950 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_994 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_158_ vssd1 vssd1 vccd1 vccd1 _158_/HI _158_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_089_ vssd1 vssd1 vccd1 vccd1 _089_/HI _089_/LO sky130_fd_sc_ls__conb_1
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput207 la_oen[20] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_ls__clkbuf_1
Xinput218 la_oen[30] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_ls__clkbuf_1
Xinput229 la_oen[40] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_ls__clkbuf_1
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_224 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_268 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_279 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
X_012_ vssd1 vssd1 vccd1 vccd1 _012_/HI _012_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_780 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_791 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_109 _167_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_81_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_191_ vssd1 vssd1 vccd1 vccd1 _191_/HI _191_/LO sky130_fd_sc_ls__conb_1
XFILLER_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_609 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput18 io_in[25] vssd1 vssd1 vccd1 vccd1 INV/A sky130_fd_sc_ls__clkbuf_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput29 io_in[35] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_ls__clkbuf_1
X_174_ vssd1 vssd1 vccd1 vccd1 _174_/HI _174_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_406 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_1005 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_439 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput480 _076_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_ls__clkbuf_2
Xoutput491 _086_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_962 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_940 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_995 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_157_ vssd1 vssd1 vccd1 vccd1 _157_/HI _157_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_088_ vssd1 vssd1 vccd1 vccd1 _088_/HI _088_/LO sky130_fd_sc_ls__conb_1
XFILLER_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput208 la_oen[21] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput219 la_oen[31] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_225 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_203 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_269 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_011_ vssd1 vssd1 vccd1 vccd1 _011_/HI _011_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_781 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_209_ vssd1 vssd1 vccd1 vccd1 _209_/HI _209_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_190_ vssd1 vssd1 vccd1 vccd1 _190_/HI _190_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_56_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput19 io_in[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_ls__clkbuf_1
X_173_ vssd1 vssd1 vccd1 vccd1 _173_/HI _173_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_407 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1028 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1006 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1039 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput470 _182_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_ls__clkbuf_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xoutput492 _087_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_ls__clkbuf_2
Xoutput481 _077_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_ls__clkbuf_2
XFILLER_47_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_930 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_70_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_963 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_996 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_974 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_156_ vssd1 vssd1 vccd1 vccd1 _156_/HI _156_/LO sky130_fd_sc_ls__conb_1
X_087_ vssd1 vssd1 vccd1 vccd1 _087_/HI _087_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput209 la_oen[22] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_215 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_204 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_259 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_010_ vssd1 vssd1 vccd1 vccd1 _010_/HI _010_/LO sky130_fd_sc_ls__conb_1
XFILLER_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_771 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_760 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_208_ vssd1 vssd1 vccd1 vccd1 _208_/HI _208_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_139_ vssd1 vssd1 vccd1 vccd1 _139_/HI _139_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_590 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_172_ vssd1 vssd1 vccd1 vccd1 _172_/HI _172_/LO sky130_fd_sc_ls__conb_1
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_408 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_419 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1029 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1007 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput460 _173_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_ls__clkbuf_2
Xoutput471 _183_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_ls__clkbuf_2
Xoutput493 _088_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_ls__clkbuf_2
Xoutput482 _078_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_ls__clkbuf_2
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XAND2X1 vccd1 vssd1 AND2X1/Y AND2X1/A input1/X AND2X1
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_920 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_997 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_155_ vssd1 vssd1 vccd1 vccd1 _155_/HI _155_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_086_ vssd1 vssd1 vccd1 vccd1 _086_/HI _086_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_216 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_205 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_249 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_772 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_750 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_794 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_783 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_207_ vssd1 vssd1 vccd1 vccd1 _207_/HI _207_/LO sky130_fd_sc_ls__conb_1
X_138_ vssd1 vssd1 vccd1 vccd1 _138_/HI _138_/LO sky130_fd_sc_ls__conb_1
X_069_ vssd1 vssd1 vccd1 vccd1 _069_/HI _069_/LO sky130_fd_sc_ls__conb_1
XFILLER_31_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_580 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput360 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input360/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput190 la_oen[120] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_171_ vssd1 vssd1 vccd1 vccd1 _171_/HI _171_/LO sky130_fd_sc_ls__conb_1
XFILLER_22_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_409 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1019 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_1008 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput450 _164_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_ls__clkbuf_2
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput461 _174_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput472 _184_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_ls__clkbuf_2
Xoutput483 _060_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_ls__clkbuf_2
Xoutput494 _061_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XAND2X2 vccd1 vssd1 AND2X2/Y AND2X2/B AND2X2/A AND2X2
XFILLER_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_921 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_910 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_954 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_987 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_998 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_154_ vssd1 vssd1 vccd1 vccd1 _154_/HI _154_/LO sky130_fd_sc_ls__conb_1
X_085_ vssd1 vssd1 vccd1 vccd1 _085_/HI _085_/LO sky130_fd_sc_ls__conb_1
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_206 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_239 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_762 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_740 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_795 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_206_ vssd1 vssd1 vccd1 vccd1 _206_/HI _206_/LO sky130_fd_sc_ls__conb_1
X_137_ vssd1 vssd1 vccd1 vccd1 _137_/HI _137_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_068_ vssd1 vssd1 vccd1 vccd1 _068_/HI _068_/LO sky130_fd_sc_ls__conb_1
XFILLER_24_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_43_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_570 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput350 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 input350/X sky130_fd_sc_ls__clkbuf_1
Xinput361 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input361/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_68_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput180 la_oen[111] vssd1 vssd1 vccd1 vccd1 input180/X sky130_fd_sc_ls__clkbuf_1
Xinput191 la_oen[121] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_170_ vssd1 vssd1 vccd1 vccd1 _170_/HI _170_/LO sky130_fd_sc_ls__conb_1
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_1009 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput440 _039_/LO vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_ls__clkbuf_2
Xoutput451 _165_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_ls__clkbuf_2
Xoutput462 _175_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_ls__clkbuf_2
Xoutput473 _185_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_ls__clkbuf_2
Xoutput495 _089_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_ls__clkbuf_2
Xoutput484 _079_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_ls__clkbuf_2
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_911 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_900 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_944 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_988 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_222_ vssd1 vssd1 vccd1 vccd1 _222_/HI _222_/LO sky130_fd_sc_ls__conb_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_999 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_153_ vssd1 vssd1 vccd1 vccd1 _153_/HI _153_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_084_ vssd1 vssd1 vccd1 vccd1 _084_/HI _084_/LO sky130_fd_sc_ls__conb_1
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_207 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_229 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_763 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_730 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_205_ vssd1 vssd1 vccd1 vccd1 _205_/HI _205_/LO sky130_fd_sc_ls__conb_1
X_136_ vssd1 vssd1 vccd1 vccd1 _136_/HI _136_/LO sky130_fd_sc_ls__conb_1
X_067_ vssd1 vssd1 vccd1 vccd1 _067_/HI _067_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_71_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_560 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_119_ vssd1 vssd1 vccd1 vccd1 _119_/HI _119_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_71_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput351 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 input351/X sky130_fd_sc_ls__clkbuf_1
Xinput362 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 input362/X sky130_fd_sc_ls__clkbuf_1
Xinput340 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 input340/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_390 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XANTENNA_0 _012_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_6_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput181 la_oen[112] vssd1 vssd1 vccd1 vccd1 input181/X sky130_fd_sc_ls__clkbuf_1
Xinput170 la_oen[102] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_ls__clkbuf_1
XFILLER_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput192 la_oen[122] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput600 _193_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_ls__clkbuf_2
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_220 _215_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput430 _054_/LO vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_ls__clkbuf_2
Xoutput441 _040_/LO vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_ls__clkbuf_2
Xoutput452 _166_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_ls__clkbuf_2
Xoutput485 _080_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_ls__clkbuf_2
Xoutput496 _090_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_ls__clkbuf_2
Xoutput463 _176_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_ls__clkbuf_2
Xoutput474 _186_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_912 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_901 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_945 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_923 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_978 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_956 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_221_ vssd1 vssd1 vccd1 vccd1 _221_/HI _221_/LO sky130_fd_sc_ls__conb_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_989 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_152_ vssd1 vssd1 vccd1 vccd1 _152_/HI _152_/LO sky130_fd_sc_ls__conb_1
X_083_ vssd1 vssd1 vccd1 vccd1 _083_/HI _083_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_219 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_208 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_720 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_731 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_786 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_764 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_204_ vssd1 vssd1 vccd1 vccd1 _204_/HI _204_/LO sky130_fd_sc_ls__conb_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_797 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_135_ vssd1 vssd1 vccd1 vccd1 _135_/HI _135_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_066_ vssd1 vssd1 vccd1 vccd1 _066_/HI _066_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_550 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_572 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_118_ vssd1 vssd1 vccd1 vccd1 _118_/HI _118_/LO sky130_fd_sc_ls__conb_1
X_049_ vssd1 vssd1 vccd1 vccd1 _049_/HI _049_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput330 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input330/X sky130_fd_sc_ls__clkbuf_1
Xinput363 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 input363/X sky130_fd_sc_ls__clkbuf_1
Xinput352 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input352/X sky130_fd_sc_ls__clkbuf_1
Xinput341 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input341/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_380 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_391 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XANTENNA_1 _012_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput171 la_oen[103] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_ls__clkbuf_1
Xinput160 la_data_in[94] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput193 la_oen[123] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_ls__clkbuf_1
Xinput182 la_oen[113] vssd1 vssd1 vccd1 vccd1 input182/X sky130_fd_sc_ls__clkbuf_1
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput601 _194_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_221 _190_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_210 _206_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput420 _050_/LO vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_ls__clkbuf_2
Xoutput431 INVX4/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_ls__clkbuf_2
Xoutput442 _041_/LO vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_ls__clkbuf_2
Xoutput453 _167_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_ls__clkbuf_2
Xoutput486 _081_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_ls__clkbuf_2
Xoutput475 _071_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_ls__clkbuf_2
Xoutput464 _177_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_ls__clkbuf_2
Xoutput497 _091_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_902 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_935 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_913 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_220_ vssd1 vssd1 vccd1 vccd1 _220_/HI _220_/LO sky130_fd_sc_ls__conb_1
X_151_ vssd1 vssd1 vccd1 vccd1 _151_/HI _151_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_10_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_082_ vssd1 vssd1 vccd1 vccd1 _082_/HI _082_/LO sky130_fd_sc_ls__conb_1
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_12_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_209 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_47_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_710 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_754 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_203_ vssd1 vssd1 vccd1 vccd1 _203_/HI _203_/LO sky130_fd_sc_ls__conb_1
XPHY_798 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_134_ vssd1 vssd1 vccd1 vccd1 _134_/HI _134_/LO sky130_fd_sc_ls__conb_1
X_065_ vssd1 vssd1 vccd1 vccd1 _065_/HI _065_/LO sky130_fd_sc_ls__conb_1
XFILLER_31_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_540 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_117_ vssd1 vssd1 vccd1 vccd1 _117_/HI _117_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_048_ vssd1 vssd1 vccd1 vccd1 _048_/HI _048_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput320 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 input320/X sky130_fd_sc_ls__clkbuf_1
Xinput353 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 input353/X sky130_fd_sc_ls__clkbuf_1
Xinput342 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 input342/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput331 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 input331/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput364 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 input364/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_370 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_392 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XANTENNA_2 _019_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_62_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_66_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_76_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput172 la_oen[104] vssd1 vssd1 vccd1 vccd1 input172/X sky130_fd_sc_ls__clkbuf_1
Xinput161 la_data_in[95] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_ls__clkbuf_1
Xinput150 la_data_in[85] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_ls__clkbuf_1
Xinput194 la_oen[124] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_ls__clkbuf_1
Xinput183 la_oen[114] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput602 _195_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_ls__clkbuf_2
XFILLER_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XANTENNA_200 _155_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_222 _190_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_211 _189_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput410 _045_/LO vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_ls__clkbuf_2
Xoutput432 _055_/LO vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_ls__clkbuf_2
Xoutput421 HAX1/YS vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_ls__clkbuf_2
Xoutput443 AOI21X1/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_ls__clkbuf_2
Xoutput454 _168_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_ls__clkbuf_2
Xoutput476 _072_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_ls__clkbuf_2
Xoutput487 _082_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_ls__clkbuf_2
Xoutput465 _178_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_ls__clkbuf_2
Xoutput498 _092_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_ls__clkbuf_2
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_903 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_936 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_914 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_150_ vssd1 vssd1 vccd1 vccd1 _150_/HI _150_/LO sky130_fd_sc_ls__conb_1
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
X_081_ vssd1 vssd1 vccd1 vccd1 _081_/HI _081_/LO sky130_fd_sc_ls__conb_1
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_28_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_700 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_755 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_202_ vssd1 vssd1 vccd1 vccd1 _202_/HI _202_/LO sky130_fd_sc_ls__conb_1
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_799 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_133_ vssd1 vssd1 vccd1 vccd1 _133_/HI _133_/LO sky130_fd_sc_ls__conb_1
X_064_ vssd1 vssd1 vccd1 vccd1 _064_/HI _064_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_25_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_541 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_116_ vssd1 vssd1 vccd1 vccd1 _116_/HI _116_/LO sky130_fd_sc_ls__conb_1
X_047_ vssd1 vssd1 vccd1 vccd1 _047_/HI _047_/LO sky130_fd_sc_ls__conb_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xinput321 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 input321/X sky130_fd_sc_ls__clkbuf_1
Xinput310 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 input310/X sky130_fd_sc_ls__clkbuf_1
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput354 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 input354/X sky130_fd_sc_ls__clkbuf_1
Xinput343 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 input343/X sky130_fd_sc_ls__clkbuf_1
Xinput332 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 input332/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
Xinput365 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 input365/X sky130_fd_sc_ls__clkbuf_1
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_360 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_371 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_3 _019_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_72_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_9_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput140 la_data_in[76] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_ls__clkbuf_1
Xinput151 la_data_in[86] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_ls__clkbuf_1
Xinput162 la_data_in[96] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_ls__clkbuf_1
Xinput184 la_oen[115] vssd1 vssd1 vccd1 vccd1 input184/X sky130_fd_sc_ls__clkbuf_1
Xinput173 la_oen[105] vssd1 vssd1 vccd1 vccd1 input173/X sky130_fd_sc_ls__clkbuf_1
Xinput195 la_oen[125] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_190 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput603 _196_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_ls__clkbuf_2
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_223 _218_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_212 _189_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XANTENNA_201 _068_/LO vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
XFILLER_26_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_13_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput400 _015_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_ls__clkbuf_2
Xoutput411 AOI22X1/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_ls__clkbuf_2
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
Xoutput433 INVX8/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_ls__clkbuf_2
Xoutput422 HAX1/YC vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_ls__clkbuf_2
Xoutput444 _059_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_ls__clkbuf_2
Xoutput466 _070_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_ls__clkbuf_2
Xoutput477 _073_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_ls__clkbuf_2
Xoutput455 _069_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_ls__clkbuf_2
XFILLER_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xoutput499 _093_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_ls__clkbuf_2
Xoutput488 _083_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_ls__clkbuf_2
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_926 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_904 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_959 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_080_ vssd1 vssd1 vccd1 vccd1 _080_/HI _080_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_2_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_45_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_68_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XPHY_701 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_712 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_201_ vssd1 vssd1 vccd1 vccd1 _201_/HI _201_/LO sky130_fd_sc_ls__conb_1
XFILLER_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_778 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_756 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XPHY_789 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
X_132_ vssd1 vssd1 vccd1 vccd1 _132_/HI _132_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_063_ vssd1 vssd1 vccd1 vccd1 _063_/HI _063_/LO sky130_fd_sc_ls__conb_1
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_78_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_73_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_520 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_34_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_564 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_597 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
X_115_ vssd1 vssd1 vccd1 vccd1 _115_/HI _115_/LO sky130_fd_sc_ls__conb_1
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
X_046_ vssd1 vssd1 vccd1 vccd1 _046_/HI _046_/LO sky130_fd_sc_ls__conb_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_55_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
Xinput311 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 input311/X sky130_fd_sc_ls__clkbuf_1
Xinput300 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input300/X sky130_fd_sc_ls__clkbuf_1
Xinput344 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 input344/X sky130_fd_sc_ls__clkbuf_1
Xinput322 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 input322/X sky130_fd_sc_ls__clkbuf_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput333 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 input333/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput366 wbs_stb_i vssd1 vssd1 vccd1 vccd1 input366/X sky130_fd_sc_ls__clkbuf_1
Xinput355 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input355/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_350 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_372 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_8_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XANTENNA_4 _020_/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__diode_2
X_029_ vssd1 vssd1 vccd1 vccd1 _029_/HI _029_/LO sky130_fd_sc_ls__conb_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_30_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XHAX1 vccd1 vssd1 HAX1/YS HAX1/YC HAX1/B HAX1/A HAX1
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_5_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput163 la_data_in[97] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_ls__clkbuf_1
Xinput152 la_data_in[87] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_ls__clkbuf_1
Xinput130 la_data_in[67] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_ls__clkbuf_1
Xinput141 la_data_in[77] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_ls__clkbuf_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xinput185 la_oen[116] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_ls__clkbuf_1
Xinput196 la_oen[126] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_ls__clkbuf_1
Xinput174 la_oen[106] vssd1 vssd1 vccd1 vccd1 input174/X sky130_fd_sc_ls__clkbuf_1
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_1
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__fill_diode_2
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XPHY_191 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XPHY_180 vssd1 vccd1 sky130_fd_sc_ls__tapvpwrvgnd_1
XFILLER_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
XFILLER_75_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_8
Xoutput604 _197_/LO vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_ls__clkbuf_2
XFILLER_4_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_ls__decap_4
.ends

