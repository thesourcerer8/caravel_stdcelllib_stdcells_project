VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 3.220 3.010 3.510 3.090 ;
        RECT 3.220 2.840 3.280 3.010 ;
        RECT 3.450 2.840 3.510 3.010 ;
        RECT 3.220 2.780 3.510 2.840 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 0.490 0.870 0.550 ;
        RECT 0.580 0.320 0.640 0.490 ;
        RECT 0.810 0.320 0.870 0.490 ;
        RECT 0.580 0.240 0.870 0.320 ;
        RECT 3.220 0.490 3.510 0.550 ;
        RECT 3.220 0.320 3.280 0.490 ;
        RECT 3.450 0.320 3.510 0.490 ;
        RECT 3.220 0.240 3.510 0.320 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.200 4.950 2.490 ;
        RECT 4.730 0.730 4.870 2.200 ;
        RECT 4.660 0.440 4.950 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.540 1.510 1.780 ;
        RECT 1.300 1.250 1.590 1.540 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 2.810 1.540 2.950 1.780 ;
        RECT 2.740 1.250 3.030 1.540 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 3.200 3.010 3.530 3.090 ;
        RECT 3.200 2.840 3.280 3.010 ;
        RECT 3.450 2.840 3.530 3.010 ;
        RECT 3.200 2.760 3.530 2.840 ;
        RECT 0.800 2.430 1.130 2.510 ;
        RECT 0.800 2.260 0.880 2.430 ;
        RECT 1.050 2.260 1.130 2.430 ;
        RECT 4.640 2.430 4.970 2.510 ;
        RECT 4.640 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.970 2.430 ;
        RECT 0.800 2.180 1.110 2.260 ;
        RECT 4.660 2.180 4.970 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 1.360 1.160 1.530 1.310 ;
        RECT 2.800 1.160 2.970 1.310 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.920 2.800 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.740 0.910 2.800 0.920 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.740 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 2.240 0.670 2.570 0.750 ;
        RECT 0.560 0.490 0.890 0.570 ;
        RECT 0.560 0.320 0.640 0.490 ;
        RECT 0.810 0.320 0.890 0.490 ;
        RECT 2.240 0.500 2.320 0.670 ;
        RECT 2.490 0.500 2.570 0.670 ;
        RECT 4.660 0.670 4.970 0.750 ;
        RECT 4.660 0.660 4.720 0.670 ;
        RECT 2.240 0.420 2.570 0.500 ;
        RECT 3.200 0.490 3.530 0.570 ;
        RECT 0.560 0.240 0.890 0.320 ;
        RECT 3.200 0.320 3.280 0.490 ;
        RECT 3.450 0.320 3.530 0.490 ;
        RECT 4.640 0.500 4.720 0.660 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
        RECT 3.200 0.240 3.530 0.320 ;
      LAYER met1 ;
        RECT 0.820 2.430 1.110 2.490 ;
        RECT 0.820 2.260 0.880 2.430 ;
        RECT 1.050 2.260 1.110 2.430 ;
        RECT 0.820 2.200 1.110 2.260 ;
        RECT 0.890 1.060 1.030 2.200 ;
        RECT 4.180 2.010 4.470 2.070 ;
        RECT 4.180 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.470 2.010 ;
        RECT 4.180 1.780 4.470 1.840 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 4.180 1.080 4.470 1.140 ;
        RECT 4.180 1.060 4.240 1.080 ;
        RECT 0.890 0.920 4.240 1.060 ;
        RECT 2.330 0.730 2.470 0.920 ;
        RECT 4.180 0.910 4.240 0.920 ;
        RECT 4.410 0.910 4.470 1.080 ;
        RECT 4.180 0.850 4.470 0.910 ;
        RECT 2.260 0.670 2.550 0.730 ;
        RECT 2.260 0.500 2.320 0.670 ;
        RECT 2.490 0.500 2.550 0.670 ;
        RECT 2.260 0.440 2.550 0.500 ;
  END
END OR2X1
END LIBRARY

