magic
tech sky130A
timestamp 1623602949
<< nwell >>
rect 0 179 1584 333
<< nmos >>
rect 137 24 152 66
rect 425 24 440 66
rect 569 24 584 66
rect 857 24 872 66
rect 1001 24 1016 66
rect 1145 24 1160 66
rect 1433 24 1448 66
<< pmos >>
rect 137 225 152 309
rect 425 225 440 309
rect 569 225 584 309
rect 857 225 872 309
rect 1001 225 1016 309
rect 1145 225 1160 309
rect 1433 225 1448 309
<< ndiff >>
rect 58 66 87 69
rect 346 66 375 69
rect 1042 66 1071 69
rect 1474 66 1503 69
rect 58 63 137 66
rect 58 46 64 63
rect 81 46 137 63
rect 58 24 137 46
rect 152 36 231 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 231 36
rect 346 63 425 66
rect 346 46 352 63
rect 369 46 425 63
rect 346 24 425 46
rect 440 24 569 66
rect 584 36 663 66
rect 584 24 616 36
rect 201 19 207 24
rect 178 13 207 19
rect 610 19 616 24
rect 633 24 663 36
rect 778 36 857 66
rect 633 19 639 24
rect 610 13 639 19
rect 778 19 784 36
rect 801 24 857 36
rect 872 36 1001 66
rect 872 24 952 36
rect 801 19 807 24
rect 778 13 807 19
rect 946 19 952 24
rect 969 24 1001 36
rect 1016 63 1145 66
rect 1016 46 1048 63
rect 1065 46 1145 63
rect 1016 24 1145 46
rect 1160 36 1239 66
rect 1160 24 1192 36
rect 969 19 975 24
rect 946 13 975 19
rect 1186 19 1192 24
rect 1209 24 1239 36
rect 1354 36 1433 66
rect 1209 19 1215 24
rect 1186 13 1215 19
rect 1354 19 1360 36
rect 1377 24 1433 36
rect 1448 63 1527 66
rect 1448 46 1480 63
rect 1497 46 1527 63
rect 1448 24 1527 46
rect 1377 19 1383 24
rect 1354 13 1383 19
<< pdiff >>
rect 178 309 207 312
rect 466 309 495 312
rect 778 309 807 312
rect 1186 309 1215 312
rect 1354 309 1383 312
rect 58 238 137 309
rect 58 221 64 238
rect 81 225 137 238
rect 152 306 231 309
rect 152 289 184 306
rect 201 289 231 306
rect 152 225 231 289
rect 346 238 425 309
rect 81 221 87 225
rect 58 215 87 221
rect 346 221 352 238
rect 369 225 425 238
rect 440 306 569 309
rect 440 289 472 306
rect 489 289 569 306
rect 440 225 569 289
rect 584 238 663 309
rect 584 225 616 238
rect 369 221 375 225
rect 346 215 375 221
rect 610 221 616 225
rect 633 225 663 238
rect 778 306 857 309
rect 778 289 784 306
rect 801 289 857 306
rect 778 225 857 289
rect 872 238 1001 309
rect 872 225 952 238
rect 633 221 639 225
rect 610 215 639 221
rect 946 221 952 225
rect 969 225 1001 238
rect 1016 225 1145 309
rect 1160 306 1239 309
rect 1160 289 1192 306
rect 1209 289 1239 306
rect 1160 225 1239 289
rect 1354 306 1433 309
rect 1354 289 1360 306
rect 1377 289 1433 306
rect 1354 225 1433 289
rect 1448 238 1527 309
rect 1448 225 1480 238
rect 969 221 975 225
rect 946 215 975 221
rect 1474 221 1480 225
rect 1497 225 1527 238
rect 1497 221 1503 225
rect 1474 215 1503 221
<< ndiffc >>
rect 64 46 81 63
rect 184 19 201 36
rect 352 46 369 63
rect 616 19 633 36
rect 784 19 801 36
rect 952 19 969 36
rect 1048 46 1065 63
rect 1192 19 1209 36
rect 1360 19 1377 36
rect 1480 46 1497 63
<< pdiffc >>
rect 64 221 81 238
rect 184 289 201 306
rect 352 221 369 238
rect 472 289 489 306
rect 616 221 633 238
rect 784 289 801 306
rect 952 221 969 238
rect 1192 289 1209 306
rect 1360 289 1377 306
rect 1480 221 1497 238
<< poly >>
rect 137 309 152 330
rect 425 309 440 330
rect 569 309 584 330
rect 857 309 872 330
rect 1001 309 1016 330
rect 1145 309 1160 330
rect 1433 309 1448 330
rect 137 206 152 225
rect 425 206 440 225
rect 569 206 584 225
rect 857 206 872 225
rect 1001 206 1016 225
rect 1145 206 1160 225
rect 1433 206 1448 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 848 198 881 206
rect 848 181 856 198
rect 873 181 881 198
rect 848 173 881 181
rect 992 198 1025 206
rect 992 181 1000 198
rect 1017 181 1025 198
rect 992 173 1025 181
rect 1136 198 1169 206
rect 1136 181 1144 198
rect 1161 181 1169 198
rect 1136 173 1169 181
rect 1424 198 1457 206
rect 1424 181 1432 198
rect 1449 181 1457 198
rect 1424 173 1457 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 848 103 881 111
rect 848 86 856 103
rect 873 86 881 103
rect 848 78 881 86
rect 992 103 1025 111
rect 992 86 1000 103
rect 1017 86 1025 103
rect 992 78 1025 86
rect 1136 103 1169 111
rect 1136 86 1144 103
rect 1161 86 1169 103
rect 1136 78 1169 86
rect 1424 103 1457 111
rect 1424 86 1432 103
rect 1449 86 1457 103
rect 1424 78 1457 86
rect 137 66 152 78
rect 425 66 440 78
rect 569 66 584 78
rect 857 66 872 78
rect 1001 66 1016 78
rect 1145 66 1160 78
rect 1433 66 1448 78
rect 137 11 152 24
rect 425 11 440 24
rect 569 11 584 24
rect 857 11 872 24
rect 1001 11 1016 24
rect 1145 11 1160 24
rect 1433 11 1448 24
<< polycont >>
rect 136 181 153 198
rect 424 181 441 198
rect 568 181 585 198
rect 856 181 873 198
rect 1000 181 1017 198
rect 1144 181 1161 198
rect 1432 181 1449 198
rect 136 86 153 103
rect 424 86 441 103
rect 568 86 585 103
rect 856 86 873 103
rect 1000 86 1017 103
rect 1144 86 1161 103
rect 1432 86 1449 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 464 306 497 314
rect 464 289 472 306
rect 489 289 497 306
rect 464 281 497 289
rect 776 289 784 314
rect 801 289 809 314
rect 776 281 809 289
rect 1184 306 1217 314
rect 1184 289 1192 306
rect 1209 289 1217 306
rect 1184 281 1217 289
rect 1352 306 1385 314
rect 1352 289 1360 306
rect 1377 289 1385 306
rect 1352 281 1385 289
rect 56 238 89 246
rect 56 221 64 238
rect 81 221 89 238
rect 56 213 89 221
rect 344 238 377 246
rect 344 221 352 238
rect 369 221 377 238
rect 344 213 377 221
rect 568 206 585 262
rect 608 238 641 246
rect 608 221 616 238
rect 633 221 641 238
rect 608 213 641 221
rect 944 238 977 246
rect 944 221 952 238
rect 969 223 977 238
rect 1472 238 1505 246
rect 1472 223 1480 238
rect 969 221 975 223
rect 944 213 975 221
rect 1474 221 1480 223
rect 1497 221 1505 238
rect 1474 213 1505 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 591 206
rect 560 181 568 198
rect 585 196 591 198
rect 848 198 881 206
rect 585 181 593 196
rect 560 173 593 181
rect 848 181 856 198
rect 873 181 881 198
rect 848 173 881 181
rect 992 198 1025 206
rect 992 181 1000 198
rect 1017 181 1025 198
rect 992 173 1025 181
rect 1136 198 1169 206
rect 1136 181 1144 198
rect 1161 181 1169 198
rect 1136 173 1169 181
rect 1424 198 1457 206
rect 1424 181 1432 198
rect 1449 181 1457 198
rect 1424 173 1457 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 848 103 881 111
rect 848 86 856 103
rect 873 86 881 103
rect 848 78 881 86
rect 992 103 1025 111
rect 992 86 1000 103
rect 1017 86 1025 103
rect 992 78 1025 86
rect 1136 103 1169 111
rect 1136 86 1144 103
rect 1161 86 1169 103
rect 1136 78 1169 86
rect 1424 103 1457 111
rect 1424 86 1432 103
rect 1449 88 1457 103
rect 1449 86 1455 88
rect 1424 78 1455 86
rect 56 63 89 71
rect 56 46 64 63
rect 81 46 89 63
rect 56 38 89 46
rect 344 63 377 71
rect 344 46 352 63
rect 369 46 377 63
rect 1042 63 1073 71
rect 1042 61 1048 63
rect 176 36 209 44
rect 344 38 377 46
rect 1040 46 1048 61
rect 1065 46 1073 63
rect 176 19 184 36
rect 201 19 209 36
rect 176 11 209 19
rect 608 36 641 44
rect 608 11 616 36
rect 633 11 641 36
rect 776 36 809 44
rect 776 11 784 36
rect 801 11 809 36
rect 944 36 977 44
rect 1040 39 1073 46
rect 1472 63 1505 71
rect 1472 46 1480 63
rect 1497 46 1505 63
rect 944 19 952 36
rect 969 22 977 36
rect 1184 36 1217 44
rect 1184 22 1192 36
rect 969 19 1192 22
rect 1209 19 1217 36
rect 944 11 1217 19
rect 1352 36 1385 44
rect 1472 38 1505 46
rect 1352 11 1360 36
rect 952 5 1209 11
rect 1377 11 1385 36
<< viali >>
rect 184 289 201 306
rect 472 289 489 306
rect 784 306 801 319
rect 784 302 801 306
rect 1192 289 1209 306
rect 1360 289 1377 306
rect 568 262 585 279
rect 64 221 81 238
rect 352 221 369 238
rect 616 221 633 238
rect 952 221 969 238
rect 1480 221 1497 238
rect 136 181 153 198
rect 424 181 441 198
rect 568 181 585 198
rect 856 181 873 198
rect 1000 181 1017 198
rect 1144 181 1161 198
rect 1432 181 1449 198
rect 136 86 153 103
rect 424 86 441 103
rect 568 86 585 103
rect 856 86 873 103
rect 1000 86 1017 103
rect 1144 86 1161 103
rect 1432 86 1449 103
rect 64 46 81 63
rect 352 46 369 63
rect 1048 46 1065 63
rect 184 19 201 36
rect 616 19 633 22
rect 616 5 633 19
rect 784 19 801 22
rect 784 5 801 19
rect 1480 46 1497 63
rect 1360 19 1377 22
rect 1360 5 1377 19
<< metal1 >>
rect 0 319 1584 357
rect 0 309 784 319
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 466 306 495 309
rect 466 289 472 306
rect 489 289 495 306
rect 778 302 784 309
rect 801 309 1584 319
rect 801 302 807 309
rect 778 296 807 302
rect 1186 306 1215 309
rect 466 283 495 289
rect 1186 289 1192 306
rect 1209 289 1215 306
rect 562 279 591 285
rect 1186 283 1215 289
rect 1354 306 1383 309
rect 1354 289 1360 306
rect 1377 289 1383 306
rect 1354 283 1383 289
rect 562 262 568 279
rect 585 277 591 279
rect 585 263 1159 277
rect 585 262 591 263
rect 562 256 591 262
rect 58 238 87 244
rect 58 221 64 238
rect 81 221 87 238
rect 58 215 87 221
rect 346 238 375 244
rect 346 221 352 238
rect 369 237 375 238
rect 610 238 639 244
rect 610 237 616 238
rect 369 223 616 237
rect 369 221 375 223
rect 346 215 375 221
rect 610 221 616 223
rect 633 237 639 238
rect 946 238 975 244
rect 633 223 871 237
rect 633 221 639 223
rect 610 215 639 221
rect 65 69 79 215
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 137 109 151 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 102 159 103
rect 353 102 367 215
rect 857 204 871 223
rect 946 221 952 238
rect 969 237 975 238
rect 969 223 1063 237
rect 969 221 975 223
rect 946 215 975 221
rect 418 198 447 204
rect 418 181 424 198
rect 441 181 447 198
rect 418 175 447 181
rect 562 198 591 204
rect 562 181 568 198
rect 585 181 591 198
rect 562 175 591 181
rect 850 198 879 204
rect 850 181 856 198
rect 873 181 879 198
rect 850 175 879 181
rect 994 198 1023 204
rect 994 181 1000 198
rect 1017 181 1023 198
rect 994 175 1023 181
rect 425 109 439 175
rect 569 109 583 175
rect 857 109 871 175
rect 1001 109 1015 175
rect 153 88 367 102
rect 153 86 159 88
rect 130 80 159 86
rect 353 69 367 88
rect 418 103 447 109
rect 418 86 424 103
rect 441 86 447 103
rect 418 80 447 86
rect 562 103 591 109
rect 562 86 568 103
rect 585 86 591 103
rect 562 80 591 86
rect 850 103 879 109
rect 850 86 856 103
rect 873 86 879 103
rect 850 80 879 86
rect 994 103 1023 109
rect 994 86 1000 103
rect 1017 86 1023 103
rect 994 80 1023 86
rect 58 63 87 69
rect 58 46 64 63
rect 81 46 87 63
rect 58 40 87 46
rect 346 63 375 69
rect 346 46 352 63
rect 369 46 375 63
rect 425 61 439 80
rect 1001 61 1015 80
rect 1049 69 1063 223
rect 1145 204 1159 263
rect 1474 238 1503 244
rect 1474 221 1480 238
rect 1497 221 1503 238
rect 1474 215 1503 221
rect 1138 198 1167 204
rect 1138 181 1144 198
rect 1161 181 1167 198
rect 1138 175 1167 181
rect 1426 198 1455 204
rect 1426 181 1432 198
rect 1449 181 1455 198
rect 1426 175 1455 181
rect 1145 109 1159 175
rect 1433 109 1447 175
rect 1138 103 1167 109
rect 1138 86 1144 103
rect 1161 86 1167 103
rect 1138 80 1167 86
rect 1426 103 1455 109
rect 1426 86 1432 103
rect 1449 86 1455 103
rect 1426 80 1455 86
rect 425 47 1015 61
rect 1042 63 1071 69
rect 178 36 207 42
rect 346 40 375 46
rect 1042 46 1048 63
rect 1065 61 1071 63
rect 1433 61 1447 80
rect 1481 69 1495 215
rect 1065 47 1447 61
rect 1474 63 1503 69
rect 1065 46 1071 47
rect 1042 40 1071 46
rect 1474 46 1480 63
rect 1497 46 1503 63
rect 1474 40 1503 46
rect 178 24 184 36
rect 0 19 184 24
rect 201 24 207 36
rect 610 24 639 28
rect 778 24 807 28
rect 1354 24 1383 28
rect 201 22 1584 24
rect 201 19 616 22
rect 0 5 616 19
rect 633 5 784 22
rect 801 5 1360 22
rect 1377 5 1584 22
rect 0 -24 1584 5
<< labels >>
rlabel metal1 0 309 1584 357 0 VDD
port 1 se
rlabel metal1 0 -24 1584 24 0 GND
port 2 se
rlabel metal1 1474 40 1503 69 0 YS
port 3 se
rlabel metal1 1481 69 1495 215 0 YS
port 4 se
rlabel metal1 1474 215 1503 244 0 YS
port 5 se
rlabel metal1 58 40 87 69 0 YC
port 6 se
rlabel metal1 65 69 79 215 0 YC
port 7 se
rlabel metal1 58 215 87 244 0 YC
port 8 se
rlabel metal1 562 80 591 109 0 A
port 9 se
rlabel metal1 569 109 583 175 0 A
port 10 se
rlabel metal1 562 175 591 204 0 A
port 11 se
rlabel metal1 425 47 1015 61 0 B
port 12 se
rlabel metal1 425 61 439 80 0 B
port 13 se
rlabel metal1 1001 61 1015 80 0 B
port 14 se
rlabel metal1 418 80 447 109 0 B
port 15 se
rlabel metal1 994 80 1023 109 0 B
port 16 se
rlabel metal1 425 109 439 175 0 B
port 17 se
rlabel metal1 1001 109 1015 175 0 B
port 18 se
rlabel metal1 418 175 447 204 0 B
port 19 se
rlabel metal1 994 175 1023 204 0 B
port 20 se
<< properties >>
string FIXED_BBOX 0 0 1584 333
<< end >>
