magic
tech sky130A
timestamp 1621277091
<< end >>
