VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 2.880 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.880 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.150 0.870 2.440 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 2.810 2.090 3.140 ;
        RECT 0.560 2.130 0.890 2.460 ;
        RECT 1.280 1.730 1.610 2.060 ;
        RECT 1.280 0.780 1.610 1.110 ;
        RECT 0.560 0.380 0.890 0.710 ;
        RECT 1.760 0.110 2.090 0.440 ;
  END
END INVX2
END LIBRARY

