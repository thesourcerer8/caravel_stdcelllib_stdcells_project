MACRO AND2X1
 CLASS CORE ;
 FOREIGN AND2X1 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 4.65500000 0.39500000 4.94500000 0.68500000 ;
        RECT 4.73000000 0.68500000 4.87000000 2.15000000 ;
        RECT 4.65500000 2.15000000 4.94500000 2.44000000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.73500000 0.80000000 3.02500000 1.09000000 ;
        RECT 2.81000000 1.09000000 2.95000000 1.74500000 ;
        RECT 2.73500000 1.74500000 3.02500000 2.03500000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.29500000 0.80000000 1.58500000 1.09000000 ;
        RECT 1.37000000 1.09000000 1.51000000 1.74500000 ;
        RECT 1.29500000 1.74500000 1.58500000 2.03500000 ;
    END
  END A


END AND2X1
