VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SUTHERLAND1989
  CLASS CORE ;
  FOREIGN SUTHERLAND1989 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 3.220 2.970 3.510 3.090 ;
        RECT 3.220 2.800 3.280 2.970 ;
        RECT 3.450 2.800 3.510 2.970 ;
        RECT 3.220 2.740 3.510 2.800 ;
        RECT 6.100 2.970 6.390 3.090 ;
        RECT 6.100 2.800 6.160 2.970 ;
        RECT 6.330 2.800 6.390 2.970 ;
        RECT 6.100 2.740 6.390 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 3.200 2.970 3.530 3.090 ;
        RECT 3.200 2.800 3.280 2.970 ;
        RECT 3.450 2.800 3.530 2.970 ;
        RECT 3.200 2.720 3.530 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.220 0.670 3.510 0.730 ;
        RECT 3.220 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.510 0.670 ;
        RECT 3.220 0.440 3.510 0.500 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.080 0.670 6.410 0.750 ;
        RECT 6.080 0.500 6.160 0.670 ;
        RECT 6.330 0.500 6.410 0.670 ;
        RECT 6.080 0.420 6.410 0.500 ;
        RECT 6.160 0.240 6.330 0.420 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
  END VGND
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.780 1.060 8.070 1.140 ;
        RECT 9.940 1.060 10.230 1.140 ;
        RECT 7.780 0.920 10.230 1.060 ;
        RECT 7.780 0.850 8.070 0.920 ;
        RECT 9.940 0.850 10.230 0.920 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 2.000 1.590 2.070 ;
        RECT 5.620 2.000 5.910 2.070 ;
        RECT 1.300 1.860 5.910 2.000 ;
        RECT 1.300 1.780 1.590 1.860 ;
        RECT 5.620 1.780 5.910 1.860 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 5.690 1.140 5.830 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
        RECT 5.620 0.850 5.910 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.060 3.030 1.140 ;
        RECT 4.180 1.060 4.470 1.140 ;
        RECT 2.740 0.920 4.470 1.060 ;
        RECT 2.740 0.850 3.030 0.920 ;
        RECT 4.180 0.850 4.470 0.920 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 6.080 2.970 6.410 3.050 ;
        RECT 6.080 2.800 6.160 2.970 ;
        RECT 6.330 2.800 6.410 2.970 ;
        RECT 6.080 2.720 6.410 2.800 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 5.120 2.430 5.450 2.510 ;
        RECT 5.120 2.260 5.200 2.430 ;
        RECT 5.370 2.260 5.450 2.430 ;
        RECT 7.760 2.430 8.090 2.510 ;
        RECT 7.760 2.260 7.840 2.430 ;
        RECT 8.010 2.260 8.090 2.430 ;
        RECT 5.120 2.180 5.430 2.260 ;
        RECT 7.760 2.180 8.090 2.260 ;
        RECT 9.200 2.430 9.530 2.510 ;
        RECT 9.200 2.260 9.280 2.430 ;
        RECT 9.450 2.260 9.530 2.430 ;
        RECT 10.400 2.430 10.730 2.510 ;
        RECT 10.400 2.260 10.480 2.430 ;
        RECT 10.650 2.260 10.730 2.430 ;
        RECT 9.200 2.180 9.530 2.260 ;
        RECT 10.420 2.180 10.730 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 2.800 1.160 2.970 1.760 ;
        RECT 4.240 1.160 4.410 1.760 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.920 3.050 1.080 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 2.970 0.910 3.030 0.920 ;
        RECT 2.720 0.830 3.030 0.910 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.920 5.930 1.080 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.840 1.080 8.010 2.180 ;
        RECT 9.920 2.010 10.250 2.090 ;
        RECT 9.920 1.840 10.000 2.010 ;
        RECT 10.170 1.840 10.250 2.010 ;
        RECT 9.920 1.760 10.250 1.840 ;
        RECT 10.000 1.160 10.170 1.760 ;
        RECT 9.920 1.080 10.250 1.160 ;
        RECT 5.850 0.910 5.910 0.920 ;
        RECT 5.600 0.830 5.910 0.910 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.370 1.080 ;
        RECT 9.920 0.910 10.000 1.080 ;
        RECT 10.170 0.910 10.250 1.080 ;
        RECT 7.040 0.830 7.370 0.910 ;
        RECT 7.840 0.750 8.010 0.910 ;
        RECT 9.920 0.830 10.250 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 3.200 0.670 3.530 0.750 ;
        RECT 3.200 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
        RECT 5.120 0.670 5.430 0.750 ;
        RECT 5.120 0.500 5.200 0.670 ;
        RECT 5.370 0.660 5.430 0.670 ;
        RECT 7.760 0.670 8.090 0.750 ;
        RECT 5.370 0.500 5.450 0.660 ;
        RECT 5.120 0.420 5.450 0.500 ;
        RECT 7.760 0.500 7.840 0.670 ;
        RECT 8.010 0.500 8.090 0.670 ;
        RECT 7.760 0.420 8.090 0.500 ;
        RECT 9.200 0.670 9.530 0.750 ;
        RECT 9.200 0.500 9.280 0.670 ;
        RECT 9.450 0.500 9.530 0.670 ;
        RECT 10.420 0.670 10.730 0.750 ;
        RECT 10.420 0.660 10.480 0.670 ;
        RECT 9.200 0.420 9.530 0.500 ;
        RECT 10.400 0.500 10.480 0.660 ;
        RECT 10.650 0.500 10.730 0.670 ;
        RECT 10.400 0.420 10.730 0.500 ;
      LAYER met1 ;
        RECT 0.580 2.430 0.870 2.490 ;
        RECT 0.580 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.870 2.430 ;
        RECT 0.580 2.200 0.870 2.260 ;
        RECT 5.140 2.430 5.430 2.490 ;
        RECT 5.140 2.260 5.200 2.430 ;
        RECT 5.370 2.410 5.430 2.430 ;
        RECT 9.220 2.430 9.510 2.490 ;
        RECT 9.220 2.410 9.280 2.430 ;
        RECT 5.370 2.270 9.280 2.410 ;
        RECT 5.370 2.260 5.430 2.270 ;
        RECT 5.140 2.200 5.430 2.260 ;
        RECT 9.220 2.260 9.280 2.270 ;
        RECT 9.450 2.260 9.510 2.430 ;
        RECT 9.220 2.200 9.510 2.260 ;
        RECT 10.420 2.430 10.710 2.490 ;
        RECT 10.420 2.260 10.480 2.430 ;
        RECT 10.650 2.260 10.710 2.430 ;
        RECT 10.420 2.200 10.710 2.260 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 7.060 2.010 7.350 2.070 ;
        RECT 7.060 1.840 7.120 2.010 ;
        RECT 7.290 2.000 7.350 2.010 ;
        RECT 10.490 2.000 10.630 2.200 ;
        RECT 7.290 1.860 10.630 2.000 ;
        RECT 7.290 1.840 7.350 1.860 ;
        RECT 7.060 1.780 7.350 1.840 ;
        RECT 7.130 1.140 7.270 1.780 ;
        RECT 7.060 1.080 7.350 1.140 ;
        RECT 7.060 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.350 1.080 ;
        RECT 7.060 0.850 7.350 0.910 ;
        RECT 10.490 0.730 10.630 1.860 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 5.140 0.670 5.430 0.730 ;
        RECT 5.140 0.500 5.200 0.670 ;
        RECT 5.370 0.660 5.430 0.670 ;
        RECT 9.220 0.670 9.510 0.730 ;
        RECT 9.220 0.660 9.280 0.670 ;
        RECT 5.370 0.520 9.280 0.660 ;
        RECT 5.370 0.500 5.430 0.520 ;
        RECT 5.140 0.440 5.430 0.500 ;
        RECT 9.220 0.500 9.280 0.520 ;
        RECT 9.450 0.500 9.510 0.670 ;
        RECT 9.220 0.440 9.510 0.500 ;
        RECT 10.420 0.670 10.710 0.730 ;
        RECT 10.420 0.500 10.480 0.670 ;
        RECT 10.650 0.500 10.710 0.670 ;
        RECT 10.420 0.440 10.710 0.500 ;
  END
END SUTHERLAND1989
END LIBRARY

