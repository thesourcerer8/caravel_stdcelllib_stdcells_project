magic
tech sky130A
timestamp 1624067235
<< nwell >>
rect 0 179 720 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
<< ndiff >>
rect 82 67 111 73
rect 82 66 88 67
rect 58 50 88 66
rect 105 66 111 67
rect 322 67 351 73
rect 322 66 328 67
rect 105 50 137 66
rect 58 24 137 50
rect 152 49 281 66
rect 152 32 184 49
rect 201 32 281 49
rect 152 24 281 32
rect 296 50 328 66
rect 345 66 351 67
rect 514 67 543 73
rect 514 66 520 67
rect 345 50 425 66
rect 296 24 425 50
rect 440 50 520 66
rect 537 66 543 67
rect 610 67 639 73
rect 610 66 616 67
rect 537 50 569 66
rect 440 24 569 50
rect 584 50 616 66
rect 633 66 639 67
rect 633 50 663 66
rect 584 24 663 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 88 243
rect 105 226 137 243
rect 58 225 137 226
rect 152 225 281 309
rect 296 301 425 309
rect 296 284 328 301
rect 345 284 425 301
rect 296 225 425 284
rect 440 225 569 309
rect 584 243 663 309
rect 584 226 616 243
rect 633 226 663 243
rect 584 225 663 226
rect 82 220 111 225
rect 610 220 639 225
<< ndiffc >>
rect 88 50 105 67
rect 184 32 201 49
rect 328 50 345 67
rect 520 50 537 67
rect 616 50 633 67
<< pdiffc >>
rect 88 226 105 243
rect 328 284 345 301
rect 616 226 633 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
<< locali >>
rect 320 301 353 309
rect 320 284 328 301
rect 345 284 353 301
rect 320 276 353 284
rect 80 243 113 251
rect 80 226 88 243
rect 105 226 113 243
rect 608 243 641 251
rect 608 226 616 243
rect 633 226 641 243
rect 80 218 111 226
rect 610 218 641 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 128 108 161 116
rect 128 92 136 108
rect 130 91 136 92
rect 153 91 161 108
rect 130 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 560 108 593 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 92 568 108
rect 520 75 537 91
rect 562 91 568 92
rect 585 91 593 108
rect 562 83 593 91
rect 80 67 113 75
rect 80 50 88 67
rect 105 50 113 67
rect 322 67 353 75
rect 322 66 328 67
rect 80 42 113 50
rect 176 49 209 57
rect 176 32 184 49
rect 201 32 209 49
rect 320 50 328 66
rect 345 50 353 67
rect 320 42 353 50
rect 512 67 545 75
rect 512 50 520 67
rect 537 50 545 67
rect 610 67 641 75
rect 610 66 616 67
rect 512 42 545 50
rect 608 50 616 66
rect 633 50 641 67
rect 608 42 641 50
rect 176 27 209 32
rect 176 24 184 27
rect 201 24 209 27
<< viali >>
rect 328 284 345 301
rect 88 226 105 243
rect 616 226 633 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 520 91 537 108
rect 568 91 585 108
rect 88 50 105 67
rect 328 50 345 67
rect 616 50 633 67
rect 184 10 201 27
<< metal1 >>
rect 0 309 720 357
rect 322 301 351 309
rect 322 284 328 301
rect 345 284 351 301
rect 322 278 351 284
rect 82 243 111 249
rect 82 226 88 243
rect 105 241 111 243
rect 610 243 639 249
rect 610 241 616 243
rect 105 227 616 241
rect 105 226 111 227
rect 82 220 111 226
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 137 114 151 178
rect 281 114 295 178
rect 425 114 439 178
rect 521 114 535 227
rect 610 226 616 227
rect 633 226 639 243
rect 610 220 639 226
rect 562 201 591 207
rect 562 184 568 201
rect 585 184 591 201
rect 562 178 591 184
rect 569 114 583 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 274 108 303 114
rect 274 91 280 108
rect 297 91 303 108
rect 274 85 303 91
rect 418 108 447 114
rect 418 91 424 108
rect 441 91 447 108
rect 418 85 447 91
rect 514 108 543 114
rect 514 91 520 108
rect 537 91 543 108
rect 514 85 543 91
rect 562 108 591 114
rect 562 91 568 108
rect 585 91 591 108
rect 562 85 591 91
rect 82 67 111 73
rect 82 50 88 67
rect 105 66 111 67
rect 322 67 351 73
rect 322 66 328 67
rect 105 52 328 66
rect 105 50 111 52
rect 82 44 111 50
rect 322 50 328 52
rect 345 66 351 67
rect 610 67 639 73
rect 610 66 616 67
rect 345 52 616 66
rect 345 50 351 52
rect 322 44 351 50
rect 610 50 616 52
rect 633 50 639 67
rect 610 44 639 50
rect 178 27 207 33
rect 178 24 184 27
rect 0 10 184 24
rect 201 24 207 27
rect 201 10 720 24
rect 0 -24 720 10
<< labels >>
rlabel metal1 0 309 720 357 0 VDD
port 1 se
rlabel metal1 0 -24 720 24 0 GND
port 2 se
rlabel metal1 514 85 543 114 0 Y
port 3 se
rlabel metal1 82 220 111 227 0 Y
port 4 se
rlabel metal1 521 114 535 227 0 Y
port 5 se
rlabel metal1 610 220 639 227 0 Y
port 6 se
rlabel metal1 82 227 639 241 0 Y
port 7 se
rlabel metal1 82 241 111 249 0 Y
port 8 se
rlabel metal1 610 241 639 249 0 Y
port 9 se
rlabel metal1 130 85 159 114 0 B
port 10 se
rlabel metal1 137 114 151 178 0 B
port 11 se
rlabel metal1 130 178 159 207 0 B
port 12 se
rlabel metal1 418 85 447 114 0 C
port 13 se
rlabel metal1 425 114 439 178 0 C
port 14 se
rlabel metal1 418 178 447 207 0 C
port 15 se
rlabel metal1 562 85 591 114 0 D
port 16 se
rlabel metal1 569 114 583 178 0 D
port 17 se
rlabel metal1 562 178 591 207 0 D
port 18 se
rlabel metal1 274 85 303 114 0 A
port 19 se
rlabel metal1 281 114 295 178 0 A
port 20 se
rlabel metal1 274 178 303 207 0 A
port 21 se
<< properties >>
string FIXED_BBOX 0 0 720 333
<< end >>
