VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.370 2.675 2.950 2.815 ;
        RECT 1.370 2.070 1.510 2.675 ;
        RECT 2.810 2.070 2.950 2.675 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 2.390500 ;
    PORT
      LAYER met1 ;
        RECT 0.575 0.440 0.865 0.730 ;
        RECT 3.215 0.440 3.505 0.730 ;
        RECT 6.095 0.440 6.385 0.730 ;
        RECT 8.975 0.440 9.265 0.730 ;
        RECT 11.855 0.440 12.145 0.730 ;
        RECT 0.650 0.240 0.790 0.440 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 6.170 0.240 6.310 0.440 ;
        RECT 9.050 0.240 9.190 0.440 ;
        RECT 11.930 0.240 12.070 0.440 ;
        RECT 0.000 -0.240 12.960 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 12.960 3.570 ;
        RECT 0.575 2.735 0.865 3.090 ;
        RECT 3.215 2.735 3.505 3.090 ;
        RECT 6.095 2.735 6.385 3.090 ;
        RECT 8.975 2.735 9.265 3.090 ;
        RECT 11.855 2.735 12.145 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 3.494400 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.155 3.215 12.805 3.245 ;
        RECT 0.155 3.090 3.025 3.215 ;
        RECT 3.695 3.090 12.805 3.215 ;
        RECT 0.555 2.715 0.885 3.090 ;
        RECT 6.075 2.715 6.405 3.090 ;
        RECT 8.955 2.715 9.285 3.090 ;
        RECT 11.835 2.715 12.165 3.090 ;
      LAYER mcon ;
        RECT 6.155 3.245 6.325 3.415 ;
        RECT 0.635 2.795 0.805 2.965 ;
        RECT 6.155 2.795 6.325 2.965 ;
        RECT 9.035 2.795 9.205 2.965 ;
        RECT 11.915 2.795 12.085 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 10.415 2.195 10.705 2.485 ;
        RECT 10.490 1.540 10.630 2.195 ;
        RECT 10.415 1.250 10.705 1.540 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 12.960 3.330 ;
      LAYER li1 ;
        RECT 3.195 2.715 3.525 3.045 ;
        RECT 1.755 2.260 2.085 2.505 ;
        RECT 1.775 2.175 2.085 2.260 ;
        RECT 4.635 2.175 4.965 2.505 ;
        RECT 7.515 2.260 7.845 2.505 ;
        RECT 10.395 2.260 10.725 2.505 ;
        RECT 7.535 2.175 7.845 2.260 ;
        RECT 10.415 2.175 10.725 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 2.005 4.465 2.090 ;
        RECT 4.155 1.760 4.485 2.005 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 11.355 1.760 11.685 2.090 ;
        RECT 2.795 1.155 2.965 1.760 ;
        RECT 5.675 1.155 5.845 1.760 ;
        RECT 8.555 1.155 8.725 1.760 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 2.715 0.825 3.025 0.920 ;
        RECT 4.155 0.825 4.485 1.155 ;
        RECT 5.595 0.920 5.925 1.155 ;
        RECT 7.035 0.920 7.365 1.155 ;
        RECT 8.475 0.920 8.805 1.155 ;
        RECT 9.915 0.920 10.245 1.155 ;
        RECT 5.595 0.825 5.905 0.920 ;
        RECT 7.035 0.825 7.345 0.920 ;
        RECT 8.475 0.825 8.785 0.920 ;
        RECT 9.915 0.825 10.225 0.920 ;
        RECT 10.475 0.750 10.645 1.480 ;
        RECT 11.355 0.920 11.685 1.155 ;
        RECT 11.355 0.825 11.665 0.920 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.775 0.655 2.085 0.750 ;
        RECT 1.755 0.420 2.085 0.655 ;
        RECT 3.195 0.420 3.525 0.750 ;
        RECT 4.655 0.655 4.965 0.750 ;
        RECT 4.635 0.420 4.965 0.655 ;
        RECT 6.075 0.420 6.405 0.750 ;
        RECT 7.515 0.420 7.845 0.750 ;
        RECT 8.955 0.420 9.285 0.750 ;
        RECT 10.395 0.420 10.725 0.750 ;
        RECT 11.835 0.420 12.165 0.750 ;
        RECT 0.155 0.085 12.805 0.240 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 3.275 2.795 3.445 2.965 ;
        RECT 1.835 2.255 2.005 2.425 ;
        RECT 4.715 2.255 4.885 2.425 ;
        RECT 7.595 2.255 7.765 2.425 ;
        RECT 10.475 2.255 10.645 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 5.675 1.840 5.845 2.010 ;
        RECT 7.115 1.840 7.285 2.010 ;
        RECT 8.555 1.840 8.725 2.010 ;
        RECT 9.995 1.840 10.165 2.010 ;
        RECT 11.435 1.840 11.605 2.010 ;
        RECT 10.475 1.310 10.645 1.480 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 7.115 0.905 7.285 1.075 ;
        RECT 9.995 0.905 10.165 1.075 ;
        RECT 11.435 0.905 11.605 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 6.155 0.500 6.325 0.670 ;
        RECT 7.595 0.500 7.765 0.670 ;
        RECT 9.035 0.500 9.205 0.670 ;
        RECT 11.915 0.500 12.085 0.670 ;
        RECT 6.155 -0.085 6.325 0.085 ;
      LAYER met1 ;
        RECT 4.250 2.675 5.830 2.815 ;
        RECT 1.775 2.195 2.065 2.485 ;
        RECT 1.850 1.060 1.990 2.195 ;
        RECT 4.250 2.070 4.390 2.675 ;
        RECT 4.655 2.195 4.945 2.485 ;
        RECT 4.175 1.780 4.465 2.070 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 1.850 0.920 4.465 1.060 ;
        RECT 1.850 0.730 1.990 0.920 ;
        RECT 4.175 0.845 4.465 0.920 ;
        RECT 4.730 1.060 4.870 2.195 ;
        RECT 5.690 2.070 5.830 2.675 ;
        RECT 7.130 2.675 8.710 2.815 ;
        RECT 7.130 2.070 7.270 2.675 ;
        RECT 7.535 2.195 7.825 2.485 ;
        RECT 5.615 1.780 5.905 2.070 ;
        RECT 7.055 1.780 7.345 2.070 ;
        RECT 7.130 1.135 7.270 1.780 ;
        RECT 7.055 1.060 7.345 1.135 ;
        RECT 4.730 0.920 7.345 1.060 ;
        RECT 4.730 0.730 4.870 0.920 ;
        RECT 7.055 0.845 7.345 0.920 ;
        RECT 7.610 1.060 7.750 2.195 ;
        RECT 8.570 2.070 8.710 2.675 ;
        RECT 8.495 1.780 8.785 2.070 ;
        RECT 9.935 1.780 10.225 2.070 ;
        RECT 11.375 1.780 11.665 2.070 ;
        RECT 10.010 1.135 10.150 1.780 ;
        RECT 11.450 1.135 11.590 1.780 ;
        RECT 9.935 1.060 10.225 1.135 ;
        RECT 11.375 1.060 11.665 1.135 ;
        RECT 7.610 0.920 11.665 1.060 ;
        RECT 7.610 0.730 7.750 0.920 ;
        RECT 9.935 0.845 10.225 0.920 ;
        RECT 11.375 0.845 11.665 0.920 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 4.655 0.440 4.945 0.730 ;
        RECT 7.535 0.440 7.825 0.730 ;
  END
END CLKBUF1
END LIBRARY

