VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO or
  CLASS BLOCK ;
  FOREIGN or ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  PIN VDD
    ANTENNAGATEAREA 0.567000 ;
    ANTENNADIFFAREA 4.227600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 3.200 2.740 3.530 3.090 ;
        RECT 0.800 2.260 1.130 2.510 ;
        RECT 0.800 2.180 1.110 2.260 ;
        RECT 4.640 2.180 4.970 2.510 ;
        RECT 1.280 1.760 1.610 2.090 ;
        RECT 2.720 1.760 3.050 2.090 ;
        RECT 4.160 2.010 4.470 2.090 ;
        RECT 4.160 1.760 4.490 2.010 ;
        RECT 1.280 0.830 1.610 1.160 ;
        RECT 2.720 0.920 3.050 1.160 ;
        RECT 2.740 0.830 3.050 0.920 ;
        RECT 4.160 0.920 4.490 1.160 ;
        RECT 4.160 0.830 4.470 0.920 ;
        RECT 0.560 0.260 0.890 0.590 ;
        RECT 2.240 0.420 2.570 0.750 ;
        RECT 3.200 0.240 3.530 0.590 ;
        RECT 4.640 0.420 4.970 0.750 ;
        RECT 0.000 0.090 0.390 0.240 ;
        RECT 1.060 0.090 5.760 0.240 ;
        RECT 0.000 -0.240 5.760 0.090 ;
      LAYER mcon ;
        RECT 0.160 3.250 0.330 3.420 ;
        RECT 0.640 3.250 0.810 3.420 ;
        RECT 1.120 3.250 1.290 3.420 ;
        RECT 1.600 3.250 1.770 3.420 ;
        RECT 2.080 3.250 2.250 3.420 ;
        RECT 2.560 3.250 2.730 3.420 ;
        RECT 3.040 3.250 3.210 3.420 ;
        RECT 3.520 3.250 3.690 3.420 ;
        RECT 4.000 3.250 4.170 3.420 ;
        RECT 4.480 3.250 4.650 3.420 ;
        RECT 4.960 3.250 5.130 3.420 ;
        RECT 5.440 3.250 5.610 3.420 ;
        RECT 3.280 2.820 3.450 2.990 ;
        RECT 0.880 2.260 1.050 2.430 ;
        RECT 4.720 2.260 4.890 2.430 ;
        RECT 1.360 1.840 1.530 2.010 ;
        RECT 2.800 1.840 2.970 2.010 ;
        RECT 4.240 1.840 4.410 2.010 ;
        RECT 1.360 0.910 1.530 1.080 ;
        RECT 2.800 0.910 2.970 1.080 ;
        RECT 4.240 0.910 4.410 1.080 ;
        RECT 0.640 0.340 0.810 0.510 ;
        RECT 2.320 0.500 2.490 0.670 ;
        RECT 4.720 0.500 4.890 0.670 ;
        RECT 0.160 -0.090 0.330 0.090 ;
        RECT 0.640 -0.090 0.810 0.090 ;
        RECT 1.120 -0.090 1.290 0.090 ;
        RECT 1.600 -0.090 1.770 0.090 ;
        RECT 2.080 -0.090 2.250 0.090 ;
        RECT 2.560 -0.090 2.730 0.090 ;
        RECT 3.040 -0.090 3.210 0.090 ;
        RECT 3.520 -0.090 3.690 0.090 ;
        RECT 4.000 -0.090 4.170 0.090 ;
        RECT 4.480 -0.090 4.650 0.090 ;
        RECT 4.960 -0.090 5.130 0.090 ;
        RECT 5.440 -0.090 5.610 0.090 ;
      LAYER met1 ;
        RECT 0.000 -0.240 5.760 3.570 ;
    END
  END VDD
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 5.760 3.330 ;
  END
END or
END LIBRARY

