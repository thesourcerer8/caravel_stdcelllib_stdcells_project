magic
tech sky130A
timestamp 1623602999
<< nwell >>
rect 0 179 720 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
<< ndiff >>
rect 82 66 111 69
rect 370 66 399 69
rect 514 66 543 69
rect 610 66 639 69
rect 58 63 137 66
rect 58 46 88 63
rect 105 46 137 63
rect 58 24 137 46
rect 152 36 281 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 281 36
rect 296 63 425 66
rect 296 46 376 63
rect 393 46 425 63
rect 296 24 425 46
rect 440 63 569 66
rect 440 46 520 63
rect 537 46 569 63
rect 440 24 569 46
rect 584 63 663 66
rect 584 46 616 63
rect 633 46 663 63
rect 584 24 663 46
rect 201 19 207 24
rect 178 13 207 19
<< pdiff >>
rect 322 309 351 312
rect 58 238 137 309
rect 58 225 88 238
rect 82 221 88 225
rect 105 225 137 238
rect 152 225 281 309
rect 296 306 425 309
rect 296 289 328 306
rect 345 289 425 306
rect 296 225 425 289
rect 440 225 569 309
rect 584 238 663 309
rect 584 225 616 238
rect 105 221 111 225
rect 82 215 111 221
rect 610 221 616 225
rect 633 225 663 238
rect 633 221 639 225
rect 610 215 639 221
<< ndiffc >>
rect 88 46 105 63
rect 184 19 201 36
rect 376 46 393 63
rect 520 46 537 63
rect 616 46 633 63
<< pdiffc >>
rect 88 221 105 238
rect 328 289 345 306
rect 616 221 633 238
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 569 309 584 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 569 206 584 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 569 66 584 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
<< locali >>
rect 320 306 353 314
rect 320 289 328 306
rect 345 289 353 306
rect 320 281 353 289
rect 80 238 113 246
rect 80 221 88 238
rect 105 223 113 238
rect 608 238 641 246
rect 608 223 616 238
rect 105 221 111 223
rect 80 213 111 221
rect 610 221 616 223
rect 633 221 641 238
rect 610 213 641 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 128 103 161 111
rect 128 88 136 103
rect 130 86 136 88
rect 153 86 161 103
rect 130 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 560 103 593 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 88 568 103
rect 520 71 537 86
rect 562 86 568 88
rect 585 86 593 103
rect 562 78 593 86
rect 80 63 113 71
rect 80 46 88 63
rect 105 46 113 63
rect 80 38 113 46
rect 368 63 399 71
rect 368 46 376 63
rect 393 61 399 63
rect 512 63 545 71
rect 393 46 401 61
rect 176 36 209 44
rect 368 38 401 46
rect 512 46 520 63
rect 537 46 545 63
rect 610 63 641 71
rect 610 61 616 63
rect 512 38 545 46
rect 608 46 616 61
rect 633 46 641 63
rect 608 38 641 46
rect 176 11 184 36
rect 201 11 209 36
<< viali >>
rect 328 289 345 306
rect 88 221 105 238
rect 616 221 633 238
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 520 86 537 103
rect 568 86 585 103
rect 88 46 105 63
rect 376 46 393 63
rect 616 46 633 63
rect 184 19 201 22
rect 184 5 201 19
<< metal1 >>
rect 0 309 720 357
rect 322 306 351 309
rect 322 289 328 306
rect 345 289 351 306
rect 322 283 351 289
rect 82 238 111 244
rect 82 221 88 238
rect 105 237 111 238
rect 610 238 639 244
rect 610 237 616 238
rect 105 223 616 237
rect 105 221 111 223
rect 82 215 111 221
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 274 198 303 204
rect 274 181 280 198
rect 297 181 303 198
rect 274 175 303 181
rect 418 198 447 204
rect 418 181 424 198
rect 441 181 447 198
rect 418 175 447 181
rect 137 109 151 175
rect 281 109 295 175
rect 425 109 439 175
rect 521 109 535 223
rect 610 221 616 223
rect 633 221 639 238
rect 610 215 639 221
rect 562 198 591 204
rect 562 181 568 198
rect 585 181 591 198
rect 562 175 591 181
rect 569 109 583 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 86 159 103
rect 130 80 159 86
rect 274 103 303 109
rect 274 86 280 103
rect 297 86 303 103
rect 274 80 303 86
rect 418 103 447 109
rect 418 86 424 103
rect 441 86 447 103
rect 418 80 447 86
rect 514 103 543 109
rect 514 86 520 103
rect 537 86 543 103
rect 514 80 543 86
rect 562 103 591 109
rect 562 86 568 103
rect 585 86 591 103
rect 562 80 591 86
rect 82 63 111 69
rect 82 46 88 63
rect 105 61 111 63
rect 370 63 399 69
rect 370 61 376 63
rect 105 47 376 61
rect 105 46 111 47
rect 82 40 111 46
rect 370 46 376 47
rect 393 61 399 63
rect 610 63 639 69
rect 610 61 616 63
rect 393 47 616 61
rect 393 46 399 47
rect 370 40 399 46
rect 610 46 616 47
rect 633 46 639 63
rect 610 40 639 46
rect 178 24 207 28
rect 0 22 720 24
rect 0 5 184 22
rect 201 5 720 22
rect 0 -24 720 5
<< labels >>
rlabel metal1 0 309 720 357 0 VDD
port 1 se
rlabel metal1 0 -24 720 24 0 GND
port 2 se
rlabel metal1 514 80 543 109 0 Y
port 3 se
rlabel metal1 82 215 111 223 0 Y
port 4 se
rlabel metal1 521 109 535 223 0 Y
port 5 se
rlabel metal1 610 215 639 223 0 Y
port 6 se
rlabel metal1 82 223 639 237 0 Y
port 7 se
rlabel metal1 82 237 111 244 0 Y
port 8 se
rlabel metal1 610 237 639 244 0 Y
port 9 se
rlabel metal1 130 80 159 109 0 B
port 10 se
rlabel metal1 137 109 151 175 0 B
port 11 se
rlabel metal1 130 175 159 204 0 B
port 12 se
rlabel metal1 562 80 591 109 0 D
port 13 se
rlabel metal1 569 109 583 175 0 D
port 14 se
rlabel metal1 562 175 591 204 0 D
port 15 se
rlabel metal1 418 80 447 109 0 C
port 16 se
rlabel metal1 425 109 439 175 0 C
port 17 se
rlabel metal1 418 175 447 204 0 C
port 18 se
rlabel metal1 274 80 303 109 0 A
port 19 se
rlabel metal1 281 109 295 175 0 A
port 20 se
rlabel metal1 274 175 303 204 0 A
port 21 se
<< properties >>
string FIXED_BBOX 0 0 720 333
<< end >>
