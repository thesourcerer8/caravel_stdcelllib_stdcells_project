MACRO VANBERKEL1991
 CLASS CORE ;
 FOREIGN VANBERKEL1991 0 0 ;
 SIZE 11.52 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
    END
  END GND

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 10.41500000 0.44000000 10.70500000 0.73000000 ;
        RECT 10.49000000 0.73000000 10.63000000 2.19500000 ;
        RECT 7.05500000 2.19500000 7.34500000 2.27000000 ;
        RECT 10.41500000 2.19500000 10.70500000 2.27000000 ;
        RECT 7.05500000 2.27000000 10.70500000 2.41000000 ;
        RECT 7.05500000 2.41000000 7.34500000 2.48500000 ;
        RECT 10.41500000 2.41000000 10.70500000 2.48500000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 2.73500000 0.84500000 3.02500000 0.92000000 ;
        RECT 8.49500000 0.84500000 8.78500000 0.92000000 ;
        RECT 2.73500000 0.92000000 8.78500000 1.06000000 ;
        RECT 2.73500000 1.06000000 3.02500000 1.13500000 ;
        RECT 8.49500000 1.06000000 8.78500000 1.13500000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 3.21500000 0.44000000 3.50500000 0.51500000 ;
        RECT 1.37000000 0.51500000 3.50500000 0.65500000 ;
        RECT 3.21500000 0.65500000 3.50500000 0.73000000 ;
        RECT 1.37000000 0.65500000 1.51000000 0.84500000 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 7.11500000 0.90500000 7.28500000 1.07500000 ;
     RECT 8.55500000 0.90500000 8.72500000 1.07500000 ;
     RECT 9.99500000 0.90500000 10.16500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 7.11500000 1.84000000 7.28500000 2.01000000 ;
     RECT 8.55500000 1.84000000 8.72500000 2.01000000 ;
     RECT 9.99500000 1.84000000 10.16500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 1.83500000 2.25500000 2.00500000 2.42500000 ;
     RECT 3.75500000 2.25500000 3.92500000 2.42500000 ;
     RECT 6.39500000 2.25500000 6.56500000 2.42500000 ;
     RECT 10.47500000 2.25500000 10.64500000 2.42500000 ;
     RECT 0.87500000 2.66000000 1.04500000 2.83000000 ;
     RECT 7.59500000 2.66000000 7.76500000 2.83000000 ;
     RECT 4.71500000 2.79500000 4.88500000 2.96500000 ;
     RECT 9.03500000 2.79500000 9.20500000 2.96500000 ;

    LAYER ndiffc ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 1.83500000 0.50000000 2.00500000 0.67000000 ;
     RECT 3.75500000 0.50000000 3.92500000 0.67000000 ;
     RECT 4.71500000 0.50000000 4.88500000 0.67000000 ;
     RECT 6.39500000 0.50000000 6.56500000 0.67000000 ;
     RECT 8.07500000 0.50000000 8.24500000 0.67000000 ;
     RECT 9.03500000 0.50000000 9.20500000 0.67000000 ;
     RECT 10.47500000 0.50000000 10.64500000 0.67000000 ;

    LAYER li1 ;
     RECT 0.55500000 0.42000000 0.88500000 0.75000000 ;
     RECT 3.67500000 0.42000000 4.00500000 0.75000000 ;
     RECT 6.31500000 0.42000000 6.64500000 0.75000000 ;
     RECT 7.99500000 0.42000000 8.32500000 0.75000000 ;
     RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
     RECT 4.71500000 0.24000000 4.88500000 0.42000000 ;
     RECT 9.03500000 0.24000000 9.20500000 0.42000000 ;
     RECT 4.63500000 0.42000000 4.96500000 0.75000000 ;
     RECT 8.95500000 0.42000000 9.28500000 0.75000000 ;
     RECT 10.39500000 0.42000000 10.72500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 9.91500000 0.82500000 10.24500000 1.15500000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 2.79500000 1.15500000 2.96500000 1.76000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 3.27500000 0.50000000 3.44500000 1.04000000 ;
     RECT 4.15500000 0.82500000 4.48500000 1.04000000 ;
     RECT 3.27500000 1.04000000 4.48500000 1.15500000 ;
     RECT 3.27500000 1.15500000 4.40500000 1.21000000 ;
     RECT 4.23500000 1.21000000 4.40500000 1.76000000 ;
     RECT 4.15500000 1.76000000 4.48500000 2.09000000 ;
     RECT 8.47500000 0.82500000 8.80500000 1.15500000 ;
     RECT 8.55500000 1.15500000 8.72500000 1.76000000 ;
     RECT 8.47500000 1.76000000 8.80500000 2.09000000 ;
     RECT 9.91500000 1.76000000 10.24500000 2.09000000 ;
     RECT 2.31500000 1.31000000 2.48500000 2.29000000 ;
     RECT 7.03500000 0.82500000 7.36500000 1.15500000 ;
     RECT 7.11500000 1.15500000 7.28500000 1.76000000 ;
     RECT 7.03500000 1.76000000 7.36500000 2.09000000 ;
     RECT 7.11500000 2.09000000 7.28500000 2.42500000 ;
     RECT 1.75500000 0.42000000 2.08500000 0.75000000 ;
     RECT 1.83500000 0.75000000 2.00500000 2.17500000 ;
     RECT 1.75500000 2.17500000 2.08500000 2.50500000 ;
     RECT 3.67500000 2.17500000 4.00500000 2.50500000 ;
     RECT 6.31500000 2.17500000 6.64500000 2.50500000 ;
     RECT 10.39500000 2.17500000 10.72500000 2.50500000 ;
     RECT 0.79500000 2.58000000 1.12500000 2.91000000 ;
     RECT 7.51500000 2.58000000 7.84500000 2.91000000 ;
     RECT 8.95500000 2.71500000 9.28500000 3.04500000 ;
     RECT 4.63500000 2.71500000 4.96500000 3.09000000 ;
     RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;

    LAYER viali ;
     RECT 9.03500000 -0.08500000 9.20500000 0.08500000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;
     RECT 3.75500000 0.50000000 3.92500000 0.67000000 ;
     RECT 6.39500000 0.50000000 6.56500000 0.67000000 ;
     RECT 8.07500000 0.50000000 8.24500000 0.67000000 ;
     RECT 10.47500000 0.50000000 10.64500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 8.55500000 0.90500000 8.72500000 1.07500000 ;
     RECT 9.99500000 0.90500000 10.16500000 1.07500000 ;
     RECT 2.31500000 1.31000000 2.48500000 1.48000000 ;
     RECT 1.83500000 1.71500000 2.00500000 1.88500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 9.99500000 1.84000000 10.16500000 2.01000000 ;
     RECT 2.31500000 2.12000000 2.48500000 2.29000000 ;
     RECT 3.75500000 2.25500000 3.92500000 2.42500000 ;
     RECT 6.39500000 2.25500000 6.56500000 2.42500000 ;
     RECT 7.11500000 2.25500000 7.28500000 2.42500000 ;
     RECT 10.47500000 2.25500000 10.64500000 2.42500000 ;
     RECT 0.87500000 2.66000000 1.04500000 2.83000000 ;
     RECT 7.59500000 2.66000000 7.76500000 2.83000000 ;
     RECT 9.03500000 2.79500000 9.20500000 2.96500000 ;
     RECT 4.71500000 3.24500000 4.88500000 3.41500000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 11.52000000 0.24000000 ;
     RECT 3.69500000 0.44000000 3.98500000 0.51500000 ;
     RECT 6.33500000 0.44000000 6.62500000 0.51500000 ;
     RECT 3.69500000 0.51500000 6.62500000 0.65500000 ;
     RECT 3.69500000 0.65500000 3.98500000 0.73000000 ;
     RECT 6.33500000 0.65500000 6.62500000 0.73000000 ;
     RECT 2.73500000 0.84500000 3.02500000 0.92000000 ;
     RECT 8.49500000 0.84500000 8.78500000 0.92000000 ;
     RECT 2.73500000 0.92000000 8.78500000 1.06000000 ;
     RECT 2.73500000 1.06000000 3.02500000 1.13500000 ;
     RECT 8.49500000 1.06000000 8.78500000 1.13500000 ;
     RECT 8.01500000 0.44000000 8.30500000 0.51500000 ;
     RECT 8.01500000 0.51500000 9.19000000 0.65500000 ;
     RECT 8.01500000 0.65500000 8.30500000 0.73000000 ;
     RECT 2.25500000 1.25000000 2.54500000 1.32500000 ;
     RECT 9.05000000 0.65500000 9.19000000 1.32500000 ;
     RECT 2.25500000 1.32500000 9.19000000 1.46500000 ;
     RECT 2.25500000 1.46500000 2.54500000 1.54000000 ;
     RECT 3.21500000 0.44000000 3.50500000 0.51500000 ;
     RECT 1.37000000 0.51500000 3.50500000 0.65500000 ;
     RECT 3.21500000 0.65500000 3.50500000 0.73000000 ;
     RECT 1.37000000 0.65500000 1.51000000 0.84500000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
     RECT 9.93500000 0.84500000 10.22500000 1.13500000 ;
     RECT 1.77500000 1.65500000 2.06500000 1.73000000 ;
     RECT 10.01000000 1.13500000 10.15000000 1.73000000 ;
     RECT 1.77500000 1.73000000 10.15000000 1.78000000 ;
     RECT 1.77500000 1.78000000 10.22500000 1.87000000 ;
     RECT 1.77500000 1.87000000 2.06500000 1.94500000 ;
     RECT 9.93500000 1.87000000 10.22500000 2.07000000 ;
     RECT 0.57500000 0.44000000 0.86500000 0.73000000 ;
     RECT 0.65000000 0.73000000 0.79000000 2.27000000 ;
     RECT 2.25500000 2.06000000 2.54500000 2.27000000 ;
     RECT 0.65000000 2.27000000 2.54500000 2.35000000 ;
     RECT 0.65000000 2.35000000 2.47000000 2.41000000 ;
     RECT 3.69500000 2.19500000 3.98500000 2.27000000 ;
     RECT 6.33500000 2.19500000 6.62500000 2.27000000 ;
     RECT 3.69500000 2.27000000 6.62500000 2.41000000 ;
     RECT 3.69500000 2.41000000 3.98500000 2.48500000 ;
     RECT 6.33500000 2.41000000 6.62500000 2.48500000 ;
     RECT 10.41500000 0.44000000 10.70500000 0.73000000 ;
     RECT 10.49000000 0.73000000 10.63000000 2.19500000 ;
     RECT 7.05500000 2.19500000 7.34500000 2.27000000 ;
     RECT 10.41500000 2.19500000 10.70500000 2.27000000 ;
     RECT 7.05500000 2.27000000 10.70500000 2.41000000 ;
     RECT 7.05500000 2.41000000 7.34500000 2.48500000 ;
     RECT 10.41500000 2.41000000 10.70500000 2.48500000 ;
     RECT 0.81500000 2.60000000 1.10500000 2.67500000 ;
     RECT 7.53500000 2.60000000 7.82500000 2.67500000 ;
     RECT 0.81500000 2.67500000 7.82500000 2.81500000 ;
     RECT 0.81500000 2.81500000 1.10500000 2.89000000 ;
     RECT 7.53500000 2.81500000 7.82500000 2.89000000 ;
     RECT 8.97500000 2.73500000 9.26500000 3.09000000 ;
     RECT 0.00000000 3.09000000 11.52000000 3.57000000 ;

 END
END VANBERKEL1991
