magic
tech sky130A
magscale 1 2
timestamp 1636809586
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 3744 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
rect 1713 48 1743 132
rect 2001 48 2031 132
rect 2289 48 2319 132
rect 2577 48 2607 132
rect 2865 48 2895 132
rect 3153 48 3183 132
rect 3441 48 3471 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
rect 1713 450 1743 618
rect 2001 450 2031 618
rect 2289 450 2319 618
rect 2577 450 2607 618
rect 2865 450 2895 618
rect 3153 450 3183 618
rect 3441 450 3471 618
<< ndiff >>
rect 115 134 173 146
rect 115 100 127 134
rect 161 132 173 134
rect 355 134 413 146
rect 355 132 367 134
rect 161 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 643 134 701 146
rect 643 132 655 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 100 655 132
rect 689 132 701 134
rect 931 134 989 146
rect 931 132 943 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 977 100 1137 132
rect 879 48 1137 100
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1507 134 1565 146
rect 1507 132 1519 134
rect 1265 100 1425 132
rect 1167 48 1425 100
rect 1455 100 1519 132
rect 1553 132 1565 134
rect 1795 134 1853 146
rect 1795 132 1807 134
rect 1553 100 1713 132
rect 1455 48 1713 100
rect 1743 100 1807 132
rect 1841 132 1853 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1841 100 2001 132
rect 1743 48 2001 100
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2371 134 2429 146
rect 2371 132 2383 134
rect 2129 100 2289 132
rect 2031 48 2289 100
rect 2319 100 2383 132
rect 2417 132 2429 134
rect 2659 134 2717 146
rect 2659 132 2671 134
rect 2417 100 2577 132
rect 2319 48 2577 100
rect 2607 100 2671 132
rect 2705 132 2717 134
rect 2947 134 3005 146
rect 2947 132 2959 134
rect 2705 100 2865 132
rect 2607 48 2865 100
rect 2895 100 2959 132
rect 2993 132 3005 134
rect 3235 134 3293 146
rect 3235 132 3247 134
rect 2993 100 3153 132
rect 2895 48 3153 100
rect 3183 100 3247 132
rect 3281 132 3293 134
rect 3523 134 3581 146
rect 3523 132 3535 134
rect 3281 100 3441 132
rect 3183 48 3441 100
rect 3471 100 3535 132
rect 3569 132 3581 134
rect 3569 100 3629 132
rect 3471 48 3629 100
<< pdiff >>
rect 115 593 273 618
rect 115 559 127 593
rect 161 559 273 593
rect 115 450 273 559
rect 303 485 561 618
rect 303 451 367 485
rect 401 451 561 485
rect 303 450 561 451
rect 591 593 849 618
rect 591 559 655 593
rect 689 559 849 593
rect 591 450 849 559
rect 879 485 1137 618
rect 879 451 943 485
rect 977 451 1137 485
rect 879 450 1137 451
rect 1167 593 1425 618
rect 1167 559 1231 593
rect 1265 559 1425 593
rect 1167 450 1425 559
rect 1455 485 1713 618
rect 1455 451 1519 485
rect 1553 451 1713 485
rect 1455 450 1713 451
rect 1743 593 2001 618
rect 1743 559 1807 593
rect 1841 559 2001 593
rect 1743 450 2001 559
rect 2031 485 2289 618
rect 2031 451 2095 485
rect 2129 451 2289 485
rect 2031 450 2289 451
rect 2319 593 2577 618
rect 2319 559 2383 593
rect 2417 559 2577 593
rect 2319 450 2577 559
rect 2607 485 2865 618
rect 2607 451 2671 485
rect 2705 451 2865 485
rect 2607 450 2865 451
rect 2895 593 3153 618
rect 2895 559 2959 593
rect 2993 559 3153 593
rect 2895 450 3153 559
rect 3183 485 3441 618
rect 3183 451 3247 485
rect 3281 451 3441 485
rect 3183 450 3441 451
rect 3471 593 3629 618
rect 3471 559 3535 593
rect 3569 559 3629 593
rect 3471 450 3629 559
rect 355 439 413 450
rect 931 439 989 450
rect 1507 439 1565 450
rect 2083 439 2141 450
rect 2659 439 2717 450
rect 3235 439 3293 450
<< ndiffc >>
rect 127 100 161 134
rect 367 100 401 134
rect 655 100 689 134
rect 943 100 977 134
rect 1231 100 1265 134
rect 1519 100 1553 134
rect 1807 100 1841 134
rect 2095 100 2129 134
rect 2383 100 2417 134
rect 2671 100 2705 134
rect 2959 100 2993 134
rect 3247 100 3281 134
rect 3535 100 3569 134
<< pdiffc >>
rect 127 559 161 593
rect 367 451 401 485
rect 655 559 689 593
rect 943 451 977 485
rect 1231 559 1265 593
rect 1519 451 1553 485
rect 1807 559 1841 593
rect 2095 451 2129 485
rect 2383 559 2417 593
rect 2671 451 2705 485
rect 2959 559 2993 593
rect 3247 451 3281 485
rect 3535 559 3569 593
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 2001 618 2031 644
rect 2289 618 2319 644
rect 2577 618 2607 644
rect 2865 618 2895 644
rect 3153 618 3183 644
rect 3441 618 3471 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 2001 418 2031 450
rect 2289 418 2319 450
rect 2577 418 2607 450
rect 2865 418 2895 450
rect 3153 418 3183 450
rect 3441 418 3471 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 2559 402 2625 418
rect 2559 368 2575 402
rect 2609 368 2625 402
rect 2559 352 2625 368
rect 2847 402 2913 418
rect 2847 368 2863 402
rect 2897 368 2913 402
rect 2847 352 2913 368
rect 3135 402 3201 418
rect 3135 368 3151 402
rect 3185 368 3201 402
rect 3135 352 3201 368
rect 3423 402 3489 418
rect 3423 368 3439 402
rect 3473 368 3489 402
rect 3423 352 3489 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 181 2337 215
rect 2271 165 2337 181
rect 2559 215 2625 231
rect 2559 181 2575 215
rect 2609 181 2625 215
rect 2559 165 2625 181
rect 2847 215 2913 231
rect 2847 181 2863 215
rect 2897 181 2913 215
rect 2847 165 2913 181
rect 3135 215 3201 231
rect 3135 181 3151 215
rect 3185 181 3201 215
rect 3135 165 3201 181
rect 3423 215 3489 231
rect 3423 181 3439 215
rect 3473 181 3489 215
rect 3423 165 3489 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 2001 132 2031 165
rect 2289 132 2319 165
rect 2577 132 2607 165
rect 2865 132 2895 165
rect 3153 132 3183 165
rect 3441 132 3471 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
rect 1713 22 1743 48
rect 2001 22 2031 48
rect 2289 22 2319 48
rect 2577 22 2607 48
rect 2865 22 2895 48
rect 3153 22 3183 48
rect 3441 22 3471 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 2287 368 2321 402
rect 2575 368 2609 402
rect 2863 368 2897 402
rect 3151 368 3185 402
rect 3439 368 3473 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 2287 181 2321 215
rect 2575 181 2609 215
rect 2863 181 2897 215
rect 3151 181 3185 215
rect 3439 181 3473 215
<< locali >>
rect 0 649 1807 683
rect 1841 649 3744 683
rect 31 643 3713 649
rect 31 618 605 643
rect 739 618 3713 643
rect 111 593 177 618
rect 111 559 127 593
rect 161 559 177 593
rect 111 543 177 559
rect 639 593 705 609
rect 639 559 655 593
rect 689 559 705 593
rect 1215 593 1281 618
rect 639 543 705 559
rect 1215 559 1231 593
rect 1265 559 1281 593
rect 1791 593 1857 618
rect 1215 543 1281 559
rect 351 485 417 501
rect 351 452 367 485
rect 355 451 367 452
rect 401 451 417 485
rect 355 435 417 451
rect 927 485 993 501
rect 927 451 943 485
rect 977 451 993 485
rect 927 435 993 451
rect 1135 418 1169 532
rect 1791 559 1807 593
rect 1841 559 1857 593
rect 2367 593 2433 618
rect 1791 543 1857 559
rect 1503 485 1569 501
rect 1503 452 1519 485
rect 1507 451 1519 452
rect 1553 451 1569 485
rect 1507 435 1569 451
rect 1711 418 1745 532
rect 2367 559 2383 593
rect 2417 559 2433 593
rect 2943 593 3009 618
rect 2367 543 2433 559
rect 2079 485 2145 501
rect 2079 452 2095 485
rect 2083 451 2095 452
rect 2129 451 2145 485
rect 2083 435 2145 451
rect 2287 418 2321 532
rect 2943 559 2959 593
rect 2993 559 3009 593
rect 2943 543 3009 559
rect 3519 593 3585 618
rect 3519 559 3535 593
rect 3569 559 3585 593
rect 3519 543 3585 559
rect 2655 485 2721 501
rect 2655 452 2671 485
rect 2659 451 2671 452
rect 2705 451 2721 485
rect 2659 435 2721 451
rect 2863 418 2897 532
rect 3231 485 3297 501
rect 3231 451 3247 485
rect 3281 451 3297 485
rect 3231 435 3297 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 893 418
rect 831 368 847 402
rect 881 401 893 402
rect 1119 402 1185 418
rect 881 368 897 401
rect 831 352 897 368
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 2559 402 2625 418
rect 2559 368 2575 402
rect 2609 368 2625 402
rect 2559 352 2625 368
rect 2847 402 2913 418
rect 2847 368 2863 402
rect 2897 368 2913 402
rect 2847 352 2913 368
rect 3135 402 3197 418
rect 3135 368 3151 402
rect 3185 401 3197 402
rect 3185 368 3201 401
rect 3135 352 3201 368
rect 559 231 593 352
rect 1135 323 1169 352
rect 1711 323 1745 352
rect 2287 323 2321 352
rect 2863 323 2897 352
rect 255 215 321 231
rect 255 181 271 215
rect 305 184 321 215
rect 543 215 609 231
rect 305 181 317 184
rect 255 165 317 181
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 1119 215 1185 231
rect 881 181 893 184
rect 831 165 893 181
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 184 1473 215
rect 1695 215 1761 231
rect 1457 181 1469 184
rect 1407 165 1469 181
rect 1695 181 1711 215
rect 1745 184 1761 215
rect 1983 215 2049 231
rect 1745 181 1757 184
rect 1695 165 1757 181
rect 1983 181 1999 215
rect 2033 184 2049 215
rect 2271 215 2337 231
rect 2033 181 2045 184
rect 1983 165 2045 181
rect 2271 181 2287 215
rect 2321 181 2337 215
rect 2271 165 2337 181
rect 2559 215 2625 231
rect 2559 181 2575 215
rect 2609 184 2625 215
rect 2847 215 2913 231
rect 2609 181 2621 184
rect 2559 165 2621 181
rect 2847 181 2863 215
rect 2897 184 2913 215
rect 3135 215 3201 231
rect 2897 181 2909 184
rect 2847 165 2909 181
rect 3135 181 3151 215
rect 3185 184 3201 215
rect 3185 181 3197 184
rect 3135 165 3197 181
rect 3247 150 3281 435
rect 3423 402 3489 418
rect 3423 368 3439 402
rect 3473 368 3489 402
rect 3423 352 3489 368
rect 3423 215 3489 231
rect 3423 181 3439 215
rect 3473 181 3489 215
rect 3423 165 3489 181
rect 111 134 177 150
rect 111 100 127 134
rect 161 100 177 134
rect 111 84 177 100
rect 351 134 417 150
rect 351 100 367 134
rect 401 100 417 134
rect 643 134 705 150
rect 643 131 655 134
rect 351 84 417 100
rect 639 100 655 131
rect 689 100 705 134
rect 639 84 705 100
rect 927 134 993 150
rect 927 100 943 134
rect 977 100 993 134
rect 1219 134 1281 150
rect 1219 131 1231 134
rect 927 84 993 100
rect 1215 100 1231 131
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 1503 134 1569 150
rect 1503 100 1519 134
rect 1553 100 1569 134
rect 1503 84 1569 100
rect 1791 134 1857 150
rect 1791 100 1807 134
rect 1841 100 1857 134
rect 1791 84 1857 100
rect 2079 134 2145 150
rect 2079 100 2095 134
rect 2129 100 2145 134
rect 2371 134 2433 150
rect 2371 131 2383 134
rect 2079 84 2145 100
rect 2367 100 2383 131
rect 2417 100 2433 134
rect 2367 84 2433 100
rect 2655 134 2721 150
rect 2655 100 2671 134
rect 2705 100 2721 134
rect 2655 84 2721 100
rect 2943 134 3009 150
rect 2943 100 2959 134
rect 2993 100 3009 134
rect 2943 84 3009 100
rect 3231 134 3297 150
rect 3231 100 3247 134
rect 3281 100 3297 134
rect 3523 134 3585 150
rect 3523 131 3535 134
rect 3231 84 3297 100
rect 3519 100 3535 131
rect 3569 100 3585 134
rect 3519 84 3585 100
rect 31 17 3713 48
rect 0 -17 655 17
rect 689 -17 3744 17
<< viali >>
rect 1807 649 1841 683
rect 127 559 161 593
rect 655 559 689 593
rect 1135 532 1169 566
rect 1231 559 1265 593
rect 367 451 401 485
rect 943 451 977 485
rect 1711 532 1745 566
rect 1807 559 1841 593
rect 1519 451 1553 485
rect 2287 532 2321 566
rect 2383 559 2417 593
rect 2095 451 2129 485
rect 2863 532 2897 566
rect 2959 559 2993 593
rect 3535 559 3569 593
rect 2671 451 2705 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1423 368 1457 402
rect 1999 368 2033 402
rect 2575 368 2609 402
rect 3151 368 3185 402
rect 1135 289 1169 323
rect 1711 289 1745 323
rect 2287 289 2321 323
rect 2863 289 2897 323
rect 271 181 305 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 2287 181 2321 215
rect 2575 181 2609 215
rect 2863 181 2897 215
rect 3151 181 3185 215
rect 3439 368 3473 402
rect 3439 181 3473 215
rect 127 100 161 134
rect 367 100 401 134
rect 655 100 689 134
rect 943 100 977 134
rect 1231 100 1265 134
rect 1519 100 1553 134
rect 1807 100 1841 134
rect 2095 100 2129 134
rect 2383 100 2417 134
rect 2671 100 2705 134
rect 2959 100 2993 134
rect 3247 100 3281 134
rect 3535 100 3569 134
rect 655 -17 689 17
<< metal1 >>
rect 0 683 3744 714
rect 0 649 1807 683
rect 1841 649 3744 683
rect 0 618 3744 649
rect 115 593 173 618
rect 115 559 127 593
rect 161 559 173 593
rect 643 593 701 618
rect 115 547 173 559
rect 274 535 590 563
rect 643 559 655 593
rect 689 559 701 593
rect 1219 593 1277 618
rect 1123 566 1181 578
rect 1123 563 1135 566
rect 643 547 701 559
rect 274 414 302 535
rect 355 485 413 497
rect 355 451 367 485
rect 401 451 413 485
rect 355 439 413 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 274 227 302 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 370 212 398 439
rect 562 414 590 535
rect 850 535 1135 563
rect 850 414 878 535
rect 1123 532 1135 535
rect 1169 532 1181 566
rect 1219 559 1231 593
rect 1265 559 1277 593
rect 1795 593 1853 618
rect 1699 566 1757 578
rect 1699 563 1711 566
rect 1219 547 1277 559
rect 1123 520 1181 532
rect 1426 535 1711 563
rect 931 485 989 497
rect 931 451 943 485
rect 977 451 989 485
rect 931 439 989 451
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 946 399 974 439
rect 1426 414 1454 535
rect 1699 532 1711 535
rect 1745 532 1757 566
rect 1795 559 1807 593
rect 1841 559 1853 593
rect 2371 593 2429 618
rect 2275 566 2333 578
rect 2275 563 2287 566
rect 1795 547 1853 559
rect 1699 520 1757 532
rect 2002 535 2287 563
rect 1507 485 1565 497
rect 1507 451 1519 485
rect 1553 451 1565 485
rect 1507 439 1565 451
rect 1411 402 1469 414
rect 1411 399 1423 402
rect 946 371 1423 399
rect 850 227 878 356
rect 835 215 893 227
rect 835 212 847 215
rect 370 184 847 212
rect 370 146 398 184
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 946 146 974 371
rect 1411 368 1423 371
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1522 399 1550 439
rect 2002 414 2030 535
rect 2275 532 2287 535
rect 2321 532 2333 566
rect 2371 559 2383 593
rect 2417 559 2429 593
rect 2947 593 3005 618
rect 2851 566 2909 578
rect 2851 563 2863 566
rect 2371 547 2429 559
rect 2275 520 2333 532
rect 2578 535 2863 563
rect 2083 485 2141 497
rect 2083 451 2095 485
rect 2129 451 2141 485
rect 2083 439 2141 451
rect 1987 402 2045 414
rect 1987 399 1999 402
rect 1522 371 1999 399
rect 1123 323 1181 335
rect 1123 289 1135 323
rect 1169 289 1181 323
rect 1123 277 1181 289
rect 1138 227 1166 277
rect 1426 227 1454 356
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 1411 215 1469 227
rect 1411 181 1423 215
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 1522 146 1550 371
rect 1987 368 1999 371
rect 2033 368 2045 402
rect 1987 356 2045 368
rect 2098 399 2126 439
rect 2578 414 2606 535
rect 2851 532 2863 535
rect 2897 532 2909 566
rect 2947 559 2959 593
rect 2993 559 3005 593
rect 2947 547 3005 559
rect 3523 593 3581 618
rect 3523 559 3535 593
rect 3569 559 3581 593
rect 3523 547 3581 559
rect 2851 520 2909 532
rect 2659 485 2717 497
rect 2659 451 2671 485
rect 2705 451 2717 485
rect 2659 439 2717 451
rect 2563 402 2621 414
rect 2563 399 2575 402
rect 2098 371 2575 399
rect 1699 323 1757 335
rect 1699 289 1711 323
rect 1745 289 1757 323
rect 1699 277 1757 289
rect 1714 227 1742 277
rect 2002 227 2030 356
rect 1699 215 1757 227
rect 1699 181 1711 215
rect 1745 181 1757 215
rect 1699 169 1757 181
rect 1987 215 2045 227
rect 1987 181 1999 215
rect 2033 181 2045 215
rect 1987 169 2045 181
rect 2098 146 2126 371
rect 2563 368 2575 371
rect 2609 368 2621 402
rect 2563 356 2621 368
rect 2674 399 2702 439
rect 3139 402 3197 414
rect 3139 399 3151 402
rect 2674 371 3151 399
rect 2275 323 2333 335
rect 2275 289 2287 323
rect 2321 289 2333 323
rect 2275 277 2333 289
rect 2290 227 2318 277
rect 2578 227 2606 356
rect 2275 215 2333 227
rect 2275 181 2287 215
rect 2321 181 2333 215
rect 2275 169 2333 181
rect 2563 215 2621 227
rect 2563 181 2575 215
rect 2609 181 2621 215
rect 2563 169 2621 181
rect 2674 146 2702 371
rect 3139 368 3151 371
rect 3185 399 3197 402
rect 3427 402 3485 414
rect 3427 399 3439 402
rect 3185 371 3439 399
rect 3185 368 3197 371
rect 3139 356 3197 368
rect 3427 368 3439 371
rect 3473 368 3485 402
rect 3427 356 3485 368
rect 2851 323 2909 335
rect 2851 289 2863 323
rect 2897 289 2909 323
rect 2851 277 2909 289
rect 2866 227 2894 277
rect 3154 227 3182 356
rect 3442 227 3470 356
rect 2851 215 2909 227
rect 2851 181 2863 215
rect 2897 181 2909 215
rect 2851 169 2909 181
rect 3139 215 3197 227
rect 3139 181 3151 215
rect 3185 181 3197 215
rect 3139 169 3197 181
rect 3427 215 3485 227
rect 3427 181 3439 215
rect 3473 181 3485 215
rect 3427 169 3485 181
rect 115 134 173 146
rect 115 100 127 134
rect 161 100 173 134
rect 115 88 173 100
rect 355 134 413 146
rect 355 100 367 134
rect 401 100 413 134
rect 355 88 413 100
rect 643 134 701 146
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 931 134 989 146
rect 931 100 943 134
rect 977 100 989 134
rect 931 88 989 100
rect 1219 134 1277 146
rect 1219 100 1231 134
rect 1265 100 1277 134
rect 1219 88 1277 100
rect 1507 134 1565 146
rect 1507 100 1519 134
rect 1553 100 1565 134
rect 1507 88 1565 100
rect 1795 134 1853 146
rect 1795 100 1807 134
rect 1841 100 1853 134
rect 1795 88 1853 100
rect 2083 134 2141 146
rect 2083 100 2095 134
rect 2129 100 2141 134
rect 2083 88 2141 100
rect 2371 134 2429 146
rect 2371 100 2383 134
rect 2417 100 2429 134
rect 2371 88 2429 100
rect 2659 134 2717 146
rect 2659 100 2671 134
rect 2705 100 2717 134
rect 2659 88 2717 100
rect 2947 134 3005 146
rect 2947 100 2959 134
rect 2993 100 3005 134
rect 2947 88 3005 100
rect 3235 134 3293 146
rect 3235 100 3247 134
rect 3281 100 3293 134
rect 3235 88 3293 100
rect 3523 134 3581 146
rect 3523 100 3535 134
rect 3569 100 3581 134
rect 3523 88 3581 100
rect 130 48 158 88
rect 658 48 686 88
rect 1234 48 1262 88
rect 1810 48 1838 88
rect 2386 48 2414 88
rect 2962 48 2990 88
rect 3538 48 3566 88
rect 0 17 3744 48
rect 0 -17 655 17
rect 689 -17 3744 17
rect 0 -48 3744 -17
<< labels >>
rlabel metal1 0 618 3744 714 0 VPWR
port 2 se
rlabel metal1 0 618 3744 714 0 VPWR
port 2 se
rlabel metal1 0 -48 3744 48 0 VGND
port 1 se
rlabel metal1 0 -48 3744 48 0 VGND
port 1 se
rlabel metal1 3235 88 3293 146 0 Y
port 3 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel metal1 547 356 605 414 0 A
port 0 se
rlabel metal1 274 414 302 535 0 A
port 0 se
rlabel metal1 562 414 590 535 0 A
port 0 se
rlabel metal1 274 535 590 563 0 A
port 0 se
rlabel locali 0 -17 3744 17 4 VGND
port 1 se ground default abutment
rlabel locali 31 17 3713 48 4 VGND
port 1 se ground default abutment
rlabel locali 0 649 3744 683 4 VPWR
port 2 se power default abutment
rlabel metal1 31 618 3713 649 4 VGND
port 1 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 3744 666
<< end >>
