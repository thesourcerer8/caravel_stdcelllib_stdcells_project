VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 1.780 3.010 2.070 3.090 ;
        RECT 1.780 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.070 3.010 ;
        RECT 1.780 2.780 2.070 2.840 ;
        RECT 4.660 3.010 4.950 3.090 ;
        RECT 4.660 2.840 4.720 3.010 ;
        RECT 4.890 2.840 4.950 3.010 ;
        RECT 4.660 2.780 4.950 2.840 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 0.490 4.950 0.550 ;
        RECT 4.660 0.320 4.720 0.490 ;
        RECT 4.890 0.320 4.950 0.490 ;
        RECT 4.660 0.240 4.950 0.320 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
  END vssd1
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.410 0.870 2.490 ;
        RECT 3.220 2.410 3.510 2.490 ;
        RECT 0.580 2.270 3.510 2.410 ;
        RECT 0.580 2.200 0.870 2.270 ;
        RECT 3.220 2.200 3.510 2.270 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 0.580 0.440 0.870 0.730 ;
    END
  END Y
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 2.740 0.850 3.030 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.780 4.470 2.070 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 4.180 0.850 4.470 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 3.010 2.090 3.090 ;
        RECT 1.760 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.090 3.010 ;
        RECT 1.760 2.760 2.090 2.840 ;
        RECT 4.640 3.010 4.970 3.090 ;
        RECT 4.640 2.840 4.720 3.010 ;
        RECT 4.890 2.840 4.970 3.010 ;
        RECT 4.640 2.760 4.970 2.840 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 3.200 2.430 3.530 2.510 ;
        RECT 3.200 2.260 3.280 2.430 ;
        RECT 3.450 2.260 3.530 2.430 ;
        RECT 3.200 2.180 3.530 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.030 2.090 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 4.640 0.490 4.970 0.570 ;
        RECT 4.640 0.320 4.720 0.490 ;
        RECT 4.890 0.320 4.970 0.490 ;
        RECT 4.640 0.240 4.970 0.320 ;
  END
END NAND3X1
END LIBRARY

