magic
tech sky130A
timestamp 1624567880
<< nwell >>
rect 0 179 288 333
<< nmos >>
rect 137 24 152 66
<< pmos >>
rect 137 225 152 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 51 231 66
rect 152 34 184 51
rect 201 34 231 51
rect 152 24 231 34
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 299 231 309
rect 152 282 184 299
rect 201 282 231 299
rect 152 225 231 282
rect 58 220 87 225
<< ndiffc >>
rect 64 50 81 67
rect 184 34 201 51
<< pdiffc >>
rect 64 226 81 243
rect 184 282 201 299
<< poly >>
rect 137 309 152 322
rect 137 209 152 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 137 66 152 83
rect 137 11 152 24
<< polycont >>
rect 136 184 153 201
rect 136 91 153 108
<< locali >>
rect 0 342 288 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 288 342
rect 0 309 288 325
rect 176 299 209 309
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 56 42 89 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 176 24 209 34
rect 0 9 288 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 288 9
rect 0 -24 288 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 184 282 201 299
rect 64 226 81 243
rect 136 184 153 201
rect 136 91 153 108
rect 64 50 81 67
rect 184 34 201 51
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
<< metal1 >>
rect 0 342 288 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 288 342
rect 0 309 288 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 65 73 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 137 114 151 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 58 44 87 50
rect 178 51 207 57
rect 178 34 184 51
rect 201 34 207 51
rect 178 24 207 34
rect 0 9 288 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 288 9
rect 0 -24 288 -9
<< labels >>
rlabel metal1 65 73 79 220 0 Y
port 6 se
rlabel metal1 137 114 151 178 0 A
port 9 se
rlabel locali 0 309 288 357 0 VDD
port 1 se
rlabel metal1 0 309 288 357 0 VDD
port 2 se
rlabel locali 0 -24 288 24 0 GND
port 3 se
rlabel metal1 0 -24 288 24 0 GND
port 4 se
rlabel metal1 58 44 87 73 0 Y
port 5 se
rlabel metal1 58 220 87 249 0 Y
port 7 se
rlabel metal1 130 85 159 114 0 A
port 8 se
rlabel metal1 130 178 159 207 0 A
port 10 se
<< properties >>
string FIXED_BBOX 0 0 288 333
<< end >>
