magic
tech sky130A
timestamp 1623602822
<< nwell >>
rect 0 179 720 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
<< ndiff >>
rect 82 66 111 69
rect 610 66 639 69
rect 58 63 137 66
rect 58 46 88 63
rect 105 46 137 63
rect 58 24 137 46
rect 152 24 281 66
rect 296 36 425 66
rect 296 24 328 36
rect 322 19 328 24
rect 345 24 425 36
rect 440 24 569 66
rect 584 63 663 66
rect 584 46 616 63
rect 633 46 663 63
rect 584 24 663 46
rect 345 19 351 24
rect 322 13 351 19
<< pdiff >>
rect 178 309 207 312
rect 58 238 137 309
rect 58 225 88 238
rect 82 221 88 225
rect 105 225 137 238
rect 152 306 281 309
rect 152 289 184 306
rect 201 289 281 306
rect 152 225 281 289
rect 296 238 425 309
rect 296 225 328 238
rect 105 221 111 225
rect 82 215 111 221
rect 322 221 328 225
rect 345 225 425 238
rect 440 238 569 309
rect 440 225 472 238
rect 345 221 351 225
rect 322 215 351 221
rect 466 221 472 225
rect 489 225 569 238
rect 584 279 663 309
rect 584 262 616 279
rect 633 262 663 279
rect 584 225 663 262
rect 489 221 495 225
rect 466 215 495 221
<< ndiffc >>
rect 88 46 105 63
rect 328 19 345 36
rect 616 46 633 63
<< pdiffc >>
rect 88 221 105 238
rect 184 289 201 306
rect 328 221 345 238
rect 472 221 489 238
rect 616 262 633 279
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 569 309 584 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 569 206 584 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 569 66 584 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 608 279 641 287
rect 608 262 616 279
rect 633 262 641 279
rect 608 254 641 262
rect 80 238 113 246
rect 80 221 88 238
rect 105 221 113 238
rect 320 238 353 246
rect 320 223 328 238
rect 80 213 113 221
rect 322 221 328 223
rect 345 221 353 238
rect 464 238 497 246
rect 464 223 472 238
rect 322 213 353 221
rect 466 221 472 223
rect 489 221 497 238
rect 466 213 497 221
rect 130 198 161 206
rect 130 196 136 198
rect 128 181 136 196
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 88 593 103
rect 585 86 591 88
rect 560 78 591 86
rect 80 63 111 71
rect 80 46 88 63
rect 105 61 111 63
rect 608 63 641 71
rect 105 46 113 61
rect 80 38 113 46
rect 608 46 616 63
rect 633 46 641 63
rect 320 36 353 44
rect 608 38 641 46
rect 320 11 328 36
rect 345 11 353 36
<< viali >>
rect 184 289 201 306
rect 616 262 633 279
rect 88 221 105 238
rect 328 221 345 238
rect 472 221 489 238
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
rect 88 46 105 63
rect 616 46 633 63
rect 328 19 345 22
rect 328 5 345 19
<< metal1 >>
rect 0 309 720 357
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 610 279 639 285
rect 610 277 616 279
rect 329 263 616 277
rect 329 244 343 263
rect 610 262 616 263
rect 633 262 639 279
rect 610 256 639 262
rect 82 238 111 244
rect 82 221 88 238
rect 105 237 111 238
rect 322 238 351 244
rect 322 237 328 238
rect 105 223 328 237
rect 105 221 111 223
rect 82 215 111 221
rect 322 221 328 223
rect 345 221 351 238
rect 322 215 351 221
rect 466 238 495 244
rect 466 221 472 238
rect 489 221 495 238
rect 466 215 495 221
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 274 198 303 204
rect 274 181 280 198
rect 297 181 303 198
rect 274 175 303 181
rect 418 198 447 204
rect 418 181 424 198
rect 441 181 447 198
rect 418 175 447 181
rect 137 109 151 175
rect 281 109 295 175
rect 425 109 439 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 86 159 103
rect 130 80 159 86
rect 274 103 303 109
rect 274 86 280 103
rect 297 86 303 103
rect 274 80 303 86
rect 418 103 447 109
rect 418 86 424 103
rect 441 86 447 103
rect 418 80 447 86
rect 82 63 111 69
rect 82 46 88 63
rect 105 61 111 63
rect 473 61 487 215
rect 562 198 591 204
rect 562 181 568 198
rect 585 181 591 198
rect 562 175 591 181
rect 569 109 583 175
rect 562 103 591 109
rect 562 86 568 103
rect 585 86 591 103
rect 562 80 591 86
rect 610 63 639 69
rect 610 61 616 63
rect 105 47 616 61
rect 105 46 111 47
rect 82 40 111 46
rect 610 46 616 47
rect 633 46 639 63
rect 610 40 639 46
rect 322 24 351 28
rect 0 22 720 24
rect 0 5 328 22
rect 345 5 720 22
rect 0 -24 720 5
<< labels >>
rlabel metal1 0 309 720 357 0 VDD
port 1 se
rlabel metal1 0 -24 720 24 0 GND
port 2 se
rlabel metal1 82 40 111 47 0 Y
port 3 se
rlabel metal1 610 40 639 47 0 Y
port 4 se
rlabel metal1 82 47 639 61 0 Y
port 5 se
rlabel metal1 82 61 111 69 0 Y
port 6 se
rlabel metal1 610 61 639 69 0 Y
port 7 se
rlabel metal1 473 61 487 215 0 Y
port 8 se
rlabel metal1 466 215 495 244 0 Y
port 9 se
rlabel metal1 130 80 159 109 0 B
port 10 se
rlabel metal1 137 109 151 175 0 B
port 11 se
rlabel metal1 130 175 159 204 0 B
port 12 se
rlabel metal1 274 80 303 109 0 A
port 13 se
rlabel metal1 281 109 295 175 0 A
port 14 se
rlabel metal1 274 175 303 204 0 A
port 15 se
rlabel metal1 418 80 447 109 0 C
port 16 se
rlabel metal1 425 109 439 175 0 C
port 17 se
rlabel metal1 418 175 447 204 0 C
port 18 se
rlabel metal1 562 80 591 109 0 D
port 19 se
rlabel metal1 569 109 583 175 0 D
port 20 se
rlabel metal1 562 175 591 204 0 D
port 21 se
<< properties >>
string FIXED_BBOX 0 0 720 333
<< end >>
