magic
tech sky130A
timestamp 1624574541
<< nwell >>
rect 0 179 576 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
<< ndiff >>
rect 82 67 111 73
rect 82 66 88 67
rect 58 50 88 66
rect 105 66 111 67
rect 466 67 495 73
rect 466 66 472 67
rect 105 50 137 66
rect 58 24 137 50
rect 152 24 281 66
rect 296 51 425 66
rect 296 34 328 51
rect 345 34 425 51
rect 296 24 425 34
rect 440 50 472 66
rect 489 66 495 67
rect 489 50 519 66
rect 440 24 519 50
<< pdiff >>
rect 58 299 137 309
rect 58 282 64 299
rect 81 282 137 299
rect 58 225 137 282
rect 152 243 281 309
rect 152 226 184 243
rect 201 226 281 243
rect 152 225 281 226
rect 296 299 425 309
rect 296 282 328 299
rect 345 282 425 299
rect 296 225 425 282
rect 440 243 519 309
rect 440 226 472 243
rect 489 226 519 243
rect 440 225 519 226
rect 178 220 207 225
rect 466 220 495 225
<< ndiffc >>
rect 88 50 105 67
rect 328 34 345 51
rect 472 50 489 67
<< pdiffc >>
rect 64 282 81 299
rect 184 226 201 243
rect 328 282 345 299
rect 472 226 489 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
<< locali >>
rect 0 342 576 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 576 342
rect 0 309 576 325
rect 56 299 89 309
rect 56 282 64 299
rect 81 282 89 299
rect 56 274 89 282
rect 320 299 353 309
rect 320 282 328 299
rect 345 282 353 299
rect 320 274 353 282
rect 176 243 209 251
rect 176 226 184 243
rect 201 226 209 243
rect 176 218 209 226
rect 464 243 497 251
rect 464 226 472 243
rect 489 226 497 243
rect 464 218 497 226
rect 128 201 159 209
rect 272 201 305 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 447 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 280 116 297 176
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 92 449 108
rect 441 91 447 92
rect 416 83 447 91
rect 80 67 111 75
rect 80 50 88 67
rect 105 66 111 67
rect 464 67 497 75
rect 105 50 113 66
rect 80 42 113 50
rect 320 51 353 59
rect 320 34 328 51
rect 345 34 353 51
rect 464 50 472 67
rect 489 50 497 67
rect 464 42 497 50
rect 320 24 353 34
rect 0 9 576 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 576 9
rect 0 -24 576 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 448 325 465 342
rect 496 325 513 342
rect 544 325 561 342
rect 64 282 81 299
rect 328 282 345 299
rect 184 226 201 243
rect 472 226 489 243
rect 136 184 153 201
rect 424 184 441 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 88 50 105 67
rect 328 34 345 51
rect 472 50 489 67
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
rect 448 -9 465 9
rect 496 -9 513 9
rect 544 -9 561 9
<< metal1 >>
rect 0 342 576 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 448 342
rect 465 325 496 342
rect 513 325 544 342
rect 561 325 576 342
rect 0 309 576 325
rect 58 299 87 309
rect 58 282 64 299
rect 81 282 87 299
rect 58 276 87 282
rect 322 299 351 309
rect 322 282 328 299
rect 345 282 351 299
rect 322 276 351 282
rect 178 243 207 249
rect 178 226 184 243
rect 201 226 207 243
rect 178 220 207 226
rect 466 243 495 249
rect 466 226 472 243
rect 489 226 495 243
rect 466 220 495 226
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 185 200 199 220
rect 418 201 447 207
rect 418 200 424 201
rect 185 186 424 200
rect 137 114 151 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 82 67 111 73
rect 82 50 88 67
rect 105 66 111 67
rect 185 66 199 186
rect 418 184 424 186
rect 441 184 447 201
rect 418 178 447 184
rect 425 114 439 178
rect 274 108 303 114
rect 274 91 280 108
rect 297 91 303 108
rect 274 85 303 91
rect 418 108 447 114
rect 418 91 424 108
rect 441 91 447 108
rect 418 85 447 91
rect 473 73 487 220
rect 105 52 199 66
rect 466 67 495 73
rect 105 50 111 52
rect 82 44 111 50
rect 322 51 351 57
rect 322 34 328 51
rect 345 34 351 51
rect 466 50 472 67
rect 489 50 495 67
rect 466 44 495 50
rect 322 24 351 34
rect 0 9 576 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 448 9
rect 465 -9 496 9
rect 513 -9 544 9
rect 561 -9 576 9
rect 0 -24 576 -9
<< labels >>
rlabel metal1 473 73 487 220 0 Y
port 6 se
rlabel metal1 137 114 151 178 0 A
port 9 se
rlabel locali 0 309 576 357 0 VDD
port 1 se
rlabel metal1 0 309 576 357 0 VDD
port 2 se
rlabel locali 0 -24 576 24 0 GND
port 3 se
rlabel metal1 0 -24 576 24 0 GND
port 4 se
rlabel metal1 466 44 495 73 0 Y
port 5 se
rlabel metal1 466 220 495 249 0 Y
port 7 se
rlabel metal1 130 85 159 114 0 A
port 8 se
rlabel metal1 130 178 159 207 0 A
port 10 se
rlabel metal1 274 85 303 114 0 B
port 11 se
<< properties >>
string FIXED_BBOX 0 0 576 333
<< end >>
