magic
tech sky130A
magscale 1 2
timestamp 1636809579
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1152 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
<< ndiff >>
rect 163 134 221 146
rect 163 132 175 134
rect 115 100 175 132
rect 209 132 221 134
rect 643 134 701 146
rect 643 132 655 134
rect 209 100 273 132
rect 115 48 273 100
rect 303 48 561 132
rect 591 100 655 132
rect 689 132 701 134
rect 931 134 989 146
rect 931 132 943 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 100 943 132
rect 977 132 989 134
rect 977 100 1037 132
rect 879 48 1037 100
<< pdiff >>
rect 115 593 273 618
rect 115 559 127 593
rect 161 559 273 593
rect 115 450 273 559
rect 303 485 561 618
rect 303 451 367 485
rect 401 451 561 485
rect 303 450 561 451
rect 591 593 849 618
rect 591 559 655 593
rect 689 559 849 593
rect 591 450 849 559
rect 879 485 1037 618
rect 879 451 943 485
rect 977 451 1037 485
rect 879 450 1037 451
rect 355 439 413 450
rect 931 439 989 450
<< ndiffc >>
rect 175 100 209 134
rect 655 100 689 134
rect 943 100 977 134
<< pdiffc >>
rect 127 559 161 593
rect 367 451 401 485
rect 655 559 689 593
rect 943 451 977 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
<< locali >>
rect 0 649 655 683
rect 689 649 1152 683
rect 31 643 1121 649
rect 31 618 605 643
rect 739 618 1121 643
rect 111 593 177 618
rect 111 559 127 593
rect 161 559 177 593
rect 111 543 177 559
rect 639 593 705 609
rect 639 559 655 593
rect 689 559 705 593
rect 639 543 705 559
rect 351 485 417 501
rect 351 452 367 485
rect 355 451 367 452
rect 401 451 417 485
rect 927 485 993 501
rect 927 452 943 485
rect 355 435 417 451
rect 931 451 943 452
rect 977 451 993 485
rect 931 435 993 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 559 323 593 352
rect 255 215 321 231
rect 255 184 271 215
rect 259 181 271 184
rect 305 181 321 215
rect 259 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 881 181 893 184
rect 831 165 893 181
rect 159 134 225 150
rect 159 100 175 134
rect 209 100 225 134
rect 643 134 705 150
rect 643 131 655 134
rect 159 84 225 100
rect 639 100 655 131
rect 689 100 705 134
rect 639 84 705 100
rect 927 134 993 150
rect 927 100 943 134
rect 977 100 993 134
rect 927 84 993 100
rect 31 17 1121 48
rect 0 -17 655 17
rect 689 -17 1152 17
<< viali >>
rect 655 649 689 683
rect 127 559 161 593
rect 655 559 689 593
rect 367 451 401 485
rect 943 451 977 485
rect 271 368 305 402
rect 847 368 881 402
rect 559 289 593 323
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 175 100 209 134
rect 655 100 689 134
rect 943 100 977 134
rect 655 -17 689 17
<< metal1 >>
rect 0 683 1152 714
rect 0 649 655 683
rect 689 649 1152 683
rect 0 618 1152 649
rect 115 593 173 618
rect 115 559 127 593
rect 161 559 173 593
rect 115 547 173 559
rect 643 593 701 618
rect 643 559 655 593
rect 689 559 701 593
rect 643 547 701 559
rect 355 485 413 497
rect 355 451 367 485
rect 401 451 413 485
rect 355 439 413 451
rect 931 485 989 497
rect 931 451 943 485
rect 977 451 989 485
rect 931 439 989 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 370 399 398 439
rect 835 402 893 414
rect 835 399 847 402
rect 370 371 847 399
rect 274 227 302 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 163 134 221 146
rect 163 100 175 134
rect 209 131 221 134
rect 370 131 398 371
rect 835 368 847 371
rect 881 368 893 402
rect 835 356 893 368
rect 547 323 605 335
rect 547 289 559 323
rect 593 289 605 323
rect 547 277 605 289
rect 562 227 590 277
rect 850 227 878 356
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 835 215 893 227
rect 835 181 847 215
rect 881 181 893 215
rect 835 169 893 181
rect 946 146 974 439
rect 209 103 398 131
rect 643 134 701 146
rect 209 100 221 103
rect 163 88 221 100
rect 643 100 655 134
rect 689 100 701 134
rect 643 88 701 100
rect 931 134 989 146
rect 931 100 943 134
rect 977 100 989 134
rect 931 88 989 100
rect 658 48 686 88
rect 0 17 1152 48
rect 0 -17 655 17
rect 689 -17 1152 17
rect 0 -48 1152 -17
<< labels >>
rlabel metal1 0 618 1152 714 0 VPWR
port 3 se
rlabel metal1 0 618 1152 714 0 VPWR
port 3 se
rlabel metal1 0 -48 1152 48 0 VGND
port 2 se
rlabel metal1 0 -48 1152 48 0 VGND
port 2 se
rlabel metal1 931 88 989 146 0 Y
port 4 se
rlabel metal1 946 146 974 439 0 Y
port 4 se
rlabel metal1 931 439 989 497 0 Y
port 4 se
rlabel metal1 547 169 605 227 0 B
port 1 se
rlabel metal1 562 227 590 277 0 B
port 1 se
rlabel metal1 547 277 605 335 0 B
port 1 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel locali 0 -17 1152 17 4 VGND
port 2 se ground default abutment
rlabel locali 31 17 1121 48 4 VGND
port 2 se ground default abutment
rlabel locali 0 649 1152 683 4 VPWR
port 3 se power default abutment
rlabel metal1 31 618 1121 649 4 VGND
port 2 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1152 666
<< end >>
