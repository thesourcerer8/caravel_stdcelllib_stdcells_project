magic
tech sky130A
timestamp 1623603012
<< nwell >>
rect 0 179 1008 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
rect 857 24 872 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
rect 857 225 872 309
<< ndiff >>
rect 58 66 87 69
rect 466 66 495 69
rect 898 66 927 69
rect 58 63 137 66
rect 58 46 64 63
rect 81 46 137 63
rect 58 24 137 46
rect 152 36 281 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 281 36
rect 296 24 425 66
rect 440 63 569 66
rect 440 46 472 63
rect 489 46 569 63
rect 440 24 569 46
rect 584 24 713 66
rect 728 36 857 66
rect 728 24 760 36
rect 201 19 207 24
rect 178 13 207 19
rect 754 19 760 24
rect 777 24 857 36
rect 872 63 951 66
rect 872 46 904 63
rect 921 46 951 63
rect 872 24 951 46
rect 777 19 783 24
rect 754 13 783 19
<< pdiff >>
rect 178 309 207 312
rect 754 309 783 312
rect 58 238 137 309
rect 58 221 64 238
rect 81 225 137 238
rect 152 306 281 309
rect 152 289 184 306
rect 201 289 281 306
rect 152 225 281 289
rect 296 225 425 309
rect 440 238 569 309
rect 440 225 472 238
rect 81 221 87 225
rect 58 215 87 221
rect 466 221 472 225
rect 489 225 569 238
rect 584 225 713 309
rect 728 306 857 309
rect 728 289 760 306
rect 777 289 857 306
rect 728 225 857 289
rect 872 238 951 309
rect 872 225 904 238
rect 489 221 495 225
rect 466 215 495 221
rect 898 221 904 225
rect 921 225 951 238
rect 921 221 927 225
rect 898 215 927 221
<< ndiffc >>
rect 64 46 81 63
rect 184 19 201 36
rect 472 46 489 63
rect 760 19 777 36
rect 904 46 921 63
<< pdiffc >>
rect 64 221 81 238
rect 184 289 201 306
rect 472 221 489 238
rect 760 289 777 306
rect 904 221 921 238
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 569 309 584 330
rect 713 309 728 330
rect 857 309 872 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 569 206 584 225
rect 713 206 728 225
rect 857 206 872 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 704 198 737 206
rect 704 181 712 198
rect 729 181 737 198
rect 704 173 737 181
rect 848 198 881 206
rect 848 181 856 198
rect 873 181 881 198
rect 848 173 881 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 704 103 737 111
rect 704 86 712 103
rect 729 86 737 103
rect 704 78 737 86
rect 848 103 881 111
rect 848 86 856 103
rect 873 86 881 103
rect 848 78 881 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 569 66 584 78
rect 713 66 728 78
rect 857 66 872 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
rect 857 11 872 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 712 181 729 198
rect 856 181 873 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
rect 712 86 729 103
rect 856 86 873 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 752 306 785 314
rect 752 289 760 306
rect 777 289 785 306
rect 752 281 785 289
rect 56 238 89 246
rect 56 221 64 238
rect 81 221 89 238
rect 56 213 89 221
rect 464 238 497 246
rect 464 221 472 238
rect 489 221 497 238
rect 896 238 929 246
rect 896 223 904 238
rect 464 218 497 221
rect 473 215 497 218
rect 898 221 904 223
rect 921 221 929 238
rect 898 213 929 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 201 447 206
rect 416 198 449 201
rect 560 198 593 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 174 449 181
rect 136 111 153 127
rect 280 111 297 173
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 56 63 89 71
rect 56 46 64 63
rect 81 46 89 63
rect 376 63 393 127
rect 424 111 441 140
rect 416 103 449 111
rect 416 86 424 103
rect 441 88 449 103
rect 441 86 447 88
rect 416 78 447 86
rect 472 71 489 181
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 704 198 737 206
rect 704 181 712 198
rect 729 181 737 198
rect 704 173 737 181
rect 848 198 881 206
rect 848 181 856 198
rect 873 181 881 198
rect 848 173 881 181
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 704 103 737 111
rect 704 86 712 103
rect 729 86 737 103
rect 704 78 737 86
rect 848 103 881 111
rect 848 86 856 103
rect 873 86 881 103
rect 848 78 881 86
rect 464 63 497 71
rect 464 46 472 63
rect 489 46 497 63
rect 568 63 585 78
rect 898 63 929 71
rect 898 61 904 63
rect 896 46 904 61
rect 921 46 929 63
rect 56 38 89 46
rect 176 36 209 44
rect 464 38 497 46
rect 176 19 184 36
rect 201 19 209 36
rect 176 11 209 19
rect 752 36 785 44
rect 896 38 929 46
rect 752 11 760 36
rect 777 11 785 36
<< viali >>
rect 184 289 201 306
rect 760 289 777 306
rect 64 221 81 238
rect 472 221 489 238
rect 904 221 921 238
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 472 181 489 198
rect 136 127 153 144
rect 376 127 393 144
rect 64 46 81 63
rect 424 140 441 157
rect 568 181 585 198
rect 712 181 729 198
rect 856 181 873 198
rect 712 86 729 103
rect 856 86 873 103
rect 376 46 393 63
rect 568 46 585 63
rect 904 46 921 63
rect 184 19 201 36
rect 760 19 777 22
rect 760 5 777 19
<< metal1 >>
rect 0 309 1008 357
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 754 306 783 309
rect 754 289 760 306
rect 777 289 783 306
rect 754 283 783 289
rect 58 238 87 244
rect 58 221 64 238
rect 81 221 87 238
rect 58 215 87 221
rect 466 238 495 244
rect 466 221 472 238
rect 489 221 495 238
rect 898 238 927 244
rect 898 237 904 238
rect 466 218 495 221
rect 569 223 904 237
rect 466 215 487 218
rect 65 102 79 215
rect 473 204 487 215
rect 569 204 583 223
rect 898 221 904 223
rect 921 221 927 238
rect 898 215 927 221
rect 130 198 159 204
rect 130 181 136 198
rect 153 196 159 198
rect 274 198 303 204
rect 274 196 280 198
rect 153 182 280 196
rect 153 181 159 182
rect 130 175 159 181
rect 274 181 280 182
rect 297 181 303 198
rect 418 198 447 204
rect 473 201 495 204
rect 418 196 424 198
rect 274 175 303 181
rect 377 182 424 196
rect 137 150 151 175
rect 377 150 391 182
rect 418 181 424 182
rect 441 181 447 198
rect 418 177 447 181
rect 466 198 495 201
rect 466 181 472 198
rect 489 181 495 198
rect 466 175 495 181
rect 562 198 591 204
rect 562 181 568 198
rect 585 181 591 198
rect 562 175 591 181
rect 706 198 735 204
rect 706 181 712 198
rect 729 181 735 198
rect 706 175 735 181
rect 850 198 879 204
rect 850 181 856 198
rect 873 181 879 198
rect 850 175 879 181
rect 418 157 447 163
rect 130 144 159 150
rect 130 127 136 144
rect 153 127 159 144
rect 130 121 159 127
rect 370 144 399 150
rect 370 127 376 144
rect 393 127 399 144
rect 418 140 424 157
rect 441 156 447 157
rect 569 156 583 175
rect 441 142 583 156
rect 441 140 447 142
rect 418 134 447 140
rect 370 121 399 127
rect 713 109 727 175
rect 857 109 871 175
rect 706 103 735 109
rect 706 102 712 103
rect 65 88 712 102
rect 65 69 79 88
rect 706 86 712 88
rect 729 86 735 103
rect 706 80 735 86
rect 850 103 879 109
rect 850 86 856 103
rect 873 86 879 103
rect 850 80 879 86
rect 58 63 87 69
rect 58 46 64 63
rect 81 46 87 63
rect 58 40 87 46
rect 370 63 399 69
rect 370 46 376 63
rect 393 61 399 63
rect 562 63 591 69
rect 562 61 568 63
rect 393 47 568 61
rect 393 46 399 47
rect 178 36 207 42
rect 370 40 399 46
rect 562 46 568 47
rect 585 61 591 63
rect 857 61 871 80
rect 905 69 919 215
rect 585 47 871 61
rect 898 63 927 69
rect 585 46 591 47
rect 562 40 591 46
rect 898 46 904 63
rect 921 46 927 63
rect 898 40 927 46
rect 178 24 184 36
rect 0 19 184 24
rect 201 24 207 36
rect 754 24 783 28
rect 201 22 1008 24
rect 201 19 760 22
rect 0 5 760 19
rect 777 5 1008 22
rect 0 -24 1008 5
<< labels >>
rlabel metal1 0 309 1008 357 0 VDD
port 1 se
rlabel metal1 0 -24 1008 24 0 GND
port 2 se
rlabel space 466 175 495 204 0 Y
port 3 se
rlabel metal1 473 204 487 215 0 Y
port 4 se
rlabel nwell 466 215 495 244 0 Y
port 5 se
rlabel metal1 370 40 399 47 0 A
port 6 se
rlabel metal1 562 40 591 47 0 A
port 7 se
rlabel metal1 370 47 871 61 0 A
port 8 se
rlabel metal1 370 61 399 69 0 A
port 9 se
rlabel metal1 562 61 591 69 0 A
port 10 se
rlabel metal1 857 61 871 80 0 A
port 11 se
rlabel metal1 850 80 879 109 0 A
port 12 se
rlabel metal1 857 109 871 175 0 A
port 13 se
rlabel metal1 850 175 879 204 0 A
port 14 se
rlabel metal1 130 121 159 150 0 B
port 15 se
rlabel metal1 137 150 151 175 0 B
port 16 se
rlabel metal1 130 175 159 182 0 B
port 17 se
rlabel metal1 274 175 303 182 0 B
port 18 se
rlabel metal1 130 182 303 196 0 B
port 19 se
rlabel metal1 130 196 159 204 0 B
port 20 se
rlabel metal1 274 196 303 204 0 B
port 21 se
<< properties >>
string FIXED_BBOX 0 0 1008 333
<< end >>
