magic
tech sky130A
timestamp 1624703114
<< nwell >>
rect 0 179 432 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 322 67 351 73
rect 322 66 328 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 51 281 66
rect 152 34 184 51
rect 201 34 281 51
rect 152 24 281 34
rect 296 50 328 66
rect 345 66 351 67
rect 345 50 375 66
rect 296 24 375 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 243 375 309
rect 296 226 328 243
rect 345 226 375 243
rect 296 225 375 226
rect 58 220 87 225
rect 322 220 351 225
<< ndiffc >>
rect 64 50 81 67
rect 184 34 201 51
rect 328 50 345 67
<< pdiffc >>
rect 64 226 81 243
rect 184 282 201 299
rect 328 226 345 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 137 209 152 225
rect 281 209 296 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 137 66 152 83
rect 281 66 296 83
rect 137 11 152 24
rect 281 11 296 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 136 91 153 108
rect 280 91 297 108
<< locali >>
rect 0 342 432 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 432 342
rect 0 309 432 325
rect 176 299 209 309
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 320 243 353 251
rect 320 226 328 243
rect 345 226 353 243
rect 320 218 353 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 303 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 92 305 108
rect 297 91 303 92
rect 272 83 303 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 320 67 353 75
rect 56 42 89 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 320 50 328 67
rect 345 50 353 67
rect 320 42 353 50
rect 176 24 209 34
rect 0 9 432 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 432 9
rect 0 -24 432 -9
<< viali >>
rect 16 325 33 342
rect 64 325 81 342
rect 112 325 129 342
rect 160 325 177 342
rect 208 325 225 342
rect 256 325 273 342
rect 304 325 321 342
rect 352 325 369 342
rect 400 325 417 342
rect 184 282 201 299
rect 64 226 81 243
rect 328 226 345 243
rect 136 184 153 201
rect 280 184 297 201
rect 136 91 153 108
rect 280 91 297 108
rect 64 50 81 67
rect 328 50 345 67
rect 16 -9 33 9
rect 64 -9 81 9
rect 112 -9 129 9
rect 160 -9 177 9
rect 208 -9 225 9
rect 256 -9 273 9
rect 304 -9 321 9
rect 352 -9 369 9
rect 400 -9 417 9
<< metal1 >>
rect 0 342 432 357
rect 0 325 16 342
rect 33 325 64 342
rect 81 325 112 342
rect 129 325 160 342
rect 177 325 208 342
rect 225 325 256 342
rect 273 325 304 342
rect 321 325 352 342
rect 369 325 400 342
rect 417 325 432 342
rect 0 309 432 325
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 322 243 351 249
rect 322 226 328 243
rect 345 226 351 243
rect 322 220 351 226
rect 65 73 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 137 114 151 178
rect 281 114 295 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 106 159 108
rect 274 108 303 114
rect 274 106 280 108
rect 153 92 280 106
rect 153 91 159 92
rect 130 85 159 91
rect 274 91 280 92
rect 297 91 303 108
rect 274 85 303 91
rect 329 73 343 220
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 322 67 351 73
rect 322 66 328 67
rect 81 52 328 66
rect 81 50 87 52
rect 58 44 87 50
rect 322 50 328 52
rect 345 50 351 67
rect 322 44 351 50
rect 0 9 432 24
rect 0 -9 16 9
rect 33 -9 64 9
rect 81 -9 112 9
rect 129 -9 160 9
rect 177 -9 208 9
rect 225 -9 256 9
rect 273 -9 304 9
rect 321 -9 352 9
rect 369 -9 400 9
rect 417 -9 432 9
rect 0 -24 432 -9
<< labels >>
rlabel locali 0 309 432 357 0 VDD
port 1 se
rlabel metal1 0 309 432 357 0 VDD
port 2 se
rlabel locali 0 -24 432 24 0 GND
port 3 se
rlabel metal1 0 -24 432 24 0 GND
port 4 se
rlabel metal1 58 44 87 52 0 Y
port 5 se
rlabel metal1 322 44 351 52 0 Y
port 6 se
rlabel metal1 58 52 351 66 0 Y
port 7 se
rlabel metal1 58 66 87 73 0 Y
port 8 se
rlabel metal1 322 66 351 73 0 Y
port 9 se
rlabel metal1 65 73 79 220 0 Y
port 10 se
rlabel metal1 329 73 343 220 0 Y
port 11 se
rlabel metal1 58 220 87 249 0 Y
port 12 se
rlabel metal1 322 220 351 249 0 Y
port 13 se
rlabel metal1 130 85 159 92 0 A
port 14 se
rlabel metal1 274 85 303 92 0 A
port 15 se
rlabel metal1 130 92 303 106 0 A
port 16 se
rlabel metal1 130 106 159 114 0 A
port 17 se
rlabel metal1 274 106 303 114 0 A
port 18 se
rlabel metal1 137 114 151 178 0 A
port 19 se
rlabel metal1 281 114 295 178 0 A
port 20 se
rlabel metal1 130 178 159 207 0 A
port 21 se
rlabel metal1 274 178 303 207 0 A
port 22 se
<< properties >>
string FIXED_BBOX 0 0 432 333
<< end >>
