magic
tech sky130A
timestamp 1624189032
<< nwell >>
rect 0 179 432 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
<< ndiff >>
rect 82 67 111 73
rect 82 66 88 67
rect 58 50 88 66
rect 105 66 111 67
rect 322 67 351 73
rect 322 66 328 67
rect 105 50 137 66
rect 58 24 137 50
rect 152 51 281 66
rect 152 34 184 51
rect 201 34 281 51
rect 152 24 281 34
rect 296 50 328 66
rect 345 66 351 67
rect 345 50 375 66
rect 296 24 375 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 88 243
rect 105 226 137 243
rect 58 225 137 226
rect 152 299 281 309
rect 152 282 184 299
rect 201 282 281 299
rect 152 225 281 282
rect 296 243 375 309
rect 296 226 328 243
rect 345 226 375 243
rect 296 225 375 226
rect 82 220 111 225
rect 322 220 351 225
<< ndiffc >>
rect 88 50 105 67
rect 184 34 201 51
rect 328 50 345 67
<< pdiffc >>
rect 88 226 105 243
rect 184 282 201 299
rect 328 226 345 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 137 209 152 225
rect 281 209 296 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 137 66 152 83
rect 281 66 296 83
rect 137 11 152 24
rect 281 11 296 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 136 91 153 108
rect 280 91 297 108
<< locali >>
rect 176 299 209 307
rect 176 282 184 299
rect 201 282 209 299
rect 176 274 209 282
rect 80 243 113 251
rect 80 226 88 243
rect 105 226 113 243
rect 320 243 353 251
rect 320 226 328 243
rect 345 226 353 243
rect 80 218 111 226
rect 322 218 353 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 128 108 161 116
rect 128 92 136 108
rect 130 91 136 92
rect 153 91 161 108
rect 130 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 80 67 113 75
rect 80 50 88 67
rect 105 50 113 67
rect 322 67 353 75
rect 322 66 328 67
rect 80 42 113 50
rect 176 51 209 59
rect 176 34 184 51
rect 201 34 209 51
rect 320 50 328 66
rect 345 50 353 67
rect 320 42 353 50
rect 176 26 209 34
rect 184 9 201 26
<< viali >>
rect 184 282 201 299
rect 88 226 105 243
rect 328 226 345 243
rect 136 184 153 201
rect 280 184 297 201
rect 136 91 153 108
rect 280 91 297 108
rect 88 50 105 67
rect 328 50 345 67
rect 184 -9 201 9
<< metal1 >>
rect 0 309 432 357
rect 178 299 207 309
rect 178 282 184 299
rect 201 282 207 299
rect 178 276 207 282
rect 82 243 111 249
rect 82 226 88 243
rect 105 241 111 243
rect 322 243 351 249
rect 322 241 328 243
rect 105 227 328 241
rect 105 226 111 227
rect 82 220 111 226
rect 322 226 328 227
rect 345 226 351 243
rect 322 220 351 226
rect 89 73 103 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 137 114 151 178
rect 281 114 295 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 106 159 108
rect 274 108 303 114
rect 274 106 280 108
rect 153 92 280 106
rect 153 91 159 92
rect 130 85 159 91
rect 274 91 280 92
rect 297 91 303 108
rect 274 85 303 91
rect 329 73 343 220
rect 82 67 111 73
rect 82 50 88 67
rect 105 50 111 67
rect 82 44 111 50
rect 322 67 351 73
rect 322 50 328 67
rect 345 50 351 67
rect 322 44 351 50
rect 0 9 432 24
rect 0 -9 184 9
rect 201 -9 432 9
rect 0 -24 432 -9
<< labels >>
rlabel metal1 0 309 432 357 0 VDD
port 1 se
rlabel metal1 0 -24 432 24 0 GND
port 2 se
rlabel metal1 82 44 111 73 0 Y
port 3 se
rlabel metal1 322 44 351 73 0 Y
port 4 se
rlabel metal1 89 73 103 220 0 Y
port 5 se
rlabel metal1 329 73 343 220 0 Y
port 6 se
rlabel metal1 82 220 111 227 0 Y
port 7 se
rlabel metal1 322 220 351 227 0 Y
port 8 se
rlabel metal1 82 227 351 241 0 Y
port 9 se
rlabel metal1 82 241 111 249 0 Y
port 10 se
rlabel metal1 322 241 351 249 0 Y
port 11 se
rlabel metal1 130 85 159 92 0 A
port 12 se
rlabel metal1 274 85 303 92 0 A
port 13 se
rlabel metal1 130 92 303 106 0 A
port 14 se
rlabel metal1 130 106 159 114 0 A
port 15 se
rlabel metal1 274 106 303 114 0 A
port 16 se
rlabel metal1 137 114 151 178 0 A
port 17 se
rlabel metal1 281 114 295 178 0 A
port 18 se
rlabel metal1 130 178 159 207 0 A
port 19 se
rlabel metal1 274 178 303 207 0 A
port 20 se
<< properties >>
string FIXED_BBOX 0 0 432 333
<< end >>
