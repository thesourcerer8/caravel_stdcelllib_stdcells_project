VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 0.580 2.970 0.870 3.090 ;
        RECT 0.580 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.870 2.970 ;
        RECT 0.580 2.740 0.870 2.800 ;
        RECT 3.220 2.970 3.510 3.090 ;
        RECT 3.220 2.800 3.280 2.970 ;
        RECT 3.450 2.800 3.510 2.970 ;
        RECT 3.220 2.740 3.510 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 0.560 2.970 0.890 3.090 ;
        RECT 0.560 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.890 2.970 ;
        RECT 0.560 2.720 0.890 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.220 0.670 3.510 0.730 ;
        RECT 3.220 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.510 0.670 ;
        RECT 3.220 0.440 3.510 0.500 ;
        RECT 3.290 0.240 3.430 0.440 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.200 4.950 2.490 ;
        RECT 4.730 0.730 4.870 2.200 ;
        RECT 4.660 0.440 4.950 0.730 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.390 3.030 1.680 ;
        RECT 2.810 1.140 2.950 1.390 ;
        RECT 2.740 0.850 3.030 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 3.200 2.970 3.530 3.050 ;
        RECT 3.200 2.800 3.280 2.970 ;
        RECT 3.450 2.800 3.530 2.970 ;
        RECT 3.200 2.720 3.530 2.800 ;
        RECT 1.760 2.430 2.090 2.510 ;
        RECT 1.760 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.090 2.430 ;
        RECT 4.640 2.430 4.970 2.510 ;
        RECT 4.640 2.260 4.720 2.430 ;
        RECT 4.890 2.260 4.970 2.430 ;
        RECT 1.780 2.180 2.090 2.260 ;
        RECT 4.660 2.180 4.970 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 2.800 1.620 2.970 1.760 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.920 1.360 1.080 ;
        RECT 1.300 0.910 1.360 0.920 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.300 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.920 4.490 1.080 ;
        RECT 4.410 0.910 4.470 0.920 ;
        RECT 4.160 0.830 4.470 0.910 ;
        RECT 0.800 0.670 1.130 0.750 ;
        RECT 0.800 0.500 0.880 0.670 ;
        RECT 1.050 0.500 1.130 0.670 ;
        RECT 3.220 0.670 3.530 0.750 ;
        RECT 3.220 0.660 3.280 0.670 ;
        RECT 0.800 0.420 1.130 0.500 ;
        RECT 3.200 0.500 3.280 0.660 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
        RECT 4.640 0.670 4.970 0.750 ;
        RECT 4.640 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
      LAYER met1 ;
        RECT 1.780 2.430 2.070 2.490 ;
        RECT 1.780 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.070 2.430 ;
        RECT 1.780 2.200 2.070 2.260 ;
        RECT 1.850 2.000 1.990 2.200 ;
        RECT 4.180 2.010 4.470 2.070 ;
        RECT 4.180 2.000 4.240 2.010 ;
        RECT 1.850 1.860 4.240 2.000 ;
        RECT 0.820 0.670 1.110 0.730 ;
        RECT 0.820 0.500 0.880 0.670 ;
        RECT 1.050 0.660 1.110 0.670 ;
        RECT 1.850 0.660 1.990 1.860 ;
        RECT 4.180 1.840 4.240 1.860 ;
        RECT 4.410 1.840 4.470 2.010 ;
        RECT 4.180 1.780 4.470 1.840 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 4.180 1.080 4.470 1.140 ;
        RECT 4.180 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.470 1.080 ;
        RECT 4.180 0.850 4.470 0.910 ;
        RECT 1.050 0.520 1.990 0.660 ;
        RECT 1.050 0.500 1.110 0.520 ;
        RECT 0.820 0.440 1.110 0.500 ;
  END
END AND2X2
END LIBRARY

