magic
tech sky130A
timestamp 1623602976
<< nwell >>
rect 0 179 864 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
<< ndiff >>
rect 58 66 87 69
rect 514 66 543 69
rect 58 63 137 66
rect 58 46 64 63
rect 81 46 137 63
rect 58 24 137 46
rect 152 36 281 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 281 36
rect 296 24 425 66
rect 440 63 569 66
rect 440 46 520 63
rect 537 46 569 63
rect 440 24 569 46
rect 584 24 713 66
rect 728 36 807 66
rect 728 24 760 36
rect 201 19 207 24
rect 178 13 207 19
rect 754 19 760 24
rect 777 24 807 36
rect 777 19 783 24
rect 754 13 783 19
<< pdiff >>
rect 178 309 207 312
rect 754 309 783 312
rect 58 238 137 309
rect 58 221 64 238
rect 81 225 137 238
rect 152 306 281 309
rect 152 289 184 306
rect 201 289 281 306
rect 152 225 281 289
rect 296 225 425 309
rect 440 238 569 309
rect 440 225 520 238
rect 81 221 87 225
rect 58 215 87 221
rect 514 221 520 225
rect 537 225 569 238
rect 584 225 713 309
rect 728 306 807 309
rect 728 289 760 306
rect 777 289 807 306
rect 728 225 807 289
rect 537 221 543 225
rect 514 215 543 221
<< ndiffc >>
rect 64 46 81 63
rect 184 19 201 36
rect 520 46 537 63
rect 760 19 777 36
<< pdiffc >>
rect 64 221 81 238
rect 184 289 201 306
rect 520 221 537 238
rect 760 289 777 306
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 425 309 440 330
rect 569 309 584 330
rect 713 309 728 330
rect 137 206 152 225
rect 281 206 296 225
rect 425 206 440 225
rect 569 206 584 225
rect 713 206 728 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 416 173 449 181
rect 560 198 593 206
rect 560 181 568 198
rect 585 181 593 198
rect 560 173 593 181
rect 704 198 737 206
rect 704 181 712 198
rect 729 181 737 198
rect 704 173 737 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 560 103 593 111
rect 560 86 568 103
rect 585 86 593 103
rect 560 78 593 86
rect 704 103 737 111
rect 704 86 712 103
rect 729 86 737 103
rect 704 78 737 86
rect 137 66 152 78
rect 281 66 296 78
rect 425 66 440 78
rect 569 66 584 78
rect 713 66 728 78
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 424 181 441 198
rect 568 181 585 198
rect 712 181 729 198
rect 136 86 153 103
rect 280 86 297 103
rect 424 86 441 103
rect 568 86 585 103
rect 712 86 729 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 752 306 785 314
rect 752 289 760 306
rect 777 289 785 306
rect 752 281 785 289
rect 56 238 89 246
rect 56 221 64 238
rect 81 221 89 238
rect 56 213 89 221
rect 512 238 545 246
rect 512 221 520 238
rect 537 221 545 238
rect 512 213 545 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 416 198 449 206
rect 416 181 424 198
rect 441 181 449 198
rect 562 198 593 206
rect 562 196 568 198
rect 416 173 449 181
rect 560 181 568 196
rect 585 181 593 198
rect 560 173 593 181
rect 704 198 737 206
rect 704 181 712 198
rect 729 181 737 198
rect 704 173 737 181
rect 136 111 153 173
rect 280 144 297 173
rect 280 111 297 127
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 416 103 449 111
rect 416 86 424 103
rect 441 86 449 103
rect 416 78 449 86
rect 520 71 537 127
rect 560 103 593 111
rect 560 88 568 103
rect 562 86 568 88
rect 585 86 593 103
rect 562 78 593 86
rect 704 103 737 111
rect 704 86 712 103
rect 729 86 737 103
rect 704 78 737 86
rect 56 63 89 71
rect 56 46 64 63
rect 81 46 89 63
rect 56 38 89 46
rect 512 63 545 71
rect 512 46 520 63
rect 537 46 545 63
rect 176 36 209 44
rect 512 38 545 46
rect 176 19 184 36
rect 201 19 209 36
rect 176 11 209 19
rect 752 36 785 44
rect 752 19 760 36
rect 777 19 785 36
rect 752 11 785 19
<< viali >>
rect 184 289 201 306
rect 760 289 777 306
rect 64 221 81 238
rect 520 221 537 238
rect 424 181 441 198
rect 568 181 585 198
rect 712 181 729 198
rect 280 127 297 144
rect 520 127 537 144
rect 136 86 153 103
rect 424 86 441 103
rect 568 86 585 103
rect 712 86 729 103
rect 64 46 81 63
rect 184 19 201 36
rect 760 19 777 36
<< metal1 >>
rect 0 309 864 357
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 754 306 783 309
rect 754 289 760 306
rect 777 289 783 306
rect 754 283 783 289
rect 58 238 87 244
rect 58 221 64 238
rect 81 221 87 238
rect 58 215 87 221
rect 514 238 543 244
rect 514 221 520 238
rect 537 221 543 238
rect 514 215 543 221
rect 65 196 79 215
rect 418 198 447 204
rect 418 196 424 198
rect 65 182 424 196
rect 65 69 79 182
rect 418 181 424 182
rect 441 196 447 198
rect 441 182 487 196
rect 441 181 447 182
rect 418 175 447 181
rect 274 144 303 150
rect 274 127 280 144
rect 297 127 303 144
rect 274 121 303 127
rect 130 103 159 109
rect 130 86 136 103
rect 153 102 159 103
rect 418 103 447 109
rect 418 102 424 103
rect 153 88 424 102
rect 153 86 159 88
rect 130 80 159 86
rect 418 86 424 88
rect 441 86 447 103
rect 473 102 487 182
rect 521 150 535 215
rect 562 198 591 204
rect 562 181 568 198
rect 585 196 591 198
rect 706 198 735 204
rect 585 182 631 196
rect 585 181 591 182
rect 562 175 591 181
rect 514 144 543 150
rect 514 127 520 144
rect 537 127 543 144
rect 514 121 543 127
rect 562 103 591 109
rect 562 102 568 103
rect 473 88 568 102
rect 418 80 447 86
rect 562 86 568 88
rect 585 86 591 103
rect 562 80 591 86
rect 58 63 87 69
rect 58 46 64 63
rect 81 46 87 63
rect 425 61 439 80
rect 617 61 631 182
rect 706 181 712 198
rect 729 181 735 198
rect 706 175 735 181
rect 713 109 727 175
rect 706 103 735 109
rect 706 86 712 103
rect 729 86 735 103
rect 706 80 735 86
rect 425 47 631 61
rect 58 40 87 46
rect 178 36 207 42
rect 178 24 184 36
rect 0 19 184 24
rect 201 24 207 36
rect 754 36 783 42
rect 754 24 760 36
rect 201 19 760 24
rect 777 24 783 36
rect 777 19 864 24
rect 0 -24 864 19
<< labels >>
rlabel metal1 0 309 864 357 0 VDD
port 1 se
rlabel metal1 0 -24 864 24 0 GND
port 2 se
rlabel metal1 514 121 543 150 0 Y
port 3 se
rlabel metal1 521 150 535 215 0 Y
port 4 se
rlabel metal1 514 215 543 244 0 Y
port 5 se
rlabel metal1 425 47 631 61 0 S
port 6 se
rlabel metal1 425 61 439 80 0 S
port 7 se
rlabel metal1 130 80 159 88 0 S
port 8 se
rlabel metal1 418 80 447 88 0 S
port 9 se
rlabel metal1 130 88 447 102 0 S
port 10 se
rlabel metal1 130 102 159 109 0 S
port 11 se
rlabel metal1 418 102 447 109 0 S
port 12 se
rlabel metal1 562 175 591 182 0 S
port 13 se
rlabel metal1 617 61 631 182 0 S
port 14 se
rlabel metal1 562 182 631 196 0 S
port 15 se
rlabel metal1 562 196 591 204 0 S
port 16 se
rlabel metal1 706 80 735 109 0 B
port 17 se
rlabel metal1 713 109 727 175 0 B
port 18 se
rlabel metal1 706 175 735 204 0 B
port 19 se
rlabel metal1 274 121 303 150 0 A
port 20 se
<< properties >>
string FIXED_BBOX 0 0 864 333
<< end >>
