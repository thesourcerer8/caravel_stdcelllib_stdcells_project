magic
tech sky130A
magscale 1 2
timestamp 1623617396
<< locali >>
rect 47551 43566 47585 43680
rect 37087 36092 37121 36206
rect 8767 27508 8801 27548
rect 8513 27474 8801 27508
rect 8383 19442 8417 19778
rect 8767 18406 8801 18446
rect 8767 18372 9055 18406
rect 8095 16926 8129 17188
rect 7745 11786 7903 11820
rect 28927 7528 28961 7642
rect 39487 6862 39521 7050
rect 45439 6196 45473 6532
rect 7999 5530 8033 5644
<< viali >>
rect 9919 57000 9953 57034
rect 13951 57000 13985 57034
rect 32671 57000 32705 57034
rect 1951 56926 1985 56960
rect 2815 56926 2849 56960
rect 5311 56926 5345 56960
rect 5791 56926 5825 56960
rect 7423 56926 7457 56960
rect 8095 56926 8129 56960
rect 11455 56926 11489 56960
rect 13183 56926 13217 56960
rect 15103 56926 15137 56960
rect 16351 56926 16385 56960
rect 18175 56926 18209 56960
rect 19519 56926 19553 56960
rect 21055 56926 21089 56960
rect 22015 56926 22049 56960
rect 24223 56926 24257 56960
rect 25951 56926 25985 56960
rect 27391 56926 27425 56960
rect 29023 56926 29057 56960
rect 30079 56926 30113 56960
rect 31711 56926 31745 56960
rect 34303 56926 34337 56960
rect 34879 56926 34913 56960
rect 38047 56926 38081 56960
rect 41983 56926 42017 56960
rect 44671 56926 44705 56960
rect 47551 56926 47585 56960
rect 53887 56926 53921 56960
rect 1759 56852 1793 56886
rect 2623 56852 2657 56886
rect 5119 56852 5153 56886
rect 7231 56852 7265 56886
rect 11263 56852 11297 56886
rect 12991 56852 13025 56886
rect 14047 56852 14081 56886
rect 16159 56852 16193 56886
rect 17983 56852 18017 56886
rect 19327 56852 19361 56886
rect 20863 56852 20897 56886
rect 24031 56852 24065 56886
rect 27199 56852 27233 56886
rect 28831 56852 28865 56886
rect 32383 56852 32417 56886
rect 32575 56852 32609 56886
rect 34111 56852 34145 56886
rect 36991 56852 37025 56886
rect 40063 56852 40097 56886
rect 40735 56852 40769 56886
rect 43231 56852 43265 56886
rect 46303 56852 46337 56886
rect 48991 56852 49025 56886
rect 51103 56852 51137 56886
rect 53119 56852 53153 56886
rect 55807 56852 55841 56886
rect 57055 56852 57089 56886
rect 9823 56704 9857 56738
rect 36703 56704 36737 56738
rect 39775 56704 39809 56738
rect 40447 56704 40481 56738
rect 40831 56704 40865 56738
rect 42943 56704 42977 56738
rect 46015 56704 46049 56738
rect 48703 56704 48737 56738
rect 50815 56704 50849 56738
rect 52831 56704 52865 56738
rect 55519 56704 55553 56738
rect 56767 56704 56801 56738
rect 1663 56482 1697 56516
rect 2431 56482 2465 56516
rect 3199 56482 3233 56516
rect 4447 56482 4481 56516
rect 5503 56482 5537 56516
rect 6271 56482 6305 56516
rect 7135 56482 7169 56516
rect 8479 56482 8513 56516
rect 10399 56482 10433 56516
rect 11071 56482 11105 56516
rect 11839 56482 11873 56516
rect 12607 56482 12641 56516
rect 13471 56482 13505 56516
rect 15007 56482 15041 56516
rect 17215 56482 17249 56516
rect 18175 56482 18209 56516
rect 19039 56482 19073 56516
rect 21343 56482 21377 56516
rect 22111 56482 22145 56516
rect 22879 56482 22913 56516
rect 24415 56482 24449 56516
rect 26047 56482 26081 56516
rect 26911 56482 26945 56516
rect 27775 56482 27809 56516
rect 28543 56482 28577 56516
rect 29695 56482 29729 56516
rect 30847 56482 30881 56516
rect 32383 56482 32417 56516
rect 33919 56482 33953 56516
rect 34687 56482 34721 56516
rect 36991 56482 37025 56516
rect 37663 56482 37697 56516
rect 38719 56482 38753 56516
rect 40159 56482 40193 56516
rect 41887 56482 41921 56516
rect 42751 56482 42785 56516
rect 43519 56482 43553 56516
rect 44191 56482 44225 56516
rect 45055 56482 45089 56516
rect 46783 56482 46817 56516
rect 48127 56482 48161 56516
rect 49759 56482 49793 56516
rect 50527 56482 50561 56516
rect 52927 56482 52961 56516
rect 53791 56482 53825 56516
rect 54559 56482 54593 56516
rect 55327 56482 55361 56516
rect 55999 56482 56033 56516
rect 6943 56334 6977 56368
rect 7231 56334 7265 56368
rect 37471 56334 37505 56368
rect 37759 56334 37793 56368
rect 45151 56334 45185 56368
rect 52063 56334 52097 56368
rect 56095 56334 56129 56368
rect 10111 56260 10145 56294
rect 10303 56260 10337 56294
rect 13567 56260 13601 56294
rect 25855 56260 25889 56294
rect 26143 56260 26177 56294
rect 38815 56260 38849 56294
rect 44287 56260 44321 56294
rect 46975 56260 47009 56294
rect 50623 56260 50657 56294
rect 57823 56260 57857 56294
rect 1759 56186 1793 56220
rect 2527 56186 2561 56220
rect 3007 56186 3041 56220
rect 3295 56186 3329 56220
rect 4255 56186 4289 56220
rect 4543 56186 4577 56220
rect 5599 56186 5633 56220
rect 6367 56186 6401 56220
rect 8575 56186 8609 56220
rect 10783 56186 10817 56220
rect 11167 56186 11201 56220
rect 11935 56186 11969 56220
rect 12415 56186 12449 56220
rect 12703 56186 12737 56220
rect 15103 56186 15137 56220
rect 15583 56186 15617 56220
rect 15775 56186 15809 56220
rect 15871 56186 15905 56220
rect 16831 56186 16865 56220
rect 17119 56186 17153 56220
rect 17983 56186 18017 56220
rect 18271 56186 18305 56220
rect 18751 56186 18785 56220
rect 18943 56186 18977 56220
rect 19999 56186 20033 56220
rect 20287 56186 20321 56220
rect 20383 56186 20417 56220
rect 21055 56186 21089 56220
rect 21439 56186 21473 56220
rect 21823 56186 21857 56220
rect 22207 56186 22241 56220
rect 22975 56186 23009 56220
rect 24127 56186 24161 56220
rect 24319 56186 24353 56220
rect 26527 56186 26561 56220
rect 26815 56186 26849 56220
rect 27487 56186 27521 56220
rect 27679 56186 27713 56220
rect 28159 56186 28193 56220
rect 28447 56186 28481 56220
rect 29407 56186 29441 56220
rect 29599 56186 29633 56220
rect 30943 56186 30977 56220
rect 31327 56186 31361 56220
rect 31615 56186 31649 56220
rect 31711 56186 31745 56220
rect 32191 56186 32225 56220
rect 32479 56186 32513 56220
rect 32863 56186 32897 56220
rect 33151 56186 33185 56220
rect 33247 56186 33281 56220
rect 34015 56186 34049 56220
rect 34783 56186 34817 56220
rect 35839 56186 35873 56220
rect 36127 56186 36161 56220
rect 36223 56186 36257 56220
rect 36607 56186 36641 56220
rect 36895 56186 36929 56220
rect 40255 56186 40289 56220
rect 41983 56186 42017 56220
rect 42367 56186 42401 56220
rect 42655 56186 42689 56220
rect 43231 56186 43265 56220
rect 43423 56186 43457 56220
rect 46495 56186 46529 56220
rect 46687 56186 46721 56220
rect 48223 56186 48257 56220
rect 48703 56186 48737 56220
rect 48895 56186 48929 56220
rect 48991 56186 49025 56220
rect 49855 56186 49889 56220
rect 51967 56186 52001 56220
rect 53023 56186 53057 56220
rect 53407 56186 53441 56220
rect 53695 56186 53729 56220
rect 54271 56186 54305 56220
rect 54463 56186 54497 56220
rect 55039 56186 55073 56220
rect 55231 56186 55265 56220
rect 55519 56186 55553 56220
rect 17983 55742 18017 55776
rect 18271 55742 18305 55776
rect 1663 55668 1697 55702
rect 4447 55668 4481 55702
rect 7615 55668 7649 55702
rect 9343 55668 9377 55702
rect 13951 55668 13985 55702
rect 20287 55668 20321 55702
rect 23551 55668 23585 55702
rect 25087 55668 25121 55702
rect 39295 55668 39329 55702
rect 40831 55668 40865 55702
rect 45631 55668 45665 55702
rect 47167 55668 47201 55702
rect 51967 55668 52001 55702
rect 56575 55668 56609 55702
rect 57727 55668 57761 55702
rect 21439 55594 21473 55628
rect 54271 55594 54305 55628
rect 54463 55594 54497 55628
rect 1759 55520 1793 55554
rect 4255 55520 4289 55554
rect 4543 55520 4577 55554
rect 7711 55520 7745 55554
rect 8191 55520 8225 55554
rect 8479 55520 8513 55554
rect 9055 55520 9089 55554
rect 9247 55520 9281 55554
rect 13759 55520 13793 55554
rect 14047 55520 14081 55554
rect 20383 55520 20417 55554
rect 23263 55520 23297 55554
rect 23455 55520 23489 55554
rect 24991 55520 25025 55554
rect 28927 55520 28961 55554
rect 30175 55520 30209 55554
rect 39199 55520 39233 55554
rect 40927 55520 40961 55554
rect 45535 55520 45569 55554
rect 47071 55520 47105 55554
rect 50527 55520 50561 55554
rect 51871 55520 51905 55554
rect 55807 55520 55841 55554
rect 56383 55520 56417 55554
rect 56671 55520 56705 55554
rect 57439 55520 57473 55554
rect 57631 55520 57665 55554
rect 1951 55372 1985 55406
rect 24703 55372 24737 55406
rect 28831 55372 28865 55406
rect 29791 55372 29825 55406
rect 38911 55372 38945 55406
rect 45247 55372 45281 55406
rect 46783 55372 46817 55406
rect 50431 55372 50465 55406
rect 51583 55372 51617 55406
rect 55615 55372 55649 55406
rect 26719 55150 26753 55184
rect 57823 55150 57857 55184
rect 54463 55002 54497 55036
rect 36703 54928 36737 54962
rect 36799 54928 36833 54962
rect 57919 54854 57953 54888
rect 22111 54706 22145 54740
rect 46591 54706 46625 54740
rect 46783 54706 46817 54740
rect 57919 54336 57953 54370
rect 30847 54188 30881 54222
rect 31135 54188 31169 54222
rect 42367 54188 42401 54222
rect 44959 54188 44993 54222
rect 45247 54188 45281 54222
rect 57823 54188 57857 54222
rect 42175 54114 42209 54148
rect 2431 54040 2465 54074
rect 57631 54040 57665 54074
rect 57919 53818 57953 53852
rect 7903 53522 7937 53556
rect 8191 53522 8225 53556
rect 57823 53522 57857 53556
rect 5215 53374 5249 53408
rect 5503 53374 5537 53408
rect 57631 53374 57665 53408
rect 12415 52856 12449 52890
rect 12607 52856 12641 52890
rect 23551 52856 23585 52890
rect 40543 52856 40577 52890
rect 40735 52856 40769 52890
rect 23455 52708 23489 52742
rect 32287 52190 32321 52224
rect 41119 51524 41153 51558
rect 41311 51524 41345 51558
rect 52735 51006 52769 51040
rect 51871 50858 51905 50892
rect 9439 50710 9473 50744
rect 9823 50710 9857 50744
rect 10687 50710 10721 50744
rect 10975 50710 11009 50744
rect 54943 50488 54977 50522
rect 10303 50414 10337 50448
rect 10015 50340 10049 50374
rect 4255 49378 4289 49412
rect 4543 49378 4577 49412
rect 33247 49378 33281 49412
rect 33439 49378 33473 49412
rect 44191 49378 44225 49412
rect 44383 49378 44417 49412
rect 27967 48860 28001 48894
rect 28255 48860 28289 48894
rect 2431 48046 2465 48080
rect 2719 48046 2753 48080
rect 41119 48046 41153 48080
rect 41311 48046 41345 48080
rect 8095 47528 8129 47562
rect 8383 47528 8417 47562
rect 49183 47454 49217 47488
rect 52735 47010 52769 47044
rect 36415 46714 36449 46748
rect 36799 46714 36833 46748
rect 17983 46196 18017 46230
rect 17695 46122 17729 46156
rect 12511 45382 12545 45416
rect 12607 45382 12641 45416
rect 48031 45382 48065 45416
rect 48799 45382 48833 45416
rect 48991 45382 49025 45416
rect 55807 45382 55841 45416
rect 55999 45382 56033 45416
rect 12127 44864 12161 44898
rect 12415 44864 12449 44898
rect 4255 44050 4289 44084
rect 4543 44050 4577 44084
rect 46399 44050 46433 44084
rect 46591 44050 46625 44084
rect 52063 44050 52097 44084
rect 52159 44050 52193 44084
rect 46303 43754 46337 43788
rect 46591 43754 46625 43788
rect 47551 43680 47585 43714
rect 17407 43532 17441 43566
rect 17695 43532 17729 43566
rect 47551 43532 47585 43566
rect 47743 43532 47777 43566
rect 47839 43532 47873 43566
rect 51295 43532 51329 43566
rect 51103 43458 51137 43492
rect 16159 42718 16193 42752
rect 16447 42718 16481 42752
rect 20095 42718 20129 42752
rect 20191 42718 20225 42752
rect 22687 42718 22721 42752
rect 22879 42718 22913 42752
rect 52543 42718 52577 42752
rect 52735 42718 52769 42752
rect 3583 42200 3617 42234
rect 29983 42200 30017 42234
rect 45343 42200 45377 42234
rect 29791 42052 29825 42086
rect 45247 42052 45281 42086
rect 33823 40868 33857 40902
rect 49759 40868 49793 40902
rect 49951 40868 49985 40902
rect 33631 40720 33665 40754
rect 57727 40720 57761 40754
rect 16543 40498 16577 40532
rect 17023 40054 17057 40088
rect 17215 40054 17249 40088
rect 23359 40054 23393 40088
rect 23551 40054 23585 40088
rect 47263 40054 47297 40088
rect 47455 40054 47489 40088
rect 47935 39536 47969 39570
rect 48223 39536 48257 39570
rect 51295 39536 51329 39570
rect 51583 39536 51617 39570
rect 34303 38870 34337 38904
rect 32095 38722 32129 38756
rect 34591 38722 34625 38756
rect 17695 38204 17729 38238
rect 36895 38204 36929 38238
rect 51679 37464 51713 37498
rect 1855 37390 1889 37424
rect 2047 37390 2081 37424
rect 5503 37390 5537 37424
rect 47455 37390 47489 37424
rect 51871 37390 51905 37424
rect 24991 37094 25025 37128
rect 6943 37020 6977 37054
rect 27967 36872 28001 36906
rect 28255 36872 28289 36906
rect 56383 36872 56417 36906
rect 24127 36798 24161 36832
rect 33439 36280 33473 36314
rect 33631 36280 33665 36314
rect 22015 36206 22049 36240
rect 37087 36206 37121 36240
rect 25567 36132 25601 36166
rect 25855 36132 25889 36166
rect 21247 36058 21281 36092
rect 21535 36058 21569 36092
rect 36703 36058 36737 36092
rect 36991 36058 37025 36092
rect 37087 36058 37121 36092
rect 50623 36058 50657 36092
rect 41503 35688 41537 35722
rect 46399 35540 46433 35574
rect 46687 35540 46721 35574
rect 12607 34800 12641 34834
rect 12895 34800 12929 34834
rect 41503 34726 41537 34760
rect 41695 34726 41729 34760
rect 17887 34356 17921 34390
rect 13855 34282 13889 34316
rect 14143 34282 14177 34316
rect 9919 34208 9953 34242
rect 21439 34208 21473 34242
rect 21151 34134 21185 34168
rect 56191 33690 56225 33724
rect 42175 33616 42209 33650
rect 42367 33616 42401 33650
rect 29311 33394 29345 33428
rect 29503 33394 29537 33428
rect 34687 33394 34721 33428
rect 37951 33394 37985 33428
rect 38239 33394 38273 33428
rect 55519 33394 55553 33428
rect 37663 33172 37697 33206
rect 44959 33098 44993 33132
rect 29407 32876 29441 32910
rect 29215 32728 29249 32762
rect 2335 32062 2369 32096
rect 6655 32062 6689 32096
rect 41311 30878 41345 30912
rect 11743 30804 11777 30838
rect 6655 30730 6689 30764
rect 28159 30730 28193 30764
rect 28351 30360 28385 30394
rect 7039 30286 7073 30320
rect 32191 30286 32225 30320
rect 7327 30212 7361 30246
rect 14815 29546 14849 29580
rect 15103 29546 15137 29580
rect 12991 29472 13025 29506
rect 1759 29028 1793 29062
rect 2047 29028 2081 29062
rect 44959 28880 44993 28914
rect 50335 28880 50369 28914
rect 22399 28066 22433 28100
rect 22591 28066 22625 28100
rect 8767 27548 8801 27582
rect 16255 27548 16289 27582
rect 22975 27548 23009 27582
rect 8479 27474 8513 27508
rect 33535 26216 33569 26250
rect 36511 26068 36545 26102
rect 36799 26068 36833 26102
rect 2239 24144 2273 24178
rect 2527 24144 2561 24178
rect 13375 24070 13409 24104
rect 36703 24070 36737 24104
rect 36895 24070 36929 24104
rect 44095 23552 44129 23586
rect 8095 22738 8129 22772
rect 28543 22738 28577 22772
rect 2623 22220 2657 22254
rect 31135 21850 31169 21884
rect 31423 21850 31457 21884
rect 32287 21406 32321 21440
rect 58015 21406 58049 21440
rect 43711 21036 43745 21070
rect 43903 21036 43937 21070
rect 41407 20962 41441 20996
rect 7135 20888 7169 20922
rect 34399 20888 34433 20922
rect 7615 20740 7649 20774
rect 9439 20518 9473 20552
rect 16255 20518 16289 20552
rect 16447 20370 16481 20404
rect 44575 20370 44609 20404
rect 44863 20370 44897 20404
rect 9631 20296 9665 20330
rect 10591 20074 10625 20108
rect 18847 20074 18881 20108
rect 42751 20074 42785 20108
rect 47167 20074 47201 20108
rect 8383 19778 8417 19812
rect 45919 19556 45953 19590
rect 52927 19556 52961 19590
rect 54751 19556 54785 19590
rect 7615 19408 7649 19442
rect 8383 19408 8417 19442
rect 36127 18890 36161 18924
rect 36319 18890 36353 18924
rect 4543 18816 4577 18850
rect 57343 18816 57377 18850
rect 15103 18742 15137 18776
rect 39967 18742 40001 18776
rect 7615 18446 7649 18480
rect 8767 18446 8801 18480
rect 9055 18372 9089 18406
rect 24031 18224 24065 18258
rect 44095 18224 44129 18258
rect 44671 18224 44705 18258
rect 9439 18150 9473 18184
rect 9727 18150 9761 18184
rect 44479 18076 44513 18110
rect 46495 17558 46529 17592
rect 46687 17558 46721 17592
rect 57343 17484 57377 17518
rect 7423 17410 7457 17444
rect 8095 17188 8129 17222
rect 8095 16892 8129 16926
rect 7615 16744 7649 16778
rect 2335 16522 2369 16556
rect 2623 16522 2657 16556
rect 54175 16226 54209 16260
rect 3871 15856 3905 15890
rect 8863 15856 8897 15890
rect 16159 15856 16193 15890
rect 26815 15856 26849 15890
rect 50143 15856 50177 15890
rect 7615 15412 7649 15446
rect 2719 14894 2753 14928
rect 2431 14820 2465 14854
rect 25663 14746 25697 14780
rect 9631 14524 9665 14558
rect 14623 14524 14657 14558
rect 49855 14450 49889 14484
rect 56383 14450 56417 14484
rect 27871 14376 27905 14410
rect 28063 14376 28097 14410
rect 7615 14080 7649 14114
rect 25279 13858 25313 13892
rect 25471 13710 25505 13744
rect 57535 13488 57569 13522
rect 54463 13414 54497 13448
rect 56671 13192 56705 13226
rect 56767 13192 56801 13226
rect 7615 13118 7649 13152
rect 57343 12526 57377 12560
rect 57631 12378 57665 12412
rect 57919 12378 57953 12412
rect 57727 12230 57761 12264
rect 37567 12082 37601 12116
rect 56191 11860 56225 11894
rect 7615 11786 7649 11820
rect 7711 11786 7745 11820
rect 7903 11786 7937 11820
rect 10879 11786 10913 11820
rect 34111 11786 34145 11820
rect 34399 11786 34433 11820
rect 56479 11712 56513 11746
rect 56575 11712 56609 11746
rect 57247 11712 57281 11746
rect 25087 11638 25121 11672
rect 57343 11638 57377 11672
rect 44287 11564 44321 11598
rect 5215 11194 5249 11228
rect 56959 11194 56993 11228
rect 5407 11046 5441 11080
rect 57247 11046 57281 11080
rect 57535 11046 57569 11080
rect 48415 10972 48449 11006
rect 56095 10972 56129 11006
rect 34591 10898 34625 10932
rect 34879 10898 34913 10932
rect 55999 10898 56033 10932
rect 57343 10898 57377 10932
rect 42655 10750 42689 10784
rect 4639 10528 4673 10562
rect 55615 10528 55649 10562
rect 56095 10528 56129 10562
rect 55807 10380 55841 10414
rect 57439 10380 57473 10414
rect 46111 10306 46145 10340
rect 56287 10306 56321 10340
rect 56575 10306 56609 10340
rect 38815 10232 38849 10266
rect 55039 10232 55073 10266
rect 57055 10232 57089 10266
rect 57343 10232 57377 10266
rect 54751 10158 54785 10192
rect 7615 10084 7649 10118
rect 55135 10084 55169 10118
rect 55903 10084 55937 10118
rect 56671 10084 56705 10118
rect 54175 9862 54209 9896
rect 54655 9862 54689 9896
rect 55615 9862 55649 9896
rect 54367 9714 54401 9748
rect 55999 9714 56033 9748
rect 57631 9640 57665 9674
rect 54463 9566 54497 9600
rect 55135 9566 55169 9600
rect 55231 9566 55265 9600
rect 55903 9566 55937 9600
rect 5695 9492 5729 9526
rect 28639 9418 28673 9452
rect 36799 9418 36833 9452
rect 54847 9418 54881 9452
rect 12031 9196 12065 9230
rect 12415 9196 12449 9230
rect 7615 9122 7649 9156
rect 9631 9122 9665 9156
rect 9919 9122 9953 9156
rect 55039 9122 55073 9156
rect 53407 9048 53441 9082
rect 55327 9048 55361 9082
rect 54271 8974 54305 9008
rect 54559 8974 54593 9008
rect 56575 8974 56609 9008
rect 57247 8974 57281 9008
rect 46303 8900 46337 8934
rect 51295 8752 51329 8786
rect 51487 8752 51521 8786
rect 53311 8752 53345 8786
rect 54655 8752 54689 8786
rect 55423 8752 55457 8786
rect 12895 8530 12929 8564
rect 15967 8530 16001 8564
rect 48607 8530 48641 8564
rect 52159 8530 52193 8564
rect 52927 8530 52961 8564
rect 1759 8382 1793 8416
rect 2239 8382 2273 8416
rect 2431 8382 2465 8416
rect 3007 8382 3041 8416
rect 3295 8382 3329 8416
rect 4543 8382 4577 8416
rect 7903 8382 7937 8416
rect 10511 8382 10545 8416
rect 11071 8382 11105 8416
rect 11359 8382 11393 8416
rect 12127 8382 12161 8416
rect 13663 8382 13697 8416
rect 16255 8382 16289 8416
rect 25663 8382 25697 8416
rect 32575 8382 32609 8416
rect 48895 8382 48929 8416
rect 52447 8382 52481 8416
rect 52735 8382 52769 8416
rect 53215 8382 53249 8416
rect 9439 8308 9473 8342
rect 9823 8308 9857 8342
rect 17023 8308 17057 8342
rect 49759 8308 49793 8342
rect 54079 8308 54113 8342
rect 55231 8308 55265 8342
rect 55999 8308 56033 8342
rect 57151 8308 57185 8342
rect 1663 8234 1697 8268
rect 2527 8234 2561 8268
rect 3199 8234 3233 8268
rect 4447 8234 4481 8268
rect 7807 8234 7841 8268
rect 9727 8234 9761 8268
rect 10591 8234 10625 8268
rect 11263 8234 11297 8268
rect 12031 8234 12065 8268
rect 12511 8234 12545 8268
rect 12799 8234 12833 8268
rect 13567 8234 13601 8268
rect 16159 8234 16193 8268
rect 16927 8234 16961 8268
rect 48127 8234 48161 8268
rect 48223 8234 48257 8268
rect 48991 8234 49025 8268
rect 49663 8234 49697 8268
rect 52543 8234 52577 8268
rect 53311 8234 53345 8268
rect 53983 8234 54017 8268
rect 5311 8160 5345 8194
rect 10303 8086 10337 8120
rect 45535 8086 45569 8120
rect 50527 8086 50561 8120
rect 2143 7864 2177 7898
rect 3679 7864 3713 7898
rect 7615 7864 7649 7898
rect 9055 7864 9089 7898
rect 29023 7864 29057 7898
rect 36511 7864 36545 7898
rect 41503 7864 41537 7898
rect 42271 7864 42305 7898
rect 45247 7864 45281 7898
rect 47551 7864 47585 7898
rect 48127 7864 48161 7898
rect 50719 7864 50753 7898
rect 10687 7790 10721 7824
rect 25087 7790 25121 7824
rect 27967 7790 28001 7824
rect 2527 7716 2561 7750
rect 4063 7716 4097 7750
rect 4831 7716 4865 7750
rect 9439 7716 9473 7750
rect 10111 7716 10145 7750
rect 10975 7716 11009 7750
rect 13855 7716 13889 7750
rect 13951 7716 13985 7750
rect 15583 7716 15617 7750
rect 15871 7716 15905 7750
rect 20959 7716 20993 7750
rect 23647 7716 23681 7750
rect 23935 7716 23969 7750
rect 24703 7716 24737 7750
rect 25471 7716 25505 7750
rect 25951 7716 25985 7750
rect 26143 7716 26177 7750
rect 27007 7716 27041 7750
rect 28255 7716 28289 7750
rect 29311 7716 29345 7750
rect 29887 7716 29921 7750
rect 30175 7716 30209 7750
rect 33535 7716 33569 7750
rect 33727 7716 33761 7750
rect 34303 7716 34337 7750
rect 34591 7716 34625 7750
rect 35359 7716 35393 7750
rect 36127 7716 36161 7750
rect 36799 7716 36833 7750
rect 38527 7716 38561 7750
rect 38719 7716 38753 7750
rect 39295 7716 39329 7750
rect 39487 7716 39521 7750
rect 39583 7716 39617 7750
rect 40351 7716 40385 7750
rect 41023 7716 41057 7750
rect 41887 7716 41921 7750
rect 42655 7716 42689 7750
rect 44863 7716 44897 7750
rect 45535 7716 45569 7750
rect 46399 7716 46433 7750
rect 47839 7716 47873 7750
rect 49375 7716 49409 7750
rect 50143 7716 50177 7750
rect 51007 7716 51041 7750
rect 51103 7716 51137 7750
rect 53407 7716 53441 7750
rect 1567 7642 1601 7676
rect 3295 7642 3329 7676
rect 10207 7642 10241 7676
rect 13183 7642 13217 7676
rect 28927 7642 28961 7676
rect 31231 7642 31265 7676
rect 46783 7642 46817 7676
rect 47071 7642 47105 7676
rect 51487 7642 51521 7676
rect 51775 7642 51809 7676
rect 55135 7642 55169 7676
rect 55807 7642 55841 7676
rect 56575 7642 56609 7676
rect 57343 7642 57377 7676
rect 5311 7568 5345 7602
rect 5599 7568 5633 7602
rect 12127 7568 12161 7602
rect 12415 7568 12449 7602
rect 31999 7568 32033 7602
rect 41119 7568 41153 7602
rect 41791 7568 41825 7602
rect 43807 7568 43841 7602
rect 44095 7568 44129 7602
rect 52639 7568 52673 7602
rect 28927 7494 28961 7528
rect 2431 7420 2465 7454
rect 3199 7420 3233 7454
rect 3967 7420 4001 7454
rect 4735 7420 4769 7454
rect 5503 7420 5537 7454
rect 9343 7420 9377 7454
rect 10879 7420 10913 7454
rect 12319 7420 12353 7454
rect 13087 7420 13121 7454
rect 15775 7420 15809 7454
rect 20863 7420 20897 7454
rect 23839 7420 23873 7454
rect 24607 7420 24641 7454
rect 25375 7420 25409 7454
rect 26239 7420 26273 7454
rect 26911 7420 26945 7454
rect 28351 7420 28385 7454
rect 29407 7420 29441 7454
rect 30079 7420 30113 7454
rect 31135 7420 31169 7454
rect 33823 7420 33857 7454
rect 34495 7420 34529 7454
rect 35263 7420 35297 7454
rect 36031 7420 36065 7454
rect 36895 7420 36929 7454
rect 38815 7420 38849 7454
rect 40255 7420 40289 7454
rect 42559 7420 42593 7454
rect 43999 7420 44033 7454
rect 44767 7420 44801 7454
rect 45631 7420 45665 7454
rect 46303 7420 46337 7454
rect 47167 7420 47201 7454
rect 47935 7420 47969 7454
rect 49279 7420 49313 7454
rect 50047 7420 50081 7454
rect 51871 7420 51905 7454
rect 52543 7420 52577 7454
rect 53311 7420 53345 7454
rect 17215 7198 17249 7232
rect 17983 7198 18017 7232
rect 18751 7198 18785 7232
rect 44575 7198 44609 7232
rect 10511 7124 10545 7158
rect 17023 7124 17057 7158
rect 23071 7124 23105 7158
rect 28351 7124 28385 7158
rect 29119 7124 29153 7158
rect 33727 7124 33761 7158
rect 39279 7124 39313 7158
rect 41119 7124 41153 7158
rect 42191 7124 42225 7158
rect 48799 7124 48833 7158
rect 49279 7124 49313 7158
rect 49951 7124 49985 7158
rect 50527 7124 50561 7158
rect 6079 7050 6113 7084
rect 13663 7050 13697 7084
rect 15103 7050 15137 7084
rect 15871 7050 15905 7084
rect 18079 7050 18113 7084
rect 18847 7050 18881 7084
rect 20383 7050 20417 7084
rect 20863 7050 20897 7084
rect 21151 7050 21185 7084
rect 21919 7050 21953 7084
rect 22687 7050 22721 7084
rect 23455 7050 23489 7084
rect 23935 7050 23969 7084
rect 24223 7050 24257 7084
rect 25663 7050 25697 7084
rect 26143 7050 26177 7084
rect 26335 7050 26369 7084
rect 26911 7050 26945 7084
rect 27199 7050 27233 7084
rect 27967 7050 28001 7084
rect 28639 7050 28673 7084
rect 29407 7050 29441 7084
rect 30943 7050 30977 7084
rect 31423 7050 31457 7084
rect 31711 7050 31745 7084
rect 32479 7050 32513 7084
rect 33247 7050 33281 7084
rect 33919 7050 33953 7084
rect 34783 7050 34817 7084
rect 36223 7050 36257 7084
rect 37471 7050 37505 7084
rect 37759 7050 37793 7084
rect 38527 7050 38561 7084
rect 39199 7050 39233 7084
rect 39487 7050 39521 7084
rect 41407 7050 41441 7084
rect 41695 7050 41729 7084
rect 43039 7050 43073 7084
rect 43807 7050 43841 7084
rect 45343 7050 45377 7084
rect 48319 7050 48353 7084
rect 48991 7050 49025 7084
rect 50239 7050 50273 7084
rect 52063 7050 52097 7084
rect 1663 6976 1697 7010
rect 2527 6976 2561 7010
rect 5023 6976 5057 7010
rect 5311 6976 5345 7010
rect 6847 6976 6881 7010
rect 11263 6976 11297 7010
rect 12703 6976 12737 7010
rect 16351 6976 16385 7010
rect 16639 6976 16673 7010
rect 36991 6976 37025 7010
rect 4447 6902 4481 6936
rect 4543 6902 4577 6936
rect 5215 6902 5249 6936
rect 5983 6902 6017 6936
rect 6751 6902 6785 6936
rect 7519 6902 7553 6936
rect 7615 6902 7649 6936
rect 8287 6902 8321 6936
rect 8383 6902 8417 6936
rect 9727 6902 9761 6936
rect 9823 6902 9857 6936
rect 10591 6902 10625 6936
rect 13567 6902 13601 6936
rect 15007 6902 15041 6936
rect 15775 6902 15809 6936
rect 17311 6902 17345 6936
rect 20287 6902 20321 6936
rect 21055 6902 21089 6936
rect 21823 6902 21857 6936
rect 22591 6902 22625 6936
rect 23359 6902 23393 6936
rect 24127 6902 24161 6936
rect 25567 6902 25601 6936
rect 26431 6902 26465 6936
rect 27103 6902 27137 6936
rect 27871 6902 27905 6936
rect 28735 6902 28769 6936
rect 29503 6902 29537 6936
rect 30847 6902 30881 6936
rect 31615 6902 31649 6936
rect 32383 6902 32417 6936
rect 33151 6902 33185 6936
rect 34015 6902 34049 6936
rect 34687 6902 34721 6936
rect 36127 6902 36161 6936
rect 36895 6902 36929 6936
rect 37663 6902 37697 6936
rect 38431 6902 38465 6936
rect 40063 6976 40097 7010
rect 47263 6976 47297 7010
rect 47551 6976 47585 7010
rect 54079 6976 54113 7010
rect 54751 6976 54785 7010
rect 55519 6976 55553 7010
rect 57823 6976 57857 7010
rect 39967 6902 40001 6936
rect 41503 6902 41537 6936
rect 42271 6902 42305 6936
rect 42943 6902 42977 6936
rect 43711 6902 43745 6936
rect 44479 6902 44513 6936
rect 45247 6902 45281 6936
rect 46399 6902 46433 6936
rect 46687 6902 46721 6936
rect 46783 6902 46817 6936
rect 47455 6902 47489 6936
rect 48223 6902 48257 6936
rect 49087 6902 49121 6936
rect 50335 6902 50369 6936
rect 51967 6902 52001 6936
rect 52735 6902 52769 6936
rect 52831 6902 52865 6936
rect 9535 6828 9569 6862
rect 39487 6828 39521 6862
rect 8095 6754 8129 6788
rect 8671 6754 8705 6788
rect 38911 6754 38945 6788
rect 44191 6754 44225 6788
rect 52447 6754 52481 6788
rect 5407 6532 5441 6566
rect 18847 6532 18881 6566
rect 20479 6532 20513 6566
rect 22591 6532 22625 6566
rect 24127 6532 24161 6566
rect 27871 6532 27905 6566
rect 31807 6532 31841 6566
rect 45439 6532 45473 6566
rect 46207 6532 46241 6566
rect 46495 6532 46529 6566
rect 50527 6532 50561 6566
rect 51295 6532 51329 6566
rect 7615 6458 7649 6492
rect 5695 6384 5729 6418
rect 7039 6384 7073 6418
rect 13663 6384 13697 6418
rect 13951 6384 13985 6418
rect 14719 6384 14753 6418
rect 15487 6384 15521 6418
rect 16255 6384 16289 6418
rect 17695 6384 17729 6418
rect 18463 6384 18497 6418
rect 19231 6384 19265 6418
rect 20767 6384 20801 6418
rect 21439 6384 21473 6418
rect 22975 6384 23009 6418
rect 23743 6384 23777 6418
rect 24415 6384 24449 6418
rect 28255 6384 28289 6418
rect 29023 6384 29057 6418
rect 30655 6384 30689 6418
rect 32191 6384 32225 6418
rect 34303 6384 34337 6418
rect 35071 6384 35105 6418
rect 37279 6384 37313 6418
rect 41311 6384 41345 6418
rect 42847 6384 42881 6418
rect 44095 6384 44129 6418
rect 44863 6384 44897 6418
rect 1567 6310 1601 6344
rect 2335 6310 2369 6344
rect 3199 6310 3233 6344
rect 3967 6310 4001 6344
rect 4735 6310 4769 6344
rect 9439 6310 9473 6344
rect 10207 6310 10241 6344
rect 10975 6310 11009 6344
rect 12223 6310 12257 6344
rect 13087 6310 13121 6344
rect 19999 6310 20033 6344
rect 21535 6310 21569 6344
rect 25663 6310 25697 6344
rect 26815 6310 26849 6344
rect 29695 6310 29729 6344
rect 31231 6310 31265 6344
rect 34223 6310 34257 6344
rect 36319 6310 36353 6344
rect 38911 6310 38945 6344
rect 40351 6310 40385 6344
rect 41887 6310 41921 6344
rect 6847 6236 6881 6270
rect 7135 6236 7169 6270
rect 33535 6236 33569 6270
rect 50911 6384 50945 6418
rect 51583 6384 51617 6418
rect 45535 6310 45569 6344
rect 46975 6310 47009 6344
rect 47743 6310 47777 6344
rect 49183 6310 49217 6344
rect 49951 6310 49985 6344
rect 50815 6310 50849 6344
rect 52063 6310 52097 6344
rect 52351 6310 52385 6344
rect 53311 6310 53345 6344
rect 54463 6310 54497 6344
rect 55231 6310 55265 6344
rect 55999 6310 56033 6344
rect 57055 6310 57089 6344
rect 57823 6310 57857 6344
rect 45439 6162 45473 6196
rect 5599 6088 5633 6122
rect 13855 6088 13889 6122
rect 14623 6088 14657 6122
rect 15391 6088 15425 6122
rect 16159 6088 16193 6122
rect 17599 6088 17633 6122
rect 18367 6088 18401 6122
rect 19135 6088 19169 6122
rect 19903 6088 19937 6122
rect 20671 6088 20705 6122
rect 22879 6088 22913 6122
rect 23647 6088 23681 6122
rect 24511 6088 24545 6122
rect 28159 6088 28193 6122
rect 28927 6088 28961 6122
rect 30559 6088 30593 6122
rect 32095 6088 32129 6122
rect 33439 6088 33473 6122
rect 34975 6088 35009 6122
rect 37183 6088 37217 6122
rect 41215 6088 41249 6122
rect 42751 6088 42785 6122
rect 43999 6088 44033 6122
rect 44767 6088 44801 6122
rect 51679 6088 51713 6122
rect 52447 6088 52481 6122
rect 12127 5718 12161 5752
rect 1567 5644 1601 5678
rect 2911 5644 2945 5678
rect 4447 5644 4481 5678
rect 5215 5644 5249 5678
rect 6847 5644 6881 5678
rect 7615 5644 7649 5678
rect 7999 5644 8033 5678
rect 8383 5644 8417 5678
rect 9631 5644 9665 5678
rect 10399 5644 10433 5678
rect 11167 5644 11201 5678
rect 12607 5644 12641 5678
rect 13471 5644 13505 5678
rect 15007 5644 15041 5678
rect 15871 5644 15905 5678
rect 16543 5644 16577 5678
rect 17311 5644 17345 5678
rect 18751 5644 18785 5678
rect 20191 5644 20225 5678
rect 20959 5644 20993 5678
rect 21727 5644 21761 5678
rect 22495 5644 22529 5678
rect 23263 5644 23297 5678
rect 24031 5644 24065 5678
rect 25471 5644 25505 5678
rect 26239 5644 26273 5678
rect 27007 5644 27041 5678
rect 27775 5644 27809 5678
rect 28543 5644 28577 5678
rect 29311 5644 29345 5678
rect 30751 5644 30785 5678
rect 31519 5644 31553 5678
rect 32287 5644 32321 5678
rect 33151 5644 33185 5678
rect 33823 5644 33857 5678
rect 34687 5644 34721 5678
rect 36127 5644 36161 5678
rect 36799 5644 36833 5678
rect 37567 5644 37601 5678
rect 38335 5644 38369 5678
rect 39103 5644 39137 5678
rect 39871 5644 39905 5678
rect 41311 5644 41345 5678
rect 42079 5644 42113 5678
rect 42847 5644 42881 5678
rect 43615 5644 43649 5678
rect 44383 5644 44417 5678
rect 45151 5644 45185 5678
rect 46591 5644 46625 5678
rect 47359 5644 47393 5678
rect 48127 5644 48161 5678
rect 48991 5644 49025 5678
rect 49663 5644 49697 5678
rect 50527 5644 50561 5678
rect 52159 5644 52193 5678
rect 52927 5644 52961 5678
rect 53695 5644 53729 5678
rect 54463 5644 54497 5678
rect 55999 5644 56033 5678
rect 57439 5644 57473 5678
rect 5983 5570 6017 5604
rect 6079 5570 6113 5604
rect 7999 5496 8033 5530
rect 17983 5422 18017 5456
rect 18271 5422 18305 5456
rect 55423 5422 55457 5456
rect 7519 5126 7553 5160
rect 1567 4978 1601 5012
rect 2335 4978 2369 5012
rect 3103 4978 3137 5012
rect 4159 4978 4193 5012
rect 5407 4978 5441 5012
rect 6943 4978 6977 5012
rect 9247 4978 9281 5012
rect 10111 4978 10145 5012
rect 10879 4978 10913 5012
rect 12223 4978 12257 5012
rect 12991 4978 13025 5012
rect 13951 4978 13985 5012
rect 14719 4978 14753 5012
rect 15487 4978 15521 5012
rect 16351 4978 16385 5012
rect 17503 4978 17537 5012
rect 18271 4978 18305 5012
rect 19039 4978 19073 5012
rect 19807 4978 19841 5012
rect 20671 4978 20705 5012
rect 21343 4978 21377 5012
rect 22783 4978 22817 5012
rect 23551 4978 23585 5012
rect 24319 4978 24353 5012
rect 25087 4978 25121 5012
rect 25855 4978 25889 5012
rect 26623 4978 26657 5012
rect 28063 4978 28097 5012
rect 28927 4978 28961 5012
rect 29599 4978 29633 5012
rect 30367 4978 30401 5012
rect 31135 4978 31169 5012
rect 31903 4978 31937 5012
rect 33343 4978 33377 5012
rect 34111 4978 34145 5012
rect 34879 4978 34913 5012
rect 35647 4978 35681 5012
rect 36415 4978 36449 5012
rect 37183 4978 37217 5012
rect 38623 4978 38657 5012
rect 39391 4978 39425 5012
rect 40159 4978 40193 5012
rect 40927 4978 40961 5012
rect 41695 4978 41729 5012
rect 42463 4978 42497 5012
rect 43903 4978 43937 5012
rect 44767 4978 44801 5012
rect 45439 4978 45473 5012
rect 46207 4978 46241 5012
rect 46975 4978 47009 5012
rect 47743 4978 47777 5012
rect 49375 4978 49409 5012
rect 50431 4978 50465 5012
rect 51103 4978 51137 5012
rect 51871 4978 51905 5012
rect 52639 4978 52673 5012
rect 54463 4978 54497 5012
rect 55615 4978 55649 5012
rect 56383 4978 56417 5012
rect 57055 4978 57089 5012
rect 15775 4534 15809 4568
rect 20575 4534 20609 4568
rect 38143 4534 38177 4568
rect 54847 4534 54881 4568
rect 55135 4534 55169 4568
rect 16543 4460 16577 4494
rect 17311 4460 17345 4494
rect 38335 4386 38369 4420
rect 1567 4312 1601 4346
rect 2335 4312 2369 4346
rect 3103 4312 3137 4346
rect 4351 4312 4385 4346
rect 5119 4312 5153 4346
rect 5887 4312 5921 4346
rect 6655 4312 6689 4346
rect 7423 4312 7457 4346
rect 8191 4312 8225 4346
rect 9631 4312 9665 4346
rect 10399 4312 10433 4346
rect 11167 4312 11201 4346
rect 11935 4312 11969 4346
rect 12703 4312 12737 4346
rect 13567 4312 13601 4346
rect 15487 4312 15521 4346
rect 16255 4312 16289 4346
rect 17023 4312 17057 4346
rect 17791 4312 17825 4346
rect 18559 4312 18593 4346
rect 20287 4312 20321 4346
rect 21055 4312 21089 4346
rect 21823 4312 21857 4346
rect 23263 4312 23297 4346
rect 24031 4312 24065 4346
rect 25471 4312 25505 4346
rect 26239 4312 26273 4346
rect 27007 4312 27041 4346
rect 28351 4312 28385 4346
rect 29119 4312 29153 4346
rect 30943 4312 30977 4346
rect 31711 4312 31745 4346
rect 32767 4312 32801 4346
rect 33919 4312 33953 4346
rect 34687 4312 34721 4346
rect 36031 4312 36065 4346
rect 36799 4312 36833 4346
rect 37567 4312 37601 4346
rect 39007 4312 39041 4346
rect 39775 4312 39809 4346
rect 41983 4312 42017 4346
rect 42751 4312 42785 4346
rect 43519 4312 43553 4346
rect 44959 4312 44993 4346
rect 46783 4312 46817 4346
rect 47551 4312 47585 4346
rect 48319 4312 48353 4346
rect 49087 4312 49121 4346
rect 49855 4312 49889 4346
rect 50623 4312 50657 4346
rect 51871 4312 51905 4346
rect 52639 4312 52673 4346
rect 53407 4312 53441 4346
rect 54175 4312 54209 4346
rect 55615 4312 55649 4346
rect 57151 4312 57185 4346
rect 13951 3868 13985 3902
rect 15487 3868 15521 3902
rect 17791 3868 17825 3902
rect 18559 3868 18593 3902
rect 20095 3720 20129 3754
rect 1567 3646 1601 3680
rect 2335 3646 2369 3680
rect 3103 3646 3137 3680
rect 3871 3646 3905 3680
rect 4639 3646 4673 3680
rect 5599 3646 5633 3680
rect 6943 3646 6977 3680
rect 7711 3646 7745 3680
rect 8479 3646 8513 3680
rect 9247 3646 9281 3680
rect 10015 3646 10049 3680
rect 10783 3646 10817 3680
rect 12991 3646 13025 3680
rect 13663 3646 13697 3680
rect 14431 3646 14465 3680
rect 15199 3646 15233 3680
rect 15967 3646 16001 3680
rect 17503 3646 17537 3680
rect 18271 3646 18305 3680
rect 19039 3646 19073 3680
rect 19807 3646 19841 3680
rect 21343 3646 21377 3680
rect 22783 3646 22817 3680
rect 23551 3646 23585 3680
rect 24319 3646 24353 3680
rect 25087 3646 25121 3680
rect 25855 3646 25889 3680
rect 26623 3646 26657 3680
rect 28063 3646 28097 3680
rect 28831 3646 28865 3680
rect 29599 3646 29633 3680
rect 30367 3646 30401 3680
rect 31135 3646 31169 3680
rect 31903 3646 31937 3680
rect 33343 3646 33377 3680
rect 34111 3646 34145 3680
rect 34879 3646 34913 3680
rect 35647 3646 35681 3680
rect 36415 3646 36449 3680
rect 37183 3646 37217 3680
rect 38623 3646 38657 3680
rect 39391 3646 39425 3680
rect 40159 3646 40193 3680
rect 40927 3646 40961 3680
rect 41695 3646 41729 3680
rect 42463 3646 42497 3680
rect 43903 3646 43937 3680
rect 44671 3646 44705 3680
rect 45439 3646 45473 3680
rect 46207 3646 46241 3680
rect 46975 3646 47009 3680
rect 47743 3646 47777 3680
rect 49183 3646 49217 3680
rect 50527 3646 50561 3680
rect 51199 3646 51233 3680
rect 51967 3646 52001 3680
rect 52735 3646 52769 3680
rect 54463 3646 54497 3680
rect 55231 3646 55265 3680
rect 55999 3646 56033 3680
rect 56767 3646 56801 3680
rect 57535 3646 57569 3680
rect 20767 3572 20801 3606
rect 20671 3424 20705 3458
rect 13279 3202 13313 3236
rect 14047 3202 14081 3236
rect 15391 3202 15425 3236
rect 18079 3202 18113 3236
rect 20767 3202 20801 3236
rect 43327 3202 43361 3236
rect 18847 3128 18881 3162
rect 51775 3054 51809 3088
rect 1567 2980 1601 3014
rect 2335 2980 2369 3014
rect 3103 2980 3137 3014
rect 4927 2980 4961 3014
rect 5695 2980 5729 3014
rect 7039 2980 7073 3014
rect 7807 2980 7841 3014
rect 9727 2980 9761 3014
rect 10495 2980 10529 3014
rect 12991 2980 13025 3014
rect 13759 2980 13793 3014
rect 15103 2980 15137 3014
rect 16639 2980 16673 3014
rect 17791 2980 17825 3014
rect 18559 2980 18593 3014
rect 20479 2980 20513 3014
rect 21247 2980 21281 3014
rect 23167 2980 23201 3014
rect 23935 2980 23969 3014
rect 25855 2980 25889 3014
rect 26623 2980 26657 3014
rect 28543 2980 28577 3014
rect 29311 2980 29345 3014
rect 31231 2980 31265 3014
rect 31999 2980 32033 3014
rect 33919 2980 33953 3014
rect 34687 2980 34721 3014
rect 36607 2980 36641 3014
rect 37375 2980 37409 3014
rect 39295 2980 39329 3014
rect 40063 2980 40097 3014
rect 41983 2980 42017 3014
rect 42751 2980 42785 3014
rect 44671 2980 44705 3014
rect 45439 2980 45473 3014
rect 47359 2980 47393 3014
rect 48127 2980 48161 3014
rect 50047 2980 50081 3014
rect 50815 2980 50849 3014
rect 52735 2980 52769 3014
rect 53503 2980 53537 3014
rect 55423 2980 55457 3014
rect 56191 2980 56225 3014
rect 19231 2906 19265 2940
rect 19519 2906 19553 2940
rect 40735 2906 40769 2940
rect 41023 2906 41057 2940
rect 43519 2906 43553 2940
rect 8767 2832 8801 2866
rect 16063 2758 16097 2792
rect 32959 2758 32993 2792
rect 54463 2758 54497 2792
<< metal1 >>
rect 1152 57302 58848 57324
rect 1152 57250 4294 57302
rect 4346 57250 4358 57302
rect 4410 57250 4422 57302
rect 4474 57250 4486 57302
rect 4538 57250 35014 57302
rect 35066 57250 35078 57302
rect 35130 57250 35142 57302
rect 35194 57250 35206 57302
rect 35258 57250 58848 57302
rect 1152 57228 58848 57250
rect 1744 56991 1750 57043
rect 1802 57031 1808 57043
rect 1802 57003 2846 57031
rect 1802 56991 1808 57003
rect 208 56917 214 56969
rect 266 56957 272 56969
rect 2818 56966 2846 57003
rect 3280 56991 3286 57043
rect 3338 57031 3344 57043
rect 3338 57003 5822 57031
rect 3338 56991 3344 57003
rect 1939 56960 1997 56966
rect 1939 56957 1951 56960
rect 266 56929 1951 56957
rect 266 56917 272 56929
rect 1939 56926 1951 56929
rect 1985 56926 1997 56960
rect 1939 56920 1997 56926
rect 2803 56960 2861 56966
rect 2803 56926 2815 56960
rect 2849 56926 2861 56960
rect 2803 56920 2861 56926
rect 4912 56917 4918 56969
rect 4970 56957 4976 56969
rect 5794 56966 5822 57003
rect 9616 56991 9622 57043
rect 9674 57031 9680 57043
rect 9907 57034 9965 57040
rect 9907 57031 9919 57034
rect 9674 57003 9919 57031
rect 9674 56991 9680 57003
rect 9907 57000 9919 57003
rect 9953 57000 9965 57034
rect 9907 56994 9965 57000
rect 11248 56991 11254 57043
rect 11306 57031 11312 57043
rect 13939 57034 13997 57040
rect 11306 57003 11486 57031
rect 11306 56991 11312 57003
rect 5299 56960 5357 56966
rect 5299 56957 5311 56960
rect 4970 56929 5311 56957
rect 4970 56917 4976 56929
rect 5299 56926 5311 56929
rect 5345 56926 5357 56960
rect 5299 56920 5357 56926
rect 5779 56960 5837 56966
rect 5779 56926 5791 56960
rect 5825 56926 5837 56960
rect 5779 56920 5837 56926
rect 6448 56917 6454 56969
rect 6506 56957 6512 56969
rect 7411 56960 7469 56966
rect 7411 56957 7423 56960
rect 6506 56929 7423 56957
rect 6506 56917 6512 56929
rect 7411 56926 7423 56929
rect 7457 56926 7469 56960
rect 8080 56957 8086 56969
rect 8041 56929 8086 56957
rect 7411 56920 7469 56926
rect 8080 56917 8086 56929
rect 8138 56917 8144 56969
rect 11458 56966 11486 57003
rect 13939 57000 13951 57034
rect 13985 57031 13997 57034
rect 16432 57031 16438 57043
rect 13985 57003 16438 57031
rect 13985 57000 13997 57003
rect 13939 56994 13997 57000
rect 16432 56991 16438 57003
rect 16490 56991 16496 57043
rect 29104 56991 29110 57043
rect 29162 57031 29168 57043
rect 32659 57034 32717 57040
rect 32659 57031 32671 57034
rect 29162 57003 32671 57031
rect 29162 56991 29168 57003
rect 32659 57000 32671 57003
rect 32705 57000 32717 57034
rect 32659 56994 32717 57000
rect 11443 56960 11501 56966
rect 11443 56926 11455 56960
rect 11489 56926 11501 56960
rect 11443 56920 11501 56926
rect 12784 56917 12790 56969
rect 12842 56957 12848 56969
rect 13171 56960 13229 56966
rect 13171 56957 13183 56960
rect 12842 56929 13183 56957
rect 12842 56917 12848 56929
rect 13171 56926 13183 56929
rect 13217 56926 13229 56960
rect 13171 56920 13229 56926
rect 14416 56917 14422 56969
rect 14474 56957 14480 56969
rect 15091 56960 15149 56966
rect 15091 56957 15103 56960
rect 14474 56929 15103 56957
rect 14474 56917 14480 56929
rect 15091 56926 15103 56929
rect 15137 56926 15149 56960
rect 15091 56920 15149 56926
rect 15952 56917 15958 56969
rect 16010 56957 16016 56969
rect 16339 56960 16397 56966
rect 16339 56957 16351 56960
rect 16010 56929 16351 56957
rect 16010 56917 16016 56929
rect 16339 56926 16351 56929
rect 16385 56926 16397 56960
rect 16339 56920 16397 56926
rect 17488 56917 17494 56969
rect 17546 56957 17552 56969
rect 18163 56960 18221 56966
rect 18163 56957 18175 56960
rect 17546 56929 18175 56957
rect 17546 56917 17552 56929
rect 18163 56926 18175 56929
rect 18209 56926 18221 56960
rect 18163 56920 18221 56926
rect 19120 56917 19126 56969
rect 19178 56957 19184 56969
rect 19507 56960 19565 56966
rect 19507 56957 19519 56960
rect 19178 56929 19519 56957
rect 19178 56917 19184 56929
rect 19507 56926 19519 56929
rect 19553 56926 19565 56960
rect 19507 56920 19565 56926
rect 20656 56917 20662 56969
rect 20714 56957 20720 56969
rect 21043 56960 21101 56966
rect 21043 56957 21055 56960
rect 20714 56929 21055 56957
rect 20714 56917 20720 56929
rect 21043 56926 21055 56929
rect 21089 56926 21101 56960
rect 21043 56920 21101 56926
rect 22003 56960 22061 56966
rect 22003 56926 22015 56960
rect 22049 56957 22061 56960
rect 22288 56957 22294 56969
rect 22049 56929 22294 56957
rect 22049 56926 22061 56929
rect 22003 56920 22061 56926
rect 22288 56917 22294 56929
rect 22346 56917 22352 56969
rect 23824 56917 23830 56969
rect 23882 56957 23888 56969
rect 24211 56960 24269 56966
rect 24211 56957 24223 56960
rect 23882 56929 24223 56957
rect 23882 56917 23888 56929
rect 24211 56926 24223 56929
rect 24257 56926 24269 56960
rect 24211 56920 24269 56926
rect 25456 56917 25462 56969
rect 25514 56957 25520 56969
rect 25939 56960 25997 56966
rect 25939 56957 25951 56960
rect 25514 56929 25951 56957
rect 25514 56917 25520 56929
rect 25939 56926 25951 56929
rect 25985 56926 25997 56960
rect 25939 56920 25997 56926
rect 26992 56917 26998 56969
rect 27050 56957 27056 56969
rect 27379 56960 27437 56966
rect 27379 56957 27391 56960
rect 27050 56929 27391 56957
rect 27050 56917 27056 56929
rect 27379 56926 27391 56929
rect 27425 56926 27437 56960
rect 27379 56920 27437 56926
rect 28624 56917 28630 56969
rect 28682 56957 28688 56969
rect 29011 56960 29069 56966
rect 29011 56957 29023 56960
rect 28682 56929 29023 56957
rect 28682 56917 28688 56929
rect 29011 56926 29023 56929
rect 29057 56926 29069 56960
rect 29011 56920 29069 56926
rect 30067 56960 30125 56966
rect 30067 56926 30079 56960
rect 30113 56957 30125 56960
rect 30160 56957 30166 56969
rect 30113 56929 30166 56957
rect 30113 56926 30125 56929
rect 30067 56920 30125 56926
rect 30160 56917 30166 56929
rect 30218 56917 30224 56969
rect 31696 56957 31702 56969
rect 31657 56929 31702 56957
rect 31696 56917 31702 56929
rect 31754 56917 31760 56969
rect 33328 56917 33334 56969
rect 33386 56957 33392 56969
rect 34291 56960 34349 56966
rect 34291 56957 34303 56960
rect 33386 56929 34303 56957
rect 33386 56917 33392 56929
rect 34291 56926 34303 56929
rect 34337 56926 34349 56960
rect 34864 56957 34870 56969
rect 34825 56929 34870 56957
rect 34291 56920 34349 56926
rect 34864 56917 34870 56929
rect 34922 56917 34928 56969
rect 38032 56957 38038 56969
rect 37993 56929 38038 56957
rect 38032 56917 38038 56929
rect 38090 56917 38096 56969
rect 41200 56917 41206 56969
rect 41258 56957 41264 56969
rect 41971 56960 42029 56966
rect 41971 56957 41983 56960
rect 41258 56929 41983 56957
rect 41258 56917 41264 56929
rect 41971 56926 41983 56929
rect 42017 56926 42029 56960
rect 41971 56920 42029 56926
rect 44368 56917 44374 56969
rect 44426 56957 44432 56969
rect 44659 56960 44717 56966
rect 44659 56957 44671 56960
rect 44426 56929 44671 56957
rect 44426 56917 44432 56929
rect 44659 56926 44671 56929
rect 44705 56926 44717 56960
rect 44659 56920 44717 56926
rect 47536 56917 47542 56969
rect 47594 56957 47600 56969
rect 47594 56929 47639 56957
rect 47594 56917 47600 56929
rect 49936 56917 49942 56969
rect 49994 56957 50000 56969
rect 52144 56957 52150 56969
rect 49994 56929 52150 56957
rect 49994 56917 50000 56929
rect 52144 56917 52150 56929
rect 52202 56917 52208 56969
rect 53872 56957 53878 56969
rect 53833 56929 53878 56957
rect 53872 56917 53878 56929
rect 53930 56917 53936 56969
rect 1747 56886 1805 56892
rect 1747 56852 1759 56886
rect 1793 56883 1805 56886
rect 2032 56883 2038 56895
rect 1793 56855 2038 56883
rect 1793 56852 1805 56855
rect 1747 56846 1805 56852
rect 2032 56843 2038 56855
rect 2090 56843 2096 56895
rect 2611 56886 2669 56892
rect 2611 56852 2623 56886
rect 2657 56883 2669 56886
rect 3568 56883 3574 56895
rect 2657 56855 3574 56883
rect 2657 56852 2669 56855
rect 2611 56846 2669 56852
rect 3568 56843 3574 56855
rect 3626 56843 3632 56895
rect 5104 56883 5110 56895
rect 5065 56855 5110 56883
rect 5104 56843 5110 56855
rect 5162 56843 5168 56895
rect 7216 56843 7222 56895
rect 7274 56883 7280 56895
rect 11248 56883 11254 56895
rect 7274 56855 7319 56883
rect 11209 56855 11254 56883
rect 7274 56843 7280 56855
rect 11248 56843 11254 56855
rect 11306 56843 11312 56895
rect 12976 56883 12982 56895
rect 12937 56855 12982 56883
rect 12976 56843 12982 56855
rect 13034 56843 13040 56895
rect 14035 56886 14093 56892
rect 14035 56852 14047 56886
rect 14081 56852 14093 56886
rect 16144 56883 16150 56895
rect 16105 56855 16150 56883
rect 14035 56846 14093 56852
rect 14050 56809 14078 56846
rect 16144 56843 16150 56855
rect 16202 56843 16208 56895
rect 17968 56883 17974 56895
rect 17929 56855 17974 56883
rect 17968 56843 17974 56855
rect 18026 56843 18032 56895
rect 19312 56883 19318 56895
rect 19273 56855 19318 56883
rect 19312 56843 19318 56855
rect 19370 56843 19376 56895
rect 20848 56883 20854 56895
rect 20809 56855 20854 56883
rect 20848 56843 20854 56855
rect 20906 56843 20912 56895
rect 24016 56883 24022 56895
rect 23977 56855 24022 56883
rect 24016 56843 24022 56855
rect 24074 56843 24080 56895
rect 27184 56883 27190 56895
rect 27145 56855 27190 56883
rect 27184 56843 27190 56855
rect 27242 56843 27248 56895
rect 28816 56883 28822 56895
rect 28777 56855 28822 56883
rect 28816 56843 28822 56855
rect 28874 56843 28880 56895
rect 32371 56886 32429 56892
rect 32371 56852 32383 56886
rect 32417 56883 32429 56886
rect 32560 56883 32566 56895
rect 32417 56855 32566 56883
rect 32417 56852 32429 56855
rect 32371 56846 32429 56852
rect 32560 56843 32566 56855
rect 32618 56843 32624 56895
rect 34096 56883 34102 56895
rect 34057 56855 34102 56883
rect 34096 56843 34102 56855
rect 34154 56843 34160 56895
rect 36496 56843 36502 56895
rect 36554 56883 36560 56895
rect 36979 56886 37037 56892
rect 36979 56883 36991 56886
rect 36554 56855 36991 56883
rect 36554 56843 36560 56855
rect 36979 56852 36991 56855
rect 37025 56852 37037 56886
rect 36979 56846 37037 56852
rect 39664 56843 39670 56895
rect 39722 56883 39728 56895
rect 40051 56886 40109 56892
rect 40051 56883 40063 56886
rect 39722 56855 40063 56883
rect 39722 56843 39728 56855
rect 40051 56852 40063 56855
rect 40097 56852 40109 56886
rect 40723 56886 40781 56892
rect 40723 56883 40735 56886
rect 40051 56846 40109 56852
rect 40450 56855 40735 56883
rect 26704 56809 26710 56821
rect 14050 56781 26710 56809
rect 26704 56769 26710 56781
rect 26762 56769 26768 56821
rect 40450 56747 40478 56855
rect 40723 56852 40735 56855
rect 40769 56852 40781 56886
rect 40723 56846 40781 56852
rect 42832 56843 42838 56895
rect 42890 56883 42896 56895
rect 43219 56886 43277 56892
rect 43219 56883 43231 56886
rect 42890 56855 43231 56883
rect 42890 56843 42896 56855
rect 43219 56852 43231 56855
rect 43265 56852 43277 56886
rect 43219 56846 43277 56852
rect 45904 56843 45910 56895
rect 45962 56883 45968 56895
rect 46291 56886 46349 56892
rect 46291 56883 46303 56886
rect 45962 56855 46303 56883
rect 45962 56843 45968 56855
rect 46291 56852 46303 56855
rect 46337 56852 46349 56886
rect 46291 56846 46349 56852
rect 48979 56886 49037 56892
rect 48979 56852 48991 56886
rect 49025 56883 49037 56886
rect 49072 56883 49078 56895
rect 49025 56855 49078 56883
rect 49025 56852 49037 56855
rect 48979 56846 49037 56852
rect 49072 56843 49078 56855
rect 49130 56843 49136 56895
rect 50704 56843 50710 56895
rect 50762 56883 50768 56895
rect 51091 56886 51149 56892
rect 51091 56883 51103 56886
rect 50762 56855 51103 56883
rect 50762 56843 50768 56855
rect 51091 56852 51103 56855
rect 51137 56852 51149 56886
rect 51091 56846 51149 56852
rect 52240 56843 52246 56895
rect 52298 56883 52304 56895
rect 53107 56886 53165 56892
rect 53107 56883 53119 56886
rect 52298 56855 53119 56883
rect 52298 56843 52304 56855
rect 53107 56852 53119 56855
rect 53153 56852 53165 56886
rect 53107 56846 53165 56852
rect 55408 56843 55414 56895
rect 55466 56883 55472 56895
rect 55795 56886 55853 56892
rect 55795 56883 55807 56886
rect 55466 56855 55807 56883
rect 55466 56843 55472 56855
rect 55795 56852 55807 56855
rect 55841 56852 55853 56886
rect 57040 56883 57046 56895
rect 57001 56855 57046 56883
rect 55795 56846 55853 56852
rect 57040 56843 57046 56855
rect 57098 56843 57104 56895
rect 47920 56769 47926 56821
rect 47978 56809 47984 56821
rect 54832 56809 54838 56821
rect 47978 56781 54838 56809
rect 47978 56769 47984 56781
rect 54832 56769 54838 56781
rect 54890 56769 54896 56821
rect 9808 56735 9814 56747
rect 9769 56707 9814 56735
rect 9808 56695 9814 56707
rect 9866 56695 9872 56747
rect 36688 56735 36694 56747
rect 36649 56707 36694 56735
rect 36688 56695 36694 56707
rect 36746 56695 36752 56747
rect 39760 56735 39766 56747
rect 39721 56707 39766 56735
rect 39760 56695 39766 56707
rect 39818 56695 39824 56747
rect 40432 56735 40438 56747
rect 40393 56707 40438 56735
rect 40432 56695 40438 56707
rect 40490 56695 40496 56747
rect 40816 56735 40822 56747
rect 40777 56707 40822 56735
rect 40816 56695 40822 56707
rect 40874 56695 40880 56747
rect 42928 56735 42934 56747
rect 42889 56707 42934 56735
rect 42928 56695 42934 56707
rect 42986 56695 42992 56747
rect 46003 56738 46061 56744
rect 46003 56704 46015 56738
rect 46049 56735 46061 56738
rect 46096 56735 46102 56747
rect 46049 56707 46102 56735
rect 46049 56704 46061 56707
rect 46003 56698 46061 56704
rect 46096 56695 46102 56707
rect 46154 56695 46160 56747
rect 48688 56735 48694 56747
rect 48649 56707 48694 56735
rect 48688 56695 48694 56707
rect 48746 56695 48752 56747
rect 50800 56735 50806 56747
rect 50761 56707 50806 56735
rect 50800 56695 50806 56707
rect 50858 56695 50864 56747
rect 52816 56735 52822 56747
rect 52777 56707 52822 56735
rect 52816 56695 52822 56707
rect 52874 56695 52880 56747
rect 55408 56695 55414 56747
rect 55466 56735 55472 56747
rect 55507 56738 55565 56744
rect 55507 56735 55519 56738
rect 55466 56707 55519 56735
rect 55466 56695 55472 56707
rect 55507 56704 55519 56707
rect 55553 56704 55565 56738
rect 56752 56735 56758 56747
rect 56713 56707 56758 56735
rect 55507 56698 55565 56704
rect 56752 56695 56758 56707
rect 56810 56695 56816 56747
rect 1152 56636 58848 56658
rect 1152 56584 19654 56636
rect 19706 56584 19718 56636
rect 19770 56584 19782 56636
rect 19834 56584 19846 56636
rect 19898 56584 50374 56636
rect 50426 56584 50438 56636
rect 50490 56584 50502 56636
rect 50554 56584 50566 56636
rect 50618 56584 58848 56636
rect 1152 56562 58848 56584
rect 688 56473 694 56525
rect 746 56513 752 56525
rect 1651 56516 1709 56522
rect 1651 56513 1663 56516
rect 746 56485 1663 56513
rect 746 56473 752 56485
rect 1651 56482 1663 56485
rect 1697 56482 1709 56516
rect 1651 56476 1709 56482
rect 2224 56473 2230 56525
rect 2282 56513 2288 56525
rect 2419 56516 2477 56522
rect 2419 56513 2431 56516
rect 2282 56485 2431 56513
rect 2282 56473 2288 56485
rect 2419 56482 2431 56485
rect 2465 56482 2477 56516
rect 2419 56476 2477 56482
rect 2800 56473 2806 56525
rect 2858 56513 2864 56525
rect 3187 56516 3245 56522
rect 3187 56513 3199 56516
rect 2858 56485 3199 56513
rect 2858 56473 2864 56485
rect 3187 56482 3199 56485
rect 3233 56482 3245 56516
rect 3187 56476 3245 56482
rect 3856 56473 3862 56525
rect 3914 56513 3920 56525
rect 4435 56516 4493 56522
rect 4435 56513 4447 56516
rect 3914 56485 4447 56513
rect 3914 56473 3920 56485
rect 4435 56482 4447 56485
rect 4481 56482 4493 56516
rect 4435 56476 4493 56482
rect 5392 56473 5398 56525
rect 5450 56513 5456 56525
rect 5491 56516 5549 56522
rect 5491 56513 5503 56516
rect 5450 56485 5503 56513
rect 5450 56473 5456 56485
rect 5491 56482 5503 56485
rect 5537 56482 5549 56516
rect 5491 56476 5549 56482
rect 5968 56473 5974 56525
rect 6026 56513 6032 56525
rect 6259 56516 6317 56522
rect 6259 56513 6271 56516
rect 6026 56485 6271 56513
rect 6026 56473 6032 56485
rect 6259 56482 6271 56485
rect 6305 56482 6317 56516
rect 6259 56476 6317 56482
rect 7024 56473 7030 56525
rect 7082 56513 7088 56525
rect 7123 56516 7181 56522
rect 7123 56513 7135 56516
rect 7082 56485 7135 56513
rect 7082 56473 7088 56485
rect 7123 56482 7135 56485
rect 7169 56482 7181 56516
rect 7123 56476 7181 56482
rect 8467 56516 8525 56522
rect 8467 56482 8479 56516
rect 8513 56513 8525 56516
rect 8560 56513 8566 56525
rect 8513 56485 8566 56513
rect 8513 56482 8525 56485
rect 8467 56476 8525 56482
rect 8560 56473 8566 56485
rect 8618 56473 8624 56525
rect 10192 56473 10198 56525
rect 10250 56513 10256 56525
rect 10387 56516 10445 56522
rect 10387 56513 10399 56516
rect 10250 56485 10399 56513
rect 10250 56473 10256 56485
rect 10387 56482 10399 56485
rect 10433 56482 10445 56516
rect 10387 56476 10445 56482
rect 10672 56473 10678 56525
rect 10730 56513 10736 56525
rect 11059 56516 11117 56522
rect 11059 56513 11071 56516
rect 10730 56485 11071 56513
rect 10730 56473 10736 56485
rect 11059 56482 11071 56485
rect 11105 56482 11117 56516
rect 11059 56476 11117 56482
rect 11728 56473 11734 56525
rect 11786 56513 11792 56525
rect 11827 56516 11885 56522
rect 11827 56513 11839 56516
rect 11786 56485 11839 56513
rect 11786 56473 11792 56485
rect 11827 56482 11839 56485
rect 11873 56482 11885 56516
rect 11827 56476 11885 56482
rect 12304 56473 12310 56525
rect 12362 56513 12368 56525
rect 12595 56516 12653 56522
rect 12595 56513 12607 56516
rect 12362 56485 12607 56513
rect 12362 56473 12368 56485
rect 12595 56482 12607 56485
rect 12641 56482 12653 56516
rect 12595 56476 12653 56482
rect 13360 56473 13366 56525
rect 13418 56513 13424 56525
rect 13459 56516 13517 56522
rect 13459 56513 13471 56516
rect 13418 56485 13471 56513
rect 13418 56473 13424 56485
rect 13459 56482 13471 56485
rect 13505 56482 13517 56516
rect 13459 56476 13517 56482
rect 14896 56473 14902 56525
rect 14954 56513 14960 56525
rect 14995 56516 15053 56522
rect 14995 56513 15007 56516
rect 14954 56485 15007 56513
rect 14954 56473 14960 56485
rect 14995 56482 15007 56485
rect 15041 56482 15053 56516
rect 14995 56476 15053 56482
rect 17008 56473 17014 56525
rect 17066 56513 17072 56525
rect 17203 56516 17261 56522
rect 17203 56513 17215 56516
rect 17066 56485 17215 56513
rect 17066 56473 17072 56485
rect 17203 56482 17215 56485
rect 17249 56482 17261 56516
rect 17203 56476 17261 56482
rect 18064 56473 18070 56525
rect 18122 56513 18128 56525
rect 18163 56516 18221 56522
rect 18163 56513 18175 56516
rect 18122 56485 18175 56513
rect 18122 56473 18128 56485
rect 18163 56482 18175 56485
rect 18209 56482 18221 56516
rect 18163 56476 18221 56482
rect 18736 56473 18742 56525
rect 18794 56513 18800 56525
rect 19027 56516 19085 56522
rect 19027 56513 19039 56516
rect 18794 56485 19039 56513
rect 18794 56473 18800 56485
rect 19027 56482 19039 56485
rect 19073 56482 19085 56516
rect 19027 56476 19085 56482
rect 21232 56473 21238 56525
rect 21290 56513 21296 56525
rect 21331 56516 21389 56522
rect 21331 56513 21343 56516
rect 21290 56485 21343 56513
rect 21290 56473 21296 56485
rect 21331 56482 21343 56485
rect 21377 56482 21389 56516
rect 21331 56476 21389 56482
rect 21712 56473 21718 56525
rect 21770 56513 21776 56525
rect 22099 56516 22157 56522
rect 22099 56513 22111 56516
rect 21770 56485 22111 56513
rect 21770 56473 21776 56485
rect 22099 56482 22111 56485
rect 22145 56482 22157 56516
rect 22099 56476 22157 56482
rect 22768 56473 22774 56525
rect 22826 56513 22832 56525
rect 22867 56516 22925 56522
rect 22867 56513 22879 56516
rect 22826 56485 22879 56513
rect 22826 56473 22832 56485
rect 22867 56482 22879 56485
rect 22913 56482 22925 56516
rect 24400 56513 24406 56525
rect 24361 56485 24406 56513
rect 22867 56476 22925 56482
rect 24400 56473 24406 56485
rect 24458 56473 24464 56525
rect 25936 56473 25942 56525
rect 25994 56513 26000 56525
rect 26035 56516 26093 56522
rect 26035 56513 26047 56516
rect 25994 56485 26047 56513
rect 25994 56473 26000 56485
rect 26035 56482 26047 56485
rect 26081 56482 26093 56516
rect 26035 56476 26093 56482
rect 26512 56473 26518 56525
rect 26570 56513 26576 56525
rect 26899 56516 26957 56522
rect 26899 56513 26911 56516
rect 26570 56485 26911 56513
rect 26570 56473 26576 56485
rect 26899 56482 26911 56485
rect 26945 56482 26957 56516
rect 26899 56476 26957 56482
rect 27568 56473 27574 56525
rect 27626 56513 27632 56525
rect 27763 56516 27821 56522
rect 27763 56513 27775 56516
rect 27626 56485 27775 56513
rect 27626 56473 27632 56485
rect 27763 56482 27775 56485
rect 27809 56482 27821 56516
rect 27763 56476 27821 56482
rect 28048 56473 28054 56525
rect 28106 56513 28112 56525
rect 28531 56516 28589 56522
rect 28531 56513 28543 56516
rect 28106 56485 28543 56513
rect 28106 56473 28112 56485
rect 28531 56482 28543 56485
rect 28577 56482 28589 56516
rect 29680 56513 29686 56525
rect 29641 56485 29686 56513
rect 28531 56476 28589 56482
rect 29680 56473 29686 56485
rect 29738 56473 29744 56525
rect 30640 56473 30646 56525
rect 30698 56513 30704 56525
rect 30835 56516 30893 56522
rect 30835 56513 30847 56516
rect 30698 56485 30847 56513
rect 30698 56473 30704 56485
rect 30835 56482 30847 56485
rect 30881 56482 30893 56516
rect 30835 56476 30893 56482
rect 32272 56473 32278 56525
rect 32330 56513 32336 56525
rect 32371 56516 32429 56522
rect 32371 56513 32383 56516
rect 32330 56485 32383 56513
rect 32330 56473 32336 56485
rect 32371 56482 32383 56485
rect 32417 56482 32429 56516
rect 32371 56476 32429 56482
rect 33808 56473 33814 56525
rect 33866 56513 33872 56525
rect 33907 56516 33965 56522
rect 33907 56513 33919 56516
rect 33866 56485 33919 56513
rect 33866 56473 33872 56485
rect 33907 56482 33919 56485
rect 33953 56482 33965 56516
rect 33907 56476 33965 56482
rect 34384 56473 34390 56525
rect 34442 56513 34448 56525
rect 34675 56516 34733 56522
rect 34675 56513 34687 56516
rect 34442 56485 34687 56513
rect 34442 56473 34448 56485
rect 34675 56482 34687 56485
rect 34721 56482 34733 56516
rect 34675 56476 34733 56482
rect 36016 56473 36022 56525
rect 36074 56513 36080 56525
rect 36979 56516 37037 56522
rect 36979 56513 36991 56516
rect 36074 56485 36991 56513
rect 36074 56473 36080 56485
rect 36979 56482 36991 56485
rect 37025 56482 37037 56516
rect 36979 56476 37037 56482
rect 37552 56473 37558 56525
rect 37610 56513 37616 56525
rect 37651 56516 37709 56522
rect 37651 56513 37663 56516
rect 37610 56485 37663 56513
rect 37610 56473 37616 56485
rect 37651 56482 37663 56485
rect 37697 56482 37709 56516
rect 37651 56476 37709 56482
rect 38608 56473 38614 56525
rect 38666 56513 38672 56525
rect 38707 56516 38765 56522
rect 38707 56513 38719 56516
rect 38666 56485 38719 56513
rect 38666 56473 38672 56485
rect 38707 56482 38719 56485
rect 38753 56482 38765 56516
rect 40144 56513 40150 56525
rect 40105 56485 40150 56513
rect 38707 56476 38765 56482
rect 40144 56473 40150 56485
rect 40202 56473 40208 56525
rect 41776 56473 41782 56525
rect 41834 56513 41840 56525
rect 41875 56516 41933 56522
rect 41875 56513 41887 56516
rect 41834 56485 41887 56513
rect 41834 56473 41840 56485
rect 41875 56482 41887 56485
rect 41921 56482 41933 56516
rect 41875 56476 41933 56482
rect 42256 56473 42262 56525
rect 42314 56513 42320 56525
rect 42739 56516 42797 56522
rect 42739 56513 42751 56516
rect 42314 56485 42751 56513
rect 42314 56473 42320 56485
rect 42739 56482 42751 56485
rect 42785 56482 42797 56516
rect 42739 56476 42797 56482
rect 43312 56473 43318 56525
rect 43370 56513 43376 56525
rect 43507 56516 43565 56522
rect 43507 56513 43519 56516
rect 43370 56485 43519 56513
rect 43370 56473 43376 56485
rect 43507 56482 43519 56485
rect 43553 56482 43565 56516
rect 43507 56476 43565 56482
rect 43888 56473 43894 56525
rect 43946 56513 43952 56525
rect 44179 56516 44237 56522
rect 44179 56513 44191 56516
rect 43946 56485 44191 56513
rect 43946 56473 43952 56485
rect 44179 56482 44191 56485
rect 44225 56482 44237 56516
rect 44179 56476 44237 56482
rect 44944 56473 44950 56525
rect 45002 56513 45008 56525
rect 45043 56516 45101 56522
rect 45043 56513 45055 56516
rect 45002 56485 45055 56513
rect 45002 56473 45008 56485
rect 45043 56482 45055 56485
rect 45089 56482 45101 56516
rect 45043 56476 45101 56482
rect 46480 56473 46486 56525
rect 46538 56513 46544 56525
rect 46771 56516 46829 56522
rect 46771 56513 46783 56516
rect 46538 56485 46783 56513
rect 46538 56473 46544 56485
rect 46771 56482 46783 56485
rect 46817 56482 46829 56516
rect 46771 56476 46829 56482
rect 48016 56473 48022 56525
rect 48074 56513 48080 56525
rect 48115 56516 48173 56522
rect 48115 56513 48127 56516
rect 48074 56485 48127 56513
rect 48074 56473 48080 56485
rect 48115 56482 48127 56485
rect 48161 56482 48173 56516
rect 48115 56476 48173 56482
rect 49648 56473 49654 56525
rect 49706 56513 49712 56525
rect 49747 56516 49805 56522
rect 49747 56513 49759 56516
rect 49706 56485 49759 56513
rect 49706 56473 49712 56485
rect 49747 56482 49759 56485
rect 49793 56482 49805 56516
rect 49747 56476 49805 56482
rect 50128 56473 50134 56525
rect 50186 56513 50192 56525
rect 50515 56516 50573 56522
rect 50515 56513 50527 56516
rect 50186 56485 50527 56513
rect 50186 56473 50192 56485
rect 50515 56482 50527 56485
rect 50561 56482 50573 56516
rect 52912 56513 52918 56525
rect 52873 56485 52918 56513
rect 50515 56476 50573 56482
rect 52912 56473 52918 56485
rect 52970 56473 52976 56525
rect 53296 56473 53302 56525
rect 53354 56513 53360 56525
rect 53779 56516 53837 56522
rect 53779 56513 53791 56516
rect 53354 56485 53791 56513
rect 53354 56473 53360 56485
rect 53779 56482 53791 56485
rect 53825 56482 53837 56516
rect 53779 56476 53837 56482
rect 54352 56473 54358 56525
rect 54410 56513 54416 56525
rect 54547 56516 54605 56522
rect 54547 56513 54559 56516
rect 54410 56485 54559 56513
rect 54410 56473 54416 56485
rect 54547 56482 54559 56485
rect 54593 56482 54605 56516
rect 54547 56476 54605 56482
rect 54928 56473 54934 56525
rect 54986 56513 54992 56525
rect 55315 56516 55373 56522
rect 55315 56513 55327 56516
rect 54986 56485 55327 56513
rect 54986 56473 54992 56485
rect 55315 56482 55327 56485
rect 55361 56482 55373 56516
rect 55984 56513 55990 56525
rect 55945 56485 55990 56513
rect 55315 56476 55373 56482
rect 55984 56473 55990 56485
rect 56042 56473 56048 56525
rect 16528 56399 16534 56451
rect 16586 56439 16592 56451
rect 56752 56439 56758 56451
rect 16586 56411 56758 56439
rect 16586 56399 16592 56411
rect 56752 56399 56758 56411
rect 56810 56399 56816 56451
rect 6931 56368 6989 56374
rect 6931 56334 6943 56368
rect 6977 56365 6989 56368
rect 7219 56368 7277 56374
rect 7219 56365 7231 56368
rect 6977 56337 7231 56365
rect 6977 56334 6989 56337
rect 6931 56328 6989 56334
rect 7219 56334 7231 56337
rect 7265 56365 7277 56368
rect 13744 56365 13750 56377
rect 7265 56337 13750 56365
rect 7265 56334 7277 56337
rect 7219 56328 7277 56334
rect 13744 56325 13750 56337
rect 13802 56325 13808 56377
rect 37459 56368 37517 56374
rect 37459 56334 37471 56368
rect 37505 56365 37517 56368
rect 37747 56368 37805 56374
rect 37747 56365 37759 56368
rect 37505 56337 37759 56365
rect 37505 56334 37517 56337
rect 37459 56328 37517 56334
rect 37747 56334 37759 56337
rect 37793 56365 37805 56368
rect 43312 56365 43318 56377
rect 37793 56337 43318 56365
rect 37793 56334 37805 56337
rect 37747 56328 37805 56334
rect 43312 56325 43318 56337
rect 43370 56325 43376 56377
rect 45139 56368 45197 56374
rect 45139 56334 45151 56368
rect 45185 56365 45197 56368
rect 45185 56337 47534 56365
rect 45185 56334 45197 56337
rect 45139 56328 45197 56334
rect 3760 56251 3766 56303
rect 3818 56291 3824 56303
rect 10099 56294 10157 56300
rect 10099 56291 10111 56294
rect 3818 56263 10111 56291
rect 3818 56251 3824 56263
rect 10099 56260 10111 56263
rect 10145 56291 10157 56294
rect 10291 56294 10349 56300
rect 10291 56291 10303 56294
rect 10145 56263 10303 56291
rect 10145 56260 10157 56263
rect 10099 56254 10157 56260
rect 10291 56260 10303 56263
rect 10337 56260 10349 56294
rect 10291 56254 10349 56260
rect 13555 56294 13613 56300
rect 13555 56260 13567 56294
rect 13601 56291 13613 56294
rect 15184 56291 15190 56303
rect 13601 56263 15190 56291
rect 13601 56260 13613 56263
rect 13555 56254 13613 56260
rect 15184 56251 15190 56263
rect 15242 56251 15248 56303
rect 25843 56294 25901 56300
rect 25843 56260 25855 56294
rect 25889 56291 25901 56294
rect 26131 56294 26189 56300
rect 26131 56291 26143 56294
rect 25889 56263 26143 56291
rect 25889 56260 25901 56263
rect 25843 56254 25901 56260
rect 26131 56260 26143 56263
rect 26177 56291 26189 56294
rect 26416 56291 26422 56303
rect 26177 56263 26422 56291
rect 26177 56260 26189 56263
rect 26131 56254 26189 56260
rect 26416 56251 26422 56263
rect 26474 56251 26480 56303
rect 36016 56251 36022 56303
rect 36074 56291 36080 56303
rect 38803 56294 38861 56300
rect 38803 56291 38815 56294
rect 36074 56263 38815 56291
rect 36074 56251 36080 56263
rect 38803 56260 38815 56263
rect 38849 56260 38861 56294
rect 38803 56254 38861 56260
rect 44275 56294 44333 56300
rect 44275 56260 44287 56294
rect 44321 56291 44333 56294
rect 44321 56263 46814 56291
rect 44321 56260 44333 56263
rect 44275 56254 44333 56260
rect 1744 56217 1750 56229
rect 1705 56189 1750 56217
rect 1744 56177 1750 56189
rect 1802 56177 1808 56229
rect 2512 56217 2518 56229
rect 2473 56189 2518 56217
rect 2512 56177 2518 56189
rect 2570 56177 2576 56229
rect 2995 56220 3053 56226
rect 2995 56186 3007 56220
rect 3041 56217 3053 56220
rect 3283 56220 3341 56226
rect 3283 56217 3295 56220
rect 3041 56189 3295 56217
rect 3041 56186 3053 56189
rect 2995 56180 3053 56186
rect 3283 56186 3295 56189
rect 3329 56217 3341 56220
rect 3376 56217 3382 56229
rect 3329 56189 3382 56217
rect 3329 56186 3341 56189
rect 3283 56180 3341 56186
rect 3376 56177 3382 56189
rect 3434 56177 3440 56229
rect 4243 56220 4301 56226
rect 4243 56186 4255 56220
rect 4289 56217 4301 56220
rect 4531 56220 4589 56226
rect 4531 56217 4543 56220
rect 4289 56189 4543 56217
rect 4289 56186 4301 56189
rect 4243 56180 4301 56186
rect 4531 56186 4543 56189
rect 4577 56217 4589 56220
rect 5200 56217 5206 56229
rect 4577 56189 5206 56217
rect 4577 56186 4589 56189
rect 4531 56180 4589 56186
rect 5200 56177 5206 56189
rect 5258 56177 5264 56229
rect 5584 56217 5590 56229
rect 5545 56189 5590 56217
rect 5584 56177 5590 56189
rect 5642 56177 5648 56229
rect 6352 56217 6358 56229
rect 6313 56189 6358 56217
rect 6352 56177 6358 56189
rect 6410 56177 6416 56229
rect 6448 56177 6454 56229
rect 6506 56217 6512 56229
rect 8563 56220 8621 56226
rect 8563 56217 8575 56220
rect 6506 56189 8575 56217
rect 6506 56177 6512 56189
rect 8563 56186 8575 56189
rect 8609 56186 8621 56220
rect 10768 56217 10774 56229
rect 10729 56189 10774 56217
rect 8563 56180 8621 56186
rect 10768 56177 10774 56189
rect 10826 56217 10832 56229
rect 11155 56220 11213 56226
rect 11155 56217 11167 56220
rect 10826 56189 11167 56217
rect 10826 56177 10832 56189
rect 11155 56186 11167 56189
rect 11201 56186 11213 56220
rect 11920 56217 11926 56229
rect 11881 56189 11926 56217
rect 11155 56180 11213 56186
rect 11920 56177 11926 56189
rect 11978 56177 11984 56229
rect 12403 56220 12461 56226
rect 12403 56186 12415 56220
rect 12449 56217 12461 56220
rect 12688 56217 12694 56229
rect 12449 56189 12694 56217
rect 12449 56186 12461 56189
rect 12403 56180 12461 56186
rect 12688 56177 12694 56189
rect 12746 56177 12752 56229
rect 15088 56177 15094 56229
rect 15146 56217 15152 56229
rect 15571 56220 15629 56226
rect 15146 56189 15191 56217
rect 15146 56177 15152 56189
rect 15571 56186 15583 56220
rect 15617 56217 15629 56220
rect 15760 56217 15766 56229
rect 15617 56189 15766 56217
rect 15617 56186 15629 56189
rect 15571 56180 15629 56186
rect 15760 56177 15766 56189
rect 15818 56177 15824 56229
rect 15859 56220 15917 56226
rect 15859 56186 15871 56220
rect 15905 56186 15917 56220
rect 15859 56180 15917 56186
rect 15376 56103 15382 56155
rect 15434 56143 15440 56155
rect 15874 56143 15902 56180
rect 16624 56177 16630 56229
rect 16682 56217 16688 56229
rect 16819 56220 16877 56226
rect 16819 56217 16831 56220
rect 16682 56189 16831 56217
rect 16682 56177 16688 56189
rect 16819 56186 16831 56189
rect 16865 56217 16877 56220
rect 17107 56220 17165 56226
rect 17107 56217 17119 56220
rect 16865 56189 17119 56217
rect 16865 56186 16877 56189
rect 16819 56180 16877 56186
rect 17107 56186 17119 56189
rect 17153 56186 17165 56220
rect 17107 56180 17165 56186
rect 17971 56220 18029 56226
rect 17971 56186 17983 56220
rect 18017 56217 18029 56220
rect 18256 56217 18262 56229
rect 18017 56189 18262 56217
rect 18017 56186 18029 56189
rect 17971 56180 18029 56186
rect 18256 56177 18262 56189
rect 18314 56177 18320 56229
rect 18736 56217 18742 56229
rect 18697 56189 18742 56217
rect 18736 56177 18742 56189
rect 18794 56217 18800 56229
rect 18931 56220 18989 56226
rect 18931 56217 18943 56220
rect 18794 56189 18943 56217
rect 18794 56177 18800 56189
rect 18931 56186 18943 56189
rect 18977 56186 18989 56220
rect 19984 56217 19990 56229
rect 19945 56189 19990 56217
rect 18931 56180 18989 56186
rect 19984 56177 19990 56189
rect 20042 56217 20048 56229
rect 20275 56220 20333 56226
rect 20275 56217 20287 56220
rect 20042 56189 20287 56217
rect 20042 56177 20048 56189
rect 20275 56186 20287 56189
rect 20321 56186 20333 56220
rect 20275 56180 20333 56186
rect 20371 56220 20429 56226
rect 20371 56186 20383 56220
rect 20417 56186 20429 56220
rect 21040 56217 21046 56229
rect 21001 56189 21046 56217
rect 20371 56180 20429 56186
rect 15434 56115 15902 56143
rect 15434 56103 15440 56115
rect 19504 56103 19510 56155
rect 19562 56143 19568 56155
rect 20386 56143 20414 56180
rect 21040 56177 21046 56189
rect 21098 56217 21104 56229
rect 21427 56220 21485 56226
rect 21427 56217 21439 56220
rect 21098 56189 21439 56217
rect 21098 56177 21104 56189
rect 21427 56186 21439 56189
rect 21473 56186 21485 56220
rect 21808 56217 21814 56229
rect 21769 56189 21814 56217
rect 21427 56180 21485 56186
rect 21808 56177 21814 56189
rect 21866 56217 21872 56229
rect 22195 56220 22253 56226
rect 22195 56217 22207 56220
rect 21866 56189 22207 56217
rect 21866 56177 21872 56189
rect 22195 56186 22207 56189
rect 22241 56186 22253 56220
rect 22195 56180 22253 56186
rect 22960 56177 22966 56229
rect 23018 56217 23024 56229
rect 24115 56220 24173 56226
rect 23018 56189 23063 56217
rect 23018 56177 23024 56189
rect 24115 56186 24127 56220
rect 24161 56217 24173 56220
rect 24304 56217 24310 56229
rect 24161 56189 24310 56217
rect 24161 56186 24173 56189
rect 24115 56180 24173 56186
rect 24304 56177 24310 56189
rect 24362 56177 24368 56229
rect 26512 56217 26518 56229
rect 26473 56189 26518 56217
rect 26512 56177 26518 56189
rect 26570 56217 26576 56229
rect 26803 56220 26861 56226
rect 26803 56217 26815 56220
rect 26570 56189 26815 56217
rect 26570 56177 26576 56189
rect 26803 56186 26815 56189
rect 26849 56186 26861 56220
rect 26803 56180 26861 56186
rect 27475 56220 27533 56226
rect 27475 56186 27487 56220
rect 27521 56217 27533 56220
rect 27664 56217 27670 56229
rect 27521 56189 27670 56217
rect 27521 56186 27533 56189
rect 27475 56180 27533 56186
rect 27664 56177 27670 56189
rect 27722 56177 27728 56229
rect 28144 56217 28150 56229
rect 28105 56189 28150 56217
rect 28144 56177 28150 56189
rect 28202 56217 28208 56229
rect 28435 56220 28493 56226
rect 28435 56217 28447 56220
rect 28202 56189 28447 56217
rect 28202 56177 28208 56189
rect 28435 56186 28447 56189
rect 28481 56186 28493 56220
rect 28435 56180 28493 56186
rect 29395 56220 29453 56226
rect 29395 56186 29407 56220
rect 29441 56217 29453 56220
rect 29584 56217 29590 56229
rect 29441 56189 29590 56217
rect 29441 56186 29453 56189
rect 29395 56180 29453 56186
rect 29584 56177 29590 56189
rect 29642 56177 29648 56229
rect 30928 56217 30934 56229
rect 30889 56189 30934 56217
rect 30928 56177 30934 56189
rect 30986 56177 30992 56229
rect 31312 56217 31318 56229
rect 31273 56189 31318 56217
rect 31312 56177 31318 56189
rect 31370 56217 31376 56229
rect 31603 56220 31661 56226
rect 31603 56217 31615 56220
rect 31370 56189 31615 56217
rect 31370 56177 31376 56189
rect 31603 56186 31615 56189
rect 31649 56186 31661 56220
rect 31603 56180 31661 56186
rect 31699 56220 31757 56226
rect 31699 56186 31711 56220
rect 31745 56186 31757 56220
rect 31699 56180 31757 56186
rect 32179 56220 32237 56226
rect 32179 56186 32191 56220
rect 32225 56217 32237 56220
rect 32464 56217 32470 56229
rect 32225 56189 32470 56217
rect 32225 56186 32237 56189
rect 32179 56180 32237 56186
rect 19562 56115 20414 56143
rect 19562 56103 19568 56115
rect 31216 56103 31222 56155
rect 31274 56143 31280 56155
rect 31714 56143 31742 56180
rect 32464 56177 32470 56189
rect 32522 56177 32528 56229
rect 32848 56217 32854 56229
rect 32809 56189 32854 56217
rect 32848 56177 32854 56189
rect 32906 56217 32912 56229
rect 33139 56220 33197 56226
rect 33139 56217 33151 56220
rect 32906 56189 33151 56217
rect 32906 56177 32912 56189
rect 33139 56186 33151 56189
rect 33185 56186 33197 56220
rect 33139 56180 33197 56186
rect 33235 56220 33293 56226
rect 33235 56186 33247 56220
rect 33281 56186 33293 56220
rect 34000 56217 34006 56229
rect 33961 56189 34006 56217
rect 33235 56180 33293 56186
rect 31274 56115 31742 56143
rect 31274 56103 31280 56115
rect 32752 56103 32758 56155
rect 32810 56143 32816 56155
rect 33250 56143 33278 56180
rect 34000 56177 34006 56189
rect 34058 56177 34064 56229
rect 34768 56217 34774 56229
rect 34729 56189 34774 56217
rect 34768 56177 34774 56189
rect 34826 56177 34832 56229
rect 35824 56217 35830 56229
rect 35785 56189 35830 56217
rect 35824 56177 35830 56189
rect 35882 56217 35888 56229
rect 36115 56220 36173 56226
rect 36115 56217 36127 56220
rect 35882 56189 36127 56217
rect 35882 56177 35888 56189
rect 36115 56186 36127 56189
rect 36161 56186 36173 56220
rect 36115 56180 36173 56186
rect 36211 56220 36269 56226
rect 36211 56186 36223 56220
rect 36257 56186 36269 56220
rect 36592 56217 36598 56229
rect 36553 56189 36598 56217
rect 36211 56180 36269 56186
rect 32810 56115 33278 56143
rect 32810 56103 32816 56115
rect 35440 56103 35446 56155
rect 35498 56143 35504 56155
rect 36226 56143 36254 56180
rect 36592 56177 36598 56189
rect 36650 56217 36656 56229
rect 36883 56220 36941 56226
rect 36883 56217 36895 56220
rect 36650 56189 36895 56217
rect 36650 56177 36656 56189
rect 36883 56186 36895 56189
rect 36929 56186 36941 56220
rect 40240 56217 40246 56229
rect 40201 56189 40246 56217
rect 36883 56180 36941 56186
rect 40240 56177 40246 56189
rect 40298 56177 40304 56229
rect 41971 56220 42029 56226
rect 41971 56186 41983 56220
rect 42017 56217 42029 56220
rect 42064 56217 42070 56229
rect 42017 56189 42070 56217
rect 42017 56186 42029 56189
rect 41971 56180 42029 56186
rect 42064 56177 42070 56189
rect 42122 56177 42128 56229
rect 42352 56217 42358 56229
rect 42313 56189 42358 56217
rect 42352 56177 42358 56189
rect 42410 56217 42416 56229
rect 42643 56220 42701 56226
rect 42643 56217 42655 56220
rect 42410 56189 42655 56217
rect 42410 56177 42416 56189
rect 42643 56186 42655 56189
rect 42689 56186 42701 56220
rect 42643 56180 42701 56186
rect 43219 56220 43277 56226
rect 43219 56186 43231 56220
rect 43265 56217 43277 56220
rect 43408 56217 43414 56229
rect 43265 56189 43414 56217
rect 43265 56186 43277 56189
rect 43219 56180 43277 56186
rect 43408 56177 43414 56189
rect 43466 56177 43472 56229
rect 46483 56220 46541 56226
rect 46483 56186 46495 56220
rect 46529 56217 46541 56220
rect 46672 56217 46678 56229
rect 46529 56189 46678 56217
rect 46529 56186 46541 56189
rect 46483 56180 46541 56186
rect 46672 56177 46678 56189
rect 46730 56177 46736 56229
rect 46786 56217 46814 56263
rect 46864 56251 46870 56303
rect 46922 56291 46928 56303
rect 46963 56294 47021 56300
rect 46963 56291 46975 56294
rect 46922 56263 46975 56291
rect 46922 56251 46928 56263
rect 46963 56260 46975 56263
rect 47009 56260 47021 56294
rect 47506 56291 47534 56337
rect 49168 56325 49174 56377
rect 49226 56365 49232 56377
rect 52051 56368 52109 56374
rect 52051 56365 52063 56368
rect 49226 56337 52063 56365
rect 49226 56325 49232 56337
rect 52051 56334 52063 56337
rect 52097 56334 52109 56368
rect 52051 56328 52109 56334
rect 52144 56325 52150 56377
rect 52202 56365 52208 56377
rect 56083 56368 56141 56374
rect 56083 56365 56095 56368
rect 52202 56337 56095 56365
rect 52202 56325 52208 56337
rect 56083 56334 56095 56337
rect 56129 56334 56141 56368
rect 56083 56328 56141 56334
rect 47506 56263 49598 56291
rect 46963 56254 47021 56260
rect 47920 56217 47926 56229
rect 46786 56189 47926 56217
rect 47920 56177 47926 56189
rect 47978 56177 47984 56229
rect 48208 56217 48214 56229
rect 48169 56189 48214 56217
rect 48208 56177 48214 56189
rect 48266 56177 48272 56229
rect 48691 56220 48749 56226
rect 48691 56186 48703 56220
rect 48737 56217 48749 56220
rect 48880 56217 48886 56229
rect 48737 56189 48886 56217
rect 48737 56186 48749 56189
rect 48691 56180 48749 56186
rect 48880 56177 48886 56189
rect 48938 56177 48944 56229
rect 48979 56220 49037 56226
rect 48979 56186 48991 56220
rect 49025 56186 49037 56220
rect 49570 56217 49598 56263
rect 49648 56251 49654 56303
rect 49706 56291 49712 56303
rect 50611 56294 50669 56300
rect 50611 56291 50623 56294
rect 49706 56263 50623 56291
rect 49706 56251 49712 56263
rect 50611 56260 50623 56263
rect 50657 56260 50669 56294
rect 54352 56291 54358 56303
rect 50611 56254 50669 56260
rect 51874 56263 54358 56291
rect 49570 56189 49790 56217
rect 48979 56180 49037 56186
rect 35498 56115 36254 56143
rect 35498 56103 35504 56115
rect 37072 56103 37078 56155
rect 37130 56143 37136 56155
rect 40816 56143 40822 56155
rect 37130 56115 40822 56143
rect 37130 56103 37136 56115
rect 40816 56103 40822 56115
rect 40874 56103 40880 56155
rect 48592 56103 48598 56155
rect 48650 56143 48656 56155
rect 48994 56143 49022 56180
rect 48650 56115 49022 56143
rect 49762 56143 49790 56189
rect 49840 56177 49846 56229
rect 49898 56217 49904 56229
rect 51874 56217 51902 56263
rect 54352 56251 54358 56263
rect 54410 56251 54416 56303
rect 57811 56294 57869 56300
rect 57811 56260 57823 56294
rect 57857 56291 57869 56294
rect 58576 56291 58582 56303
rect 57857 56263 58582 56291
rect 57857 56260 57869 56263
rect 57811 56254 57869 56260
rect 58576 56251 58582 56263
rect 58634 56251 58640 56303
rect 49898 56189 49943 56217
rect 50050 56189 51902 56217
rect 51955 56220 52013 56226
rect 49898 56177 49904 56189
rect 50050 56143 50078 56189
rect 51955 56186 51967 56220
rect 52001 56186 52013 56220
rect 53008 56217 53014 56229
rect 52969 56189 53014 56217
rect 51955 56180 52013 56186
rect 49762 56115 50078 56143
rect 48650 56103 48656 56115
rect 51184 56103 51190 56155
rect 51242 56143 51248 56155
rect 51970 56143 51998 56180
rect 53008 56177 53014 56189
rect 53066 56177 53072 56229
rect 53392 56217 53398 56229
rect 53353 56189 53398 56217
rect 53392 56177 53398 56189
rect 53450 56217 53456 56229
rect 53683 56220 53741 56226
rect 53683 56217 53695 56220
rect 53450 56189 53695 56217
rect 53450 56177 53456 56189
rect 53683 56186 53695 56189
rect 53729 56186 53741 56220
rect 53683 56180 53741 56186
rect 54259 56220 54317 56226
rect 54259 56186 54271 56220
rect 54305 56217 54317 56220
rect 54448 56217 54454 56229
rect 54305 56189 54454 56217
rect 54305 56186 54317 56189
rect 54259 56180 54317 56186
rect 54448 56177 54454 56189
rect 54506 56177 54512 56229
rect 55027 56220 55085 56226
rect 55027 56186 55039 56220
rect 55073 56217 55085 56220
rect 55219 56220 55277 56226
rect 55219 56217 55231 56220
rect 55073 56189 55231 56217
rect 55073 56186 55085 56189
rect 55027 56180 55085 56186
rect 55219 56186 55231 56189
rect 55265 56217 55277 56220
rect 55504 56217 55510 56229
rect 55265 56189 55510 56217
rect 55265 56186 55277 56189
rect 55219 56180 55277 56186
rect 55504 56177 55510 56189
rect 55562 56177 55568 56229
rect 51242 56115 51998 56143
rect 51242 56103 51248 56115
rect 1152 55970 58848 55992
rect 1152 55918 4294 55970
rect 4346 55918 4358 55970
rect 4410 55918 4422 55970
rect 4474 55918 4486 55970
rect 4538 55918 35014 55970
rect 35066 55918 35078 55970
rect 35130 55918 35142 55970
rect 35194 55918 35206 55970
rect 35258 55918 58848 55970
rect 1152 55896 58848 55918
rect 17971 55776 18029 55782
rect 17971 55742 17983 55776
rect 18017 55773 18029 55776
rect 18259 55776 18317 55782
rect 18259 55773 18271 55776
rect 18017 55745 18271 55773
rect 18017 55742 18029 55745
rect 17971 55736 18029 55742
rect 18259 55742 18271 55745
rect 18305 55773 18317 55776
rect 26320 55773 26326 55785
rect 18305 55745 26326 55773
rect 18305 55742 18317 55745
rect 18259 55736 18317 55742
rect 26320 55733 26326 55745
rect 26378 55733 26384 55785
rect 1168 55659 1174 55711
rect 1226 55699 1232 55711
rect 1651 55702 1709 55708
rect 1651 55699 1663 55702
rect 1226 55671 1663 55699
rect 1226 55659 1232 55671
rect 1651 55668 1663 55671
rect 1697 55668 1709 55702
rect 1651 55662 1709 55668
rect 4435 55702 4493 55708
rect 4435 55668 4447 55702
rect 4481 55699 4493 55702
rect 4624 55699 4630 55711
rect 4481 55671 4630 55699
rect 4481 55668 4493 55671
rect 4435 55662 4493 55668
rect 4624 55659 4630 55671
rect 4682 55659 4688 55711
rect 7504 55659 7510 55711
rect 7562 55699 7568 55711
rect 7603 55702 7661 55708
rect 7603 55699 7615 55702
rect 7562 55671 7615 55699
rect 7562 55659 7568 55671
rect 7603 55668 7615 55671
rect 7649 55668 7661 55702
rect 7603 55662 7661 55668
rect 9136 55659 9142 55711
rect 9194 55699 9200 55711
rect 9331 55702 9389 55708
rect 9331 55699 9343 55702
rect 9194 55671 9343 55699
rect 9194 55659 9200 55671
rect 9331 55668 9343 55671
rect 9377 55668 9389 55702
rect 9331 55662 9389 55668
rect 13840 55659 13846 55711
rect 13898 55699 13904 55711
rect 13939 55702 13997 55708
rect 13939 55699 13951 55702
rect 13898 55671 13951 55699
rect 13898 55659 13904 55671
rect 13939 55668 13951 55671
rect 13985 55668 13997 55702
rect 13939 55662 13997 55668
rect 20176 55659 20182 55711
rect 20234 55699 20240 55711
rect 20275 55702 20333 55708
rect 20275 55699 20287 55702
rect 20234 55671 20287 55699
rect 20234 55659 20240 55671
rect 20275 55668 20287 55671
rect 20321 55668 20333 55702
rect 20275 55662 20333 55668
rect 23344 55659 23350 55711
rect 23402 55699 23408 55711
rect 23539 55702 23597 55708
rect 23539 55699 23551 55702
rect 23402 55671 23551 55699
rect 23402 55659 23408 55671
rect 23539 55668 23551 55671
rect 23585 55668 23597 55702
rect 23539 55662 23597 55668
rect 24880 55659 24886 55711
rect 24938 55699 24944 55711
rect 25075 55702 25133 55708
rect 25075 55699 25087 55702
rect 24938 55671 25087 55699
rect 24938 55659 24944 55671
rect 25075 55668 25087 55671
rect 25121 55668 25133 55702
rect 25075 55662 25133 55668
rect 39088 55659 39094 55711
rect 39146 55699 39152 55711
rect 39283 55702 39341 55708
rect 39283 55699 39295 55702
rect 39146 55671 39295 55699
rect 39146 55659 39152 55671
rect 39283 55668 39295 55671
rect 39329 55668 39341 55702
rect 39283 55662 39341 55668
rect 40720 55659 40726 55711
rect 40778 55699 40784 55711
rect 40819 55702 40877 55708
rect 40819 55699 40831 55702
rect 40778 55671 40831 55699
rect 40778 55659 40784 55671
rect 40819 55668 40831 55671
rect 40865 55668 40877 55702
rect 40819 55662 40877 55668
rect 45424 55659 45430 55711
rect 45482 55699 45488 55711
rect 45619 55702 45677 55708
rect 45619 55699 45631 55702
rect 45482 55671 45631 55699
rect 45482 55659 45488 55671
rect 45619 55668 45631 55671
rect 45665 55668 45677 55702
rect 45619 55662 45677 55668
rect 46960 55659 46966 55711
rect 47018 55699 47024 55711
rect 47155 55702 47213 55708
rect 47155 55699 47167 55702
rect 47018 55671 47167 55699
rect 47018 55659 47024 55671
rect 47155 55668 47167 55671
rect 47201 55668 47213 55702
rect 47155 55662 47213 55668
rect 51760 55659 51766 55711
rect 51818 55699 51824 55711
rect 51955 55702 52013 55708
rect 51955 55699 51967 55702
rect 51818 55671 51967 55699
rect 51818 55659 51824 55671
rect 51955 55668 51967 55671
rect 52001 55668 52013 55702
rect 51955 55662 52013 55668
rect 56464 55659 56470 55711
rect 56522 55699 56528 55711
rect 56563 55702 56621 55708
rect 56563 55699 56575 55702
rect 56522 55671 56575 55699
rect 56522 55659 56528 55671
rect 56563 55668 56575 55671
rect 56609 55668 56621 55702
rect 56563 55662 56621 55668
rect 57520 55659 57526 55711
rect 57578 55699 57584 55711
rect 57715 55702 57773 55708
rect 57715 55699 57727 55702
rect 57578 55671 57727 55699
rect 57578 55659 57584 55671
rect 57715 55668 57727 55671
rect 57761 55668 57773 55702
rect 57715 55662 57773 55668
rect 21427 55628 21485 55634
rect 21427 55594 21439 55628
rect 21473 55625 21485 55628
rect 36016 55625 36022 55637
rect 21473 55597 36022 55625
rect 21473 55594 21485 55597
rect 21427 55588 21485 55594
rect 36016 55585 36022 55597
rect 36074 55585 36080 55637
rect 54259 55628 54317 55634
rect 54259 55625 54271 55628
rect 47506 55597 54271 55625
rect 1747 55554 1805 55560
rect 1747 55520 1759 55554
rect 1793 55520 1805 55554
rect 1747 55514 1805 55520
rect 4243 55554 4301 55560
rect 4243 55520 4255 55554
rect 4289 55551 4301 55554
rect 4531 55554 4589 55560
rect 4531 55551 4543 55554
rect 4289 55523 4543 55551
rect 4289 55520 4301 55523
rect 4243 55514 4301 55520
rect 4531 55520 4543 55523
rect 4577 55551 4589 55554
rect 4624 55551 4630 55563
rect 4577 55523 4630 55551
rect 4577 55520 4589 55523
rect 4531 55514 4589 55520
rect 1762 55403 1790 55514
rect 4624 55511 4630 55523
rect 4682 55511 4688 55563
rect 7696 55551 7702 55563
rect 7657 55523 7702 55551
rect 7696 55511 7702 55523
rect 7754 55511 7760 55563
rect 8179 55554 8237 55560
rect 8179 55520 8191 55554
rect 8225 55551 8237 55554
rect 8464 55551 8470 55563
rect 8225 55523 8470 55551
rect 8225 55520 8237 55523
rect 8179 55514 8237 55520
rect 8464 55511 8470 55523
rect 8522 55511 8528 55563
rect 9043 55554 9101 55560
rect 9043 55520 9055 55554
rect 9089 55551 9101 55554
rect 9232 55551 9238 55563
rect 9089 55523 9238 55551
rect 9089 55520 9101 55523
rect 9043 55514 9101 55520
rect 9232 55511 9238 55523
rect 9290 55511 9296 55563
rect 13747 55554 13805 55560
rect 13747 55520 13759 55554
rect 13793 55551 13805 55554
rect 14032 55551 14038 55563
rect 13793 55523 14038 55551
rect 13793 55520 13805 55523
rect 13747 55514 13805 55520
rect 14032 55511 14038 55523
rect 14090 55511 14096 55563
rect 20371 55554 20429 55560
rect 20371 55520 20383 55554
rect 20417 55551 20429 55554
rect 20464 55551 20470 55563
rect 20417 55523 20470 55551
rect 20417 55520 20429 55523
rect 20371 55514 20429 55520
rect 20464 55511 20470 55523
rect 20522 55511 20528 55563
rect 23251 55554 23309 55560
rect 23251 55520 23263 55554
rect 23297 55551 23309 55554
rect 23440 55551 23446 55563
rect 23297 55523 23446 55551
rect 23297 55520 23309 55523
rect 23251 55514 23309 55520
rect 23440 55511 23446 55523
rect 23498 55511 23504 55563
rect 24979 55554 25037 55560
rect 24979 55551 24991 55554
rect 24706 55523 24991 55551
rect 24706 55415 24734 55523
rect 24979 55520 24991 55523
rect 25025 55520 25037 55554
rect 28915 55554 28973 55560
rect 28915 55551 28927 55554
rect 24979 55514 25037 55520
rect 28834 55523 28927 55551
rect 1840 55403 1846 55415
rect 1762 55375 1846 55403
rect 1840 55363 1846 55375
rect 1898 55403 1904 55415
rect 1939 55406 1997 55412
rect 1939 55403 1951 55406
rect 1898 55375 1951 55403
rect 1898 55363 1904 55375
rect 1939 55372 1951 55375
rect 1985 55372 1997 55406
rect 24688 55403 24694 55415
rect 24649 55375 24694 55403
rect 1939 55366 1997 55372
rect 24688 55363 24694 55375
rect 24746 55363 24752 55415
rect 28624 55363 28630 55415
rect 28682 55403 28688 55415
rect 28834 55412 28862 55523
rect 28915 55520 28927 55523
rect 28961 55520 28973 55554
rect 30163 55554 30221 55560
rect 30163 55551 30175 55554
rect 28915 55514 28973 55520
rect 29794 55523 30175 55551
rect 29794 55415 29822 55523
rect 30163 55520 30175 55523
rect 30209 55520 30221 55554
rect 30163 55514 30221 55520
rect 38896 55511 38902 55563
rect 38954 55551 38960 55563
rect 39187 55554 39245 55560
rect 39187 55551 39199 55554
rect 38954 55523 39199 55551
rect 38954 55511 38960 55523
rect 39187 55520 39199 55523
rect 39233 55520 39245 55554
rect 40912 55551 40918 55563
rect 40873 55523 40918 55551
rect 39187 55514 39245 55520
rect 40912 55511 40918 55523
rect 40970 55511 40976 55563
rect 45232 55511 45238 55563
rect 45290 55551 45296 55563
rect 45523 55554 45581 55560
rect 45523 55551 45535 55554
rect 45290 55523 45535 55551
rect 45290 55511 45296 55523
rect 45523 55520 45535 55523
rect 45569 55520 45581 55554
rect 45523 55514 45581 55520
rect 46480 55511 46486 55563
rect 46538 55551 46544 55563
rect 47059 55554 47117 55560
rect 47059 55551 47071 55554
rect 46538 55523 47071 55551
rect 46538 55511 46544 55523
rect 47059 55520 47071 55523
rect 47105 55520 47117 55554
rect 47059 55514 47117 55520
rect 32368 55437 32374 55489
rect 32426 55477 32432 55489
rect 47506 55477 47534 55597
rect 54259 55594 54271 55597
rect 54305 55625 54317 55628
rect 54451 55628 54509 55634
rect 54451 55625 54463 55628
rect 54305 55597 54463 55625
rect 54305 55594 54317 55597
rect 54259 55588 54317 55594
rect 54451 55594 54463 55597
rect 54497 55594 54509 55628
rect 54451 55588 54509 55594
rect 50515 55554 50573 55560
rect 50515 55520 50527 55554
rect 50561 55520 50573 55554
rect 51859 55554 51917 55560
rect 51859 55551 51871 55554
rect 50515 55514 50573 55520
rect 51586 55523 51871 55551
rect 32426 55449 47534 55477
rect 32426 55437 32432 55449
rect 28819 55406 28877 55412
rect 28819 55403 28831 55406
rect 28682 55375 28831 55403
rect 28682 55363 28688 55375
rect 28819 55372 28831 55375
rect 28865 55372 28877 55406
rect 29776 55403 29782 55415
rect 29737 55375 29782 55403
rect 28819 55366 28877 55372
rect 29776 55363 29782 55375
rect 29834 55363 29840 55415
rect 38896 55403 38902 55415
rect 38857 55375 38902 55403
rect 38896 55363 38902 55375
rect 38954 55363 38960 55415
rect 45232 55403 45238 55415
rect 45193 55375 45238 55403
rect 45232 55363 45238 55375
rect 45290 55363 45296 55415
rect 46480 55363 46486 55415
rect 46538 55403 46544 55415
rect 46771 55406 46829 55412
rect 46771 55403 46783 55406
rect 46538 55375 46783 55403
rect 46538 55363 46544 55375
rect 46771 55372 46783 55375
rect 46817 55372 46829 55406
rect 46771 55366 46829 55372
rect 50419 55406 50477 55412
rect 50419 55372 50431 55406
rect 50465 55403 50477 55406
rect 50530 55403 50558 55514
rect 51586 55415 51614 55523
rect 51859 55520 51871 55523
rect 51905 55520 51917 55554
rect 55795 55554 55853 55560
rect 55795 55551 55807 55554
rect 51859 55514 51917 55520
rect 55618 55523 55807 55551
rect 55618 55415 55646 55523
rect 55795 55520 55807 55523
rect 55841 55520 55853 55554
rect 55795 55514 55853 55520
rect 56371 55554 56429 55560
rect 56371 55520 56383 55554
rect 56417 55551 56429 55554
rect 56656 55551 56662 55563
rect 56417 55523 56662 55551
rect 56417 55520 56429 55523
rect 56371 55514 56429 55520
rect 56656 55511 56662 55523
rect 56714 55511 56720 55563
rect 57427 55554 57485 55560
rect 57427 55520 57439 55554
rect 57473 55551 57485 55554
rect 57520 55551 57526 55563
rect 57473 55523 57526 55551
rect 57473 55520 57485 55523
rect 57427 55514 57485 55520
rect 57520 55511 57526 55523
rect 57578 55551 57584 55563
rect 57619 55554 57677 55560
rect 57619 55551 57631 55554
rect 57578 55523 57631 55551
rect 57578 55511 57584 55523
rect 57619 55520 57631 55523
rect 57665 55520 57677 55554
rect 57619 55514 57677 55520
rect 50704 55403 50710 55415
rect 50465 55375 50710 55403
rect 50465 55372 50477 55375
rect 50419 55366 50477 55372
rect 50704 55363 50710 55375
rect 50762 55363 50768 55415
rect 51568 55403 51574 55415
rect 51529 55375 51574 55403
rect 51568 55363 51574 55375
rect 51626 55363 51632 55415
rect 55600 55403 55606 55415
rect 55561 55375 55606 55403
rect 55600 55363 55606 55375
rect 55658 55363 55664 55415
rect 1152 55304 58848 55326
rect 1152 55252 19654 55304
rect 19706 55252 19718 55304
rect 19770 55252 19782 55304
rect 19834 55252 19846 55304
rect 19898 55252 50374 55304
rect 50426 55252 50438 55304
rect 50490 55252 50502 55304
rect 50554 55252 50566 55304
rect 50618 55252 58848 55304
rect 1152 55230 58848 55252
rect 12016 55141 12022 55193
rect 12074 55181 12080 55193
rect 24688 55181 24694 55193
rect 12074 55153 24694 55181
rect 12074 55141 12080 55153
rect 24688 55141 24694 55153
rect 24746 55141 24752 55193
rect 26704 55181 26710 55193
rect 26665 55153 26710 55181
rect 26704 55141 26710 55153
rect 26762 55141 26768 55193
rect 57811 55184 57869 55190
rect 57811 55150 57823 55184
rect 57857 55181 57869 55184
rect 59152 55181 59158 55193
rect 57857 55153 59158 55181
rect 57857 55150 57869 55153
rect 57811 55144 57869 55150
rect 59152 55141 59158 55153
rect 59210 55141 59216 55193
rect 30160 55067 30166 55119
rect 30218 55107 30224 55119
rect 55600 55107 55606 55119
rect 30218 55079 55606 55107
rect 30218 55067 30224 55079
rect 55600 55067 55606 55079
rect 55658 55067 55664 55119
rect 20560 54993 20566 55045
rect 20618 55033 20624 55045
rect 32368 55033 32374 55045
rect 20618 55005 32374 55033
rect 20618 54993 20624 55005
rect 32368 54993 32374 55005
rect 32426 54993 32432 55045
rect 54352 54993 54358 55045
rect 54410 55033 54416 55045
rect 54451 55036 54509 55042
rect 54451 55033 54463 55036
rect 54410 55005 54463 55033
rect 54410 54993 54416 55005
rect 54451 55002 54463 55005
rect 54497 55002 54509 55036
rect 54451 54996 54509 55002
rect 5296 54919 5302 54971
rect 5354 54959 5360 54971
rect 28624 54959 28630 54971
rect 5354 54931 28630 54959
rect 5354 54919 5360 54931
rect 28624 54919 28630 54931
rect 28682 54919 28688 54971
rect 36691 54962 36749 54968
rect 36691 54928 36703 54962
rect 36737 54959 36749 54962
rect 36784 54959 36790 54971
rect 36737 54931 36790 54959
rect 36737 54928 36749 54931
rect 36691 54922 36749 54928
rect 36784 54919 36790 54931
rect 36842 54919 36848 54971
rect 57904 54885 57910 54897
rect 27394 54857 37454 54885
rect 57865 54857 57910 54885
rect 8464 54771 8470 54823
rect 8522 54811 8528 54823
rect 27394 54811 27422 54857
rect 8522 54783 27422 54811
rect 37426 54811 37454 54857
rect 57904 54845 57910 54857
rect 57962 54845 57968 54897
rect 51088 54811 51094 54823
rect 37426 54783 51094 54811
rect 8522 54771 8528 54783
rect 51088 54771 51094 54783
rect 51146 54771 51152 54823
rect 22099 54740 22157 54746
rect 22099 54706 22111 54740
rect 22145 54737 22157 54740
rect 40912 54737 40918 54749
rect 22145 54709 40918 54737
rect 22145 54706 22157 54709
rect 22099 54700 22157 54706
rect 40912 54697 40918 54709
rect 40970 54697 40976 54749
rect 46576 54737 46582 54749
rect 46537 54709 46582 54737
rect 46576 54697 46582 54709
rect 46634 54737 46640 54749
rect 46771 54740 46829 54746
rect 46771 54737 46783 54740
rect 46634 54709 46783 54737
rect 46634 54697 46640 54709
rect 46771 54706 46783 54709
rect 46817 54706 46829 54740
rect 46771 54700 46829 54706
rect 1152 54638 58848 54660
rect 1152 54586 4294 54638
rect 4346 54586 4358 54638
rect 4410 54586 4422 54638
rect 4474 54586 4486 54638
rect 4538 54586 35014 54638
rect 35066 54586 35078 54638
rect 35130 54586 35142 54638
rect 35194 54586 35206 54638
rect 35258 54586 58848 54638
rect 1152 54564 58848 54586
rect 57907 54370 57965 54376
rect 57907 54336 57919 54370
rect 57953 54367 57965 54370
rect 58096 54367 58102 54379
rect 57953 54339 58102 54367
rect 57953 54336 57965 54339
rect 57907 54330 57965 54336
rect 58096 54327 58102 54339
rect 58154 54327 58160 54379
rect 30835 54222 30893 54228
rect 30835 54188 30847 54222
rect 30881 54219 30893 54222
rect 31123 54222 31181 54228
rect 31123 54219 31135 54222
rect 30881 54191 31135 54219
rect 30881 54188 30893 54191
rect 30835 54182 30893 54188
rect 31123 54188 31135 54191
rect 31169 54219 31181 54222
rect 33616 54219 33622 54231
rect 31169 54191 33622 54219
rect 31169 54188 31181 54191
rect 31123 54182 31181 54188
rect 33616 54179 33622 54191
rect 33674 54179 33680 54231
rect 42355 54222 42413 54228
rect 42355 54188 42367 54222
rect 42401 54188 42413 54222
rect 42355 54182 42413 54188
rect 44947 54222 45005 54228
rect 44947 54188 44959 54222
rect 44993 54219 45005 54222
rect 45235 54222 45293 54228
rect 45235 54219 45247 54222
rect 44993 54191 45247 54219
rect 44993 54188 45005 54191
rect 44947 54182 45005 54188
rect 45235 54188 45247 54191
rect 45281 54219 45293 54222
rect 49744 54219 49750 54231
rect 45281 54191 49750 54219
rect 45281 54188 45293 54191
rect 45235 54182 45293 54188
rect 2128 54105 2134 54157
rect 2186 54145 2192 54157
rect 42163 54148 42221 54154
rect 42163 54145 42175 54148
rect 2186 54117 42175 54145
rect 2186 54105 2192 54117
rect 42163 54114 42175 54117
rect 42209 54145 42221 54148
rect 42370 54145 42398 54182
rect 49744 54179 49750 54191
rect 49802 54179 49808 54231
rect 57811 54222 57869 54228
rect 57811 54219 57823 54222
rect 57634 54191 57823 54219
rect 42209 54117 42398 54145
rect 42209 54114 42221 54117
rect 42163 54108 42221 54114
rect 57634 54083 57662 54191
rect 57811 54188 57823 54191
rect 57857 54188 57869 54222
rect 57811 54182 57869 54188
rect 2419 54074 2477 54080
rect 2419 54040 2431 54074
rect 2465 54071 2477 54074
rect 34000 54071 34006 54083
rect 2465 54043 34006 54071
rect 2465 54040 2477 54043
rect 2419 54034 2477 54040
rect 34000 54031 34006 54043
rect 34058 54031 34064 54083
rect 57616 54031 57622 54083
rect 57674 54071 57680 54083
rect 57674 54043 57719 54071
rect 57674 54031 57680 54043
rect 1152 53972 58848 53994
rect 1152 53920 19654 53972
rect 19706 53920 19718 53972
rect 19770 53920 19782 53972
rect 19834 53920 19846 53972
rect 19898 53920 50374 53972
rect 50426 53920 50438 53972
rect 50490 53920 50502 53972
rect 50554 53920 50566 53972
rect 50618 53920 58848 53972
rect 1152 53898 58848 53920
rect 57907 53852 57965 53858
rect 57907 53818 57919 53852
rect 57953 53849 57965 53852
rect 59632 53849 59638 53861
rect 57953 53821 59638 53849
rect 57953 53818 57965 53821
rect 57907 53812 57965 53818
rect 59632 53809 59638 53821
rect 59690 53809 59696 53861
rect 7891 53556 7949 53562
rect 7891 53522 7903 53556
rect 7937 53553 7949 53556
rect 8179 53556 8237 53562
rect 8179 53553 8191 53556
rect 7937 53525 8191 53553
rect 7937 53522 7949 53525
rect 7891 53516 7949 53522
rect 8179 53522 8191 53525
rect 8225 53553 8237 53556
rect 57811 53556 57869 53562
rect 57811 53553 57823 53556
rect 8225 53525 17294 53553
rect 8225 53522 8237 53525
rect 8179 53516 8237 53522
rect 17266 53479 17294 53525
rect 57730 53525 57823 53553
rect 26128 53479 26134 53491
rect 7186 53451 8510 53479
rect 17266 53451 26134 53479
rect 5203 53408 5261 53414
rect 5203 53374 5215 53408
rect 5249 53405 5261 53408
rect 5491 53408 5549 53414
rect 5491 53405 5503 53408
rect 5249 53377 5503 53405
rect 5249 53374 5261 53377
rect 5203 53368 5261 53374
rect 5491 53374 5503 53377
rect 5537 53405 5549 53408
rect 7186 53405 7214 53451
rect 5537 53377 7214 53405
rect 8482 53405 8510 53451
rect 26128 53439 26134 53451
rect 26186 53439 26192 53491
rect 57730 53417 57758 53525
rect 57811 53522 57823 53525
rect 57857 53522 57869 53556
rect 57811 53516 57869 53522
rect 57328 53405 57334 53417
rect 8482 53377 57334 53405
rect 5537 53374 5549 53377
rect 5491 53368 5549 53374
rect 57328 53365 57334 53377
rect 57386 53365 57392 53417
rect 57619 53408 57677 53414
rect 57619 53374 57631 53408
rect 57665 53405 57677 53408
rect 57712 53405 57718 53417
rect 57665 53377 57718 53405
rect 57665 53374 57677 53377
rect 57619 53368 57677 53374
rect 57712 53365 57718 53377
rect 57770 53365 57776 53417
rect 1152 53306 58848 53328
rect 1152 53254 4294 53306
rect 4346 53254 4358 53306
rect 4410 53254 4422 53306
rect 4474 53254 4486 53306
rect 4538 53254 35014 53306
rect 35066 53254 35078 53306
rect 35130 53254 35142 53306
rect 35194 53254 35206 53306
rect 35258 53254 58848 53306
rect 1152 53232 58848 53254
rect 3280 52847 3286 52899
rect 3338 52887 3344 52899
rect 12403 52890 12461 52896
rect 12403 52887 12415 52890
rect 3338 52859 12415 52887
rect 3338 52847 3344 52859
rect 12403 52856 12415 52859
rect 12449 52887 12461 52890
rect 12595 52890 12653 52896
rect 12595 52887 12607 52890
rect 12449 52859 12607 52887
rect 12449 52856 12461 52859
rect 12403 52850 12461 52856
rect 12595 52856 12607 52859
rect 12641 52856 12653 52890
rect 12595 52850 12653 52856
rect 23539 52890 23597 52896
rect 23539 52856 23551 52890
rect 23585 52856 23597 52890
rect 23539 52850 23597 52856
rect 23554 52751 23582 52850
rect 25072 52847 25078 52899
rect 25130 52887 25136 52899
rect 40531 52890 40589 52896
rect 40531 52887 40543 52890
rect 25130 52859 40543 52887
rect 25130 52847 25136 52859
rect 40531 52856 40543 52859
rect 40577 52887 40589 52890
rect 40723 52890 40781 52896
rect 40723 52887 40735 52890
rect 40577 52859 40735 52887
rect 40577 52856 40589 52859
rect 40531 52850 40589 52856
rect 40723 52856 40735 52859
rect 40769 52856 40781 52890
rect 40723 52850 40781 52856
rect 23443 52742 23501 52748
rect 23443 52708 23455 52742
rect 23489 52739 23501 52742
rect 23536 52739 23542 52751
rect 23489 52711 23542 52739
rect 23489 52708 23501 52711
rect 23443 52702 23501 52708
rect 23536 52699 23542 52711
rect 23594 52699 23600 52751
rect 1152 52640 58848 52662
rect 1152 52588 19654 52640
rect 19706 52588 19718 52640
rect 19770 52588 19782 52640
rect 19834 52588 19846 52640
rect 19898 52588 50374 52640
rect 50426 52588 50438 52640
rect 50490 52588 50502 52640
rect 50554 52588 50566 52640
rect 50618 52588 58848 52640
rect 1152 52566 58848 52588
rect 11920 52181 11926 52233
rect 11978 52221 11984 52233
rect 32275 52224 32333 52230
rect 32275 52221 32287 52224
rect 11978 52193 32287 52221
rect 11978 52181 11984 52193
rect 32275 52190 32287 52193
rect 32321 52190 32333 52224
rect 32275 52184 32333 52190
rect 1152 51974 58848 51996
rect 1152 51922 4294 51974
rect 4346 51922 4358 51974
rect 4410 51922 4422 51974
rect 4474 51922 4486 51974
rect 4538 51922 35014 51974
rect 35066 51922 35078 51974
rect 35130 51922 35142 51974
rect 35194 51922 35206 51974
rect 35258 51922 58848 51974
rect 1152 51900 58848 51922
rect 23056 51515 23062 51567
rect 23114 51555 23120 51567
rect 41107 51558 41165 51564
rect 41107 51555 41119 51558
rect 23114 51527 41119 51555
rect 23114 51515 23120 51527
rect 41107 51524 41119 51527
rect 41153 51555 41165 51558
rect 41299 51558 41357 51564
rect 41299 51555 41311 51558
rect 41153 51527 41311 51555
rect 41153 51524 41165 51527
rect 41107 51518 41165 51524
rect 41299 51524 41311 51527
rect 41345 51524 41357 51558
rect 41299 51518 41357 51524
rect 1152 51308 58848 51330
rect 1152 51256 19654 51308
rect 19706 51256 19718 51308
rect 19770 51256 19782 51308
rect 19834 51256 19846 51308
rect 19898 51256 50374 51308
rect 50426 51256 50438 51308
rect 50490 51256 50502 51308
rect 50554 51256 50566 51308
rect 50618 51256 58848 51308
rect 1152 51234 58848 51256
rect 52723 51040 52781 51046
rect 52723 51006 52735 51040
rect 52769 51037 52781 51040
rect 57904 51037 57910 51049
rect 52769 51009 57910 51037
rect 52769 51006 52781 51009
rect 52723 51000 52781 51006
rect 57904 50997 57910 51009
rect 57962 50997 57968 51049
rect 1744 50849 1750 50901
rect 1802 50889 1808 50901
rect 51859 50892 51917 50898
rect 51859 50889 51871 50892
rect 1802 50861 51871 50889
rect 1802 50849 1808 50861
rect 51859 50858 51871 50861
rect 51905 50858 51917 50892
rect 51859 50852 51917 50858
rect 9424 50741 9430 50753
rect 9385 50713 9430 50741
rect 9424 50701 9430 50713
rect 9482 50741 9488 50753
rect 9811 50744 9869 50750
rect 9811 50741 9823 50744
rect 9482 50713 9823 50741
rect 9482 50701 9488 50713
rect 9811 50710 9823 50713
rect 9857 50710 9869 50744
rect 9811 50704 9869 50710
rect 10675 50744 10733 50750
rect 10675 50710 10687 50744
rect 10721 50741 10733 50744
rect 10963 50744 11021 50750
rect 10963 50741 10975 50744
rect 10721 50713 10975 50741
rect 10721 50710 10733 50713
rect 10675 50704 10733 50710
rect 10963 50710 10975 50713
rect 11009 50741 11021 50744
rect 50224 50741 50230 50753
rect 11009 50713 50230 50741
rect 11009 50710 11021 50713
rect 10963 50704 11021 50710
rect 50224 50701 50230 50713
rect 50282 50701 50288 50753
rect 1152 50642 58848 50664
rect 1152 50590 4294 50642
rect 4346 50590 4358 50642
rect 4410 50590 4422 50642
rect 4474 50590 4486 50642
rect 4538 50590 35014 50642
rect 35066 50590 35078 50642
rect 35130 50590 35142 50642
rect 35194 50590 35206 50642
rect 35258 50590 58848 50642
rect 1152 50568 58848 50590
rect 54832 50479 54838 50531
rect 54890 50519 54896 50531
rect 54931 50522 54989 50528
rect 54931 50519 54943 50522
rect 54890 50491 54943 50519
rect 54890 50479 54896 50491
rect 54931 50488 54943 50491
rect 54977 50488 54989 50522
rect 54931 50482 54989 50488
rect 10288 50445 10294 50457
rect 10249 50417 10294 50445
rect 10288 50405 10294 50417
rect 10346 50405 10352 50457
rect 10003 50374 10061 50380
rect 10003 50340 10015 50374
rect 10049 50371 10061 50374
rect 10306 50371 10334 50405
rect 10049 50343 10334 50371
rect 10049 50340 10061 50343
rect 10003 50334 10061 50340
rect 1152 49976 58848 49998
rect 1152 49924 19654 49976
rect 19706 49924 19718 49976
rect 19770 49924 19782 49976
rect 19834 49924 19846 49976
rect 19898 49924 50374 49976
rect 50426 49924 50438 49976
rect 50490 49924 50502 49976
rect 50554 49924 50566 49976
rect 50618 49924 58848 49976
rect 1152 49902 58848 49924
rect 10288 49665 10294 49717
rect 10346 49705 10352 49717
rect 29104 49705 29110 49717
rect 10346 49677 29110 49705
rect 10346 49665 10352 49677
rect 29104 49665 29110 49677
rect 29162 49665 29168 49717
rect 47536 49483 47542 49495
rect 27346 49455 47542 49483
rect 4243 49412 4301 49418
rect 4243 49378 4255 49412
rect 4289 49409 4301 49412
rect 4531 49412 4589 49418
rect 4531 49409 4543 49412
rect 4289 49381 4543 49409
rect 4289 49378 4301 49381
rect 4243 49372 4301 49378
rect 4531 49378 4543 49381
rect 4577 49409 4589 49412
rect 27346 49409 27374 49455
rect 47536 49443 47542 49455
rect 47594 49443 47600 49495
rect 33232 49409 33238 49421
rect 4577 49381 27374 49409
rect 33193 49381 33238 49409
rect 4577 49378 4589 49381
rect 4531 49372 4589 49378
rect 33232 49369 33238 49381
rect 33290 49409 33296 49421
rect 33427 49412 33485 49418
rect 33427 49409 33439 49412
rect 33290 49381 33439 49409
rect 33290 49369 33296 49381
rect 33427 49378 33439 49381
rect 33473 49378 33485 49412
rect 44176 49409 44182 49421
rect 44137 49381 44182 49409
rect 33427 49372 33485 49378
rect 44176 49369 44182 49381
rect 44234 49409 44240 49421
rect 44371 49412 44429 49418
rect 44371 49409 44383 49412
rect 44234 49381 44383 49409
rect 44234 49369 44240 49381
rect 44371 49378 44383 49381
rect 44417 49378 44429 49412
rect 44371 49372 44429 49378
rect 1152 49310 58848 49332
rect 1152 49258 4294 49310
rect 4346 49258 4358 49310
rect 4410 49258 4422 49310
rect 4474 49258 4486 49310
rect 4538 49258 35014 49310
rect 35066 49258 35078 49310
rect 35130 49258 35142 49310
rect 35194 49258 35206 49310
rect 35258 49258 58848 49310
rect 1152 49236 58848 49258
rect 9040 49147 9046 49199
rect 9098 49187 9104 49199
rect 44176 49187 44182 49199
rect 9098 49159 44182 49187
rect 9098 49147 9104 49159
rect 44176 49147 44182 49159
rect 44234 49147 44240 49199
rect 27280 49073 27286 49125
rect 27338 49113 27344 49125
rect 33232 49113 33238 49125
rect 27338 49085 33238 49113
rect 27338 49073 27344 49085
rect 33232 49073 33238 49085
rect 33290 49073 33296 49125
rect 27955 48894 28013 48900
rect 27955 48860 27967 48894
rect 28001 48891 28013 48894
rect 28243 48894 28301 48900
rect 28243 48891 28255 48894
rect 28001 48863 28255 48891
rect 28001 48860 28013 48863
rect 27955 48854 28013 48860
rect 28243 48860 28255 48863
rect 28289 48891 28301 48894
rect 39472 48891 39478 48903
rect 28289 48863 39478 48891
rect 28289 48860 28301 48863
rect 28243 48854 28301 48860
rect 39472 48851 39478 48863
rect 39530 48851 39536 48903
rect 1152 48644 58848 48666
rect 1152 48592 19654 48644
rect 19706 48592 19718 48644
rect 19770 48592 19782 48644
rect 19834 48592 19846 48644
rect 19898 48592 50374 48644
rect 50426 48592 50438 48644
rect 50490 48592 50502 48644
rect 50554 48592 50566 48644
rect 50618 48592 58848 48644
rect 1152 48570 58848 48592
rect 2419 48080 2477 48086
rect 2419 48046 2431 48080
rect 2465 48077 2477 48080
rect 2704 48077 2710 48089
rect 2465 48049 2710 48077
rect 2465 48046 2477 48049
rect 2419 48040 2477 48046
rect 2704 48037 2710 48049
rect 2762 48037 2768 48089
rect 37744 48037 37750 48089
rect 37802 48077 37808 48089
rect 41107 48080 41165 48086
rect 41107 48077 41119 48080
rect 37802 48049 41119 48077
rect 37802 48037 37808 48049
rect 41107 48046 41119 48049
rect 41153 48077 41165 48080
rect 41299 48080 41357 48086
rect 41299 48077 41311 48080
rect 41153 48049 41311 48077
rect 41153 48046 41165 48049
rect 41107 48040 41165 48046
rect 41299 48046 41311 48049
rect 41345 48046 41357 48080
rect 41299 48040 41357 48046
rect 1152 47978 58848 48000
rect 1152 47926 4294 47978
rect 4346 47926 4358 47978
rect 4410 47926 4422 47978
rect 4474 47926 4486 47978
rect 4538 47926 35014 47978
rect 35066 47926 35078 47978
rect 35130 47926 35142 47978
rect 35194 47926 35206 47978
rect 35258 47926 58848 47978
rect 1152 47904 58848 47926
rect 2704 47815 2710 47867
rect 2762 47855 2768 47867
rect 56944 47855 56950 47867
rect 2762 47827 56950 47855
rect 2762 47815 2768 47827
rect 56944 47815 56950 47827
rect 57002 47815 57008 47867
rect 8083 47562 8141 47568
rect 8083 47528 8095 47562
rect 8129 47559 8141 47562
rect 8371 47562 8429 47568
rect 8371 47559 8383 47562
rect 8129 47531 8383 47559
rect 8129 47528 8141 47531
rect 8083 47522 8141 47528
rect 8371 47528 8383 47531
rect 8417 47559 8429 47562
rect 28336 47559 28342 47571
rect 8417 47531 28342 47559
rect 8417 47528 8429 47531
rect 8371 47522 8429 47528
rect 28336 47519 28342 47531
rect 28394 47519 28400 47571
rect 49168 47485 49174 47497
rect 49129 47457 49174 47485
rect 49168 47445 49174 47457
rect 49226 47445 49232 47497
rect 1152 47312 58848 47334
rect 1152 47260 19654 47312
rect 19706 47260 19718 47312
rect 19770 47260 19782 47312
rect 19834 47260 19846 47312
rect 19898 47260 50374 47312
rect 50426 47260 50438 47312
rect 50490 47260 50502 47312
rect 50554 47260 50566 47312
rect 50618 47260 58848 47312
rect 1152 47238 58848 47260
rect 48208 47001 48214 47053
rect 48266 47041 48272 47053
rect 52723 47044 52781 47050
rect 52723 47041 52735 47044
rect 48266 47013 52735 47041
rect 48266 47001 48272 47013
rect 52723 47010 52735 47013
rect 52769 47010 52781 47044
rect 52723 47004 52781 47010
rect 36400 46745 36406 46757
rect 36361 46717 36406 46745
rect 36400 46705 36406 46717
rect 36458 46745 36464 46757
rect 36787 46748 36845 46754
rect 36787 46745 36799 46748
rect 36458 46717 36799 46745
rect 36458 46705 36464 46717
rect 36787 46714 36799 46717
rect 36833 46714 36845 46748
rect 36787 46708 36845 46714
rect 1152 46646 58848 46668
rect 1152 46594 4294 46646
rect 4346 46594 4358 46646
rect 4410 46594 4422 46646
rect 4474 46594 4486 46646
rect 4538 46594 35014 46646
rect 35066 46594 35078 46646
rect 35130 46594 35142 46646
rect 35194 46594 35206 46646
rect 35258 46594 58848 46646
rect 1152 46572 58848 46594
rect 17971 46230 18029 46236
rect 17971 46196 17983 46230
rect 18017 46196 18029 46230
rect 17971 46190 18029 46196
rect 17683 46156 17741 46162
rect 17683 46122 17695 46156
rect 17729 46153 17741 46156
rect 17986 46153 18014 46190
rect 54640 46153 54646 46165
rect 17729 46125 54646 46153
rect 17729 46122 17741 46125
rect 17683 46116 17741 46122
rect 54640 46113 54646 46125
rect 54698 46113 54704 46165
rect 1152 45980 58848 46002
rect 1152 45928 19654 45980
rect 19706 45928 19718 45980
rect 19770 45928 19782 45980
rect 19834 45928 19846 45980
rect 19898 45928 50374 45980
rect 50426 45928 50438 45980
rect 50490 45928 50502 45980
rect 50554 45928 50566 45980
rect 50618 45928 58848 45980
rect 1152 45906 58848 45928
rect 7696 45447 7702 45499
rect 7754 45487 7760 45499
rect 7754 45459 17294 45487
rect 7754 45447 7760 45459
rect 12499 45416 12557 45422
rect 12499 45382 12511 45416
rect 12545 45413 12557 45416
rect 12592 45413 12598 45425
rect 12545 45385 12598 45413
rect 12545 45382 12557 45385
rect 12499 45376 12557 45382
rect 12592 45373 12598 45385
rect 12650 45373 12656 45425
rect 17266 45413 17294 45459
rect 48019 45416 48077 45422
rect 48019 45413 48031 45416
rect 17266 45385 48031 45413
rect 48019 45382 48031 45385
rect 48065 45382 48077 45416
rect 48784 45413 48790 45425
rect 48745 45385 48790 45413
rect 48019 45376 48077 45382
rect 48784 45373 48790 45385
rect 48842 45413 48848 45425
rect 48979 45416 49037 45422
rect 48979 45413 48991 45416
rect 48842 45385 48991 45413
rect 48842 45373 48848 45385
rect 48979 45382 48991 45385
rect 49025 45382 49037 45416
rect 48979 45376 49037 45382
rect 55600 45373 55606 45425
rect 55658 45413 55664 45425
rect 55795 45416 55853 45422
rect 55795 45413 55807 45416
rect 55658 45385 55807 45413
rect 55658 45373 55664 45385
rect 55795 45382 55807 45385
rect 55841 45413 55853 45416
rect 55987 45416 56045 45422
rect 55987 45413 55999 45416
rect 55841 45385 55999 45413
rect 55841 45382 55853 45385
rect 55795 45376 55853 45382
rect 55987 45382 55999 45385
rect 56033 45382 56045 45416
rect 55987 45376 56045 45382
rect 1152 45314 58848 45336
rect 1152 45262 4294 45314
rect 4346 45262 4358 45314
rect 4410 45262 4422 45314
rect 4474 45262 4486 45314
rect 4538 45262 35014 45314
rect 35066 45262 35078 45314
rect 35130 45262 35142 45314
rect 35194 45262 35206 45314
rect 35258 45262 58848 45314
rect 1152 45240 58848 45262
rect 31792 45151 31798 45203
rect 31850 45191 31856 45203
rect 48784 45191 48790 45203
rect 31850 45163 48790 45191
rect 31850 45151 31856 45163
rect 48784 45151 48790 45163
rect 48842 45151 48848 45203
rect 12115 44898 12173 44904
rect 12115 44864 12127 44898
rect 12161 44895 12173 44898
rect 12403 44898 12461 44904
rect 12403 44895 12415 44898
rect 12161 44867 12415 44895
rect 12161 44864 12173 44867
rect 12115 44858 12173 44864
rect 12403 44864 12415 44867
rect 12449 44895 12461 44898
rect 12449 44867 17294 44895
rect 12449 44864 12461 44867
rect 12403 44858 12461 44864
rect 17266 44747 17294 44867
rect 29008 44747 29014 44759
rect 17266 44719 29014 44747
rect 29008 44707 29014 44719
rect 29066 44707 29072 44759
rect 1152 44648 58848 44670
rect 1152 44596 19654 44648
rect 19706 44596 19718 44648
rect 19770 44596 19782 44648
rect 19834 44596 19846 44648
rect 19898 44596 50374 44648
rect 50426 44596 50438 44648
rect 50490 44596 50502 44648
rect 50554 44596 50566 44648
rect 50618 44596 58848 44648
rect 1152 44574 58848 44596
rect 4243 44084 4301 44090
rect 4243 44050 4255 44084
rect 4289 44081 4301 44084
rect 4531 44084 4589 44090
rect 4531 44081 4543 44084
rect 4289 44053 4543 44081
rect 4289 44050 4301 44053
rect 4243 44044 4301 44050
rect 4531 44050 4543 44053
rect 4577 44081 4589 44084
rect 41104 44081 41110 44093
rect 4577 44053 41110 44081
rect 4577 44050 4589 44053
rect 4531 44044 4589 44050
rect 41104 44041 41110 44053
rect 41162 44041 41168 44093
rect 42256 44041 42262 44093
rect 42314 44081 42320 44093
rect 46387 44084 46445 44090
rect 46387 44081 46399 44084
rect 42314 44053 46399 44081
rect 42314 44041 42320 44053
rect 46387 44050 46399 44053
rect 46433 44081 46445 44084
rect 46579 44084 46637 44090
rect 46579 44081 46591 44084
rect 46433 44053 46591 44081
rect 46433 44050 46445 44053
rect 46387 44044 46445 44050
rect 46579 44050 46591 44053
rect 46625 44050 46637 44084
rect 46579 44044 46637 44050
rect 52051 44084 52109 44090
rect 52051 44050 52063 44084
rect 52097 44081 52109 44084
rect 52144 44081 52150 44093
rect 52097 44053 52150 44081
rect 52097 44050 52109 44053
rect 52051 44044 52109 44050
rect 52144 44041 52150 44053
rect 52202 44041 52208 44093
rect 1152 43982 58848 44004
rect 1152 43930 4294 43982
rect 4346 43930 4358 43982
rect 4410 43930 4422 43982
rect 4474 43930 4486 43982
rect 4538 43930 35014 43982
rect 35066 43930 35078 43982
rect 35130 43930 35142 43982
rect 35194 43930 35206 43982
rect 35258 43930 58848 43982
rect 1152 43908 58848 43930
rect 46291 43788 46349 43794
rect 46291 43754 46303 43788
rect 46337 43785 46349 43788
rect 46579 43788 46637 43794
rect 46579 43785 46591 43788
rect 46337 43757 46591 43785
rect 46337 43754 46349 43757
rect 46291 43748 46349 43754
rect 46579 43754 46591 43757
rect 46625 43785 46637 43788
rect 49552 43785 49558 43797
rect 46625 43757 49558 43785
rect 46625 43754 46637 43757
rect 46579 43748 46637 43754
rect 49552 43745 49558 43757
rect 49610 43745 49616 43797
rect 34576 43671 34582 43723
rect 34634 43711 34640 43723
rect 47539 43714 47597 43720
rect 47539 43711 47551 43714
rect 34634 43683 47551 43711
rect 34634 43671 34640 43683
rect 47539 43680 47551 43683
rect 47585 43680 47597 43714
rect 47539 43674 47597 43680
rect 56080 43637 56086 43649
rect 42082 43609 56086 43637
rect 17395 43566 17453 43572
rect 17395 43532 17407 43566
rect 17441 43563 17453 43566
rect 17683 43566 17741 43572
rect 17683 43563 17695 43566
rect 17441 43535 17695 43563
rect 17441 43532 17453 43535
rect 17395 43526 17453 43532
rect 17683 43532 17695 43535
rect 17729 43563 17741 43566
rect 42082 43563 42110 43609
rect 56080 43597 56086 43609
rect 56138 43597 56144 43649
rect 17729 43535 42110 43563
rect 47539 43566 47597 43572
rect 17729 43532 17741 43535
rect 17683 43526 17741 43532
rect 47539 43532 47551 43566
rect 47585 43563 47597 43566
rect 47731 43566 47789 43572
rect 47731 43563 47743 43566
rect 47585 43535 47743 43563
rect 47585 43532 47597 43535
rect 47539 43526 47597 43532
rect 47731 43532 47743 43535
rect 47777 43563 47789 43566
rect 47827 43566 47885 43572
rect 47827 43563 47839 43566
rect 47777 43535 47839 43563
rect 47777 43532 47789 43535
rect 47731 43526 47789 43532
rect 47827 43532 47839 43535
rect 47873 43532 47885 43566
rect 47827 43526 47885 43532
rect 51283 43566 51341 43572
rect 51283 43532 51295 43566
rect 51329 43532 51341 43566
rect 51283 43526 51341 43532
rect 23920 43449 23926 43501
rect 23978 43489 23984 43501
rect 51091 43492 51149 43498
rect 51091 43489 51103 43492
rect 23978 43461 51103 43489
rect 23978 43449 23984 43461
rect 51091 43458 51103 43461
rect 51137 43489 51149 43492
rect 51298 43489 51326 43526
rect 51137 43461 51326 43489
rect 51137 43458 51149 43461
rect 51091 43452 51149 43458
rect 1152 43316 58848 43338
rect 1152 43264 19654 43316
rect 19706 43264 19718 43316
rect 19770 43264 19782 43316
rect 19834 43264 19846 43316
rect 19898 43264 50374 43316
rect 50426 43264 50438 43316
rect 50490 43264 50502 43316
rect 50554 43264 50566 43316
rect 50618 43264 58848 43316
rect 1152 43242 58848 43264
rect 16147 42752 16205 42758
rect 16147 42718 16159 42752
rect 16193 42749 16205 42752
rect 16432 42749 16438 42761
rect 16193 42721 16438 42749
rect 16193 42718 16205 42721
rect 16147 42712 16205 42718
rect 16432 42709 16438 42721
rect 16490 42709 16496 42761
rect 20080 42749 20086 42761
rect 20041 42721 20086 42749
rect 20080 42709 20086 42721
rect 20138 42749 20144 42761
rect 20179 42752 20237 42758
rect 20179 42749 20191 42752
rect 20138 42721 20191 42749
rect 20138 42709 20144 42721
rect 20179 42718 20191 42721
rect 20225 42718 20237 42752
rect 20179 42712 20237 42718
rect 21136 42709 21142 42761
rect 21194 42749 21200 42761
rect 22675 42752 22733 42758
rect 22675 42749 22687 42752
rect 21194 42721 22687 42749
rect 21194 42709 21200 42721
rect 22675 42718 22687 42721
rect 22721 42749 22733 42752
rect 22867 42752 22925 42758
rect 22867 42749 22879 42752
rect 22721 42721 22879 42749
rect 22721 42718 22733 42721
rect 22675 42712 22733 42718
rect 22867 42718 22879 42721
rect 22913 42718 22925 42752
rect 52528 42749 52534 42761
rect 52489 42721 52534 42749
rect 22867 42712 22925 42718
rect 52528 42709 52534 42721
rect 52586 42749 52592 42761
rect 52723 42752 52781 42758
rect 52723 42749 52735 42752
rect 52586 42721 52735 42749
rect 52586 42709 52592 42721
rect 52723 42718 52735 42721
rect 52769 42718 52781 42752
rect 52723 42712 52781 42718
rect 1152 42650 58848 42672
rect 1152 42598 4294 42650
rect 4346 42598 4358 42650
rect 4410 42598 4422 42650
rect 4474 42598 4486 42650
rect 4538 42598 35014 42650
rect 35066 42598 35078 42650
rect 35130 42598 35142 42650
rect 35194 42598 35206 42650
rect 35258 42598 58848 42650
rect 1152 42576 58848 42598
rect 16432 42487 16438 42539
rect 16490 42527 16496 42539
rect 27760 42527 27766 42539
rect 16490 42499 27766 42527
rect 16490 42487 16496 42499
rect 27760 42487 27766 42499
rect 27818 42487 27824 42539
rect 3571 42234 3629 42240
rect 3571 42200 3583 42234
rect 3617 42231 3629 42234
rect 16720 42231 16726 42243
rect 3617 42203 16726 42231
rect 3617 42200 3629 42203
rect 3571 42194 3629 42200
rect 16720 42191 16726 42203
rect 16778 42191 16784 42243
rect 29971 42234 30029 42240
rect 29971 42231 29983 42234
rect 29794 42203 29983 42231
rect 3664 42043 3670 42095
rect 3722 42083 3728 42095
rect 29794 42092 29822 42203
rect 29971 42200 29983 42203
rect 30017 42200 30029 42234
rect 29971 42194 30029 42200
rect 45331 42234 45389 42240
rect 45331 42200 45343 42234
rect 45377 42200 45389 42234
rect 45331 42194 45389 42200
rect 45346 42095 45374 42194
rect 29779 42086 29837 42092
rect 29779 42083 29791 42086
rect 3722 42055 29791 42083
rect 3722 42043 3728 42055
rect 29779 42052 29791 42055
rect 29825 42052 29837 42086
rect 29779 42046 29837 42052
rect 45235 42086 45293 42092
rect 45235 42052 45247 42086
rect 45281 42083 45293 42086
rect 45328 42083 45334 42095
rect 45281 42055 45334 42083
rect 45281 42052 45293 42055
rect 45235 42046 45293 42052
rect 45328 42043 45334 42055
rect 45386 42043 45392 42095
rect 1152 41984 58848 42006
rect 1152 41932 19654 41984
rect 19706 41932 19718 41984
rect 19770 41932 19782 41984
rect 19834 41932 19846 41984
rect 19898 41932 50374 41984
rect 50426 41932 50438 41984
rect 50490 41932 50502 41984
rect 50554 41932 50566 41984
rect 50618 41932 58848 41984
rect 1152 41910 58848 41932
rect 1152 41318 58848 41340
rect 1152 41266 4294 41318
rect 4346 41266 4358 41318
rect 4410 41266 4422 41318
rect 4474 41266 4486 41318
rect 4538 41266 35014 41318
rect 35066 41266 35078 41318
rect 35130 41266 35142 41318
rect 35194 41266 35206 41318
rect 35258 41266 58848 41318
rect 1152 41244 58848 41266
rect 33328 40859 33334 40911
rect 33386 40899 33392 40911
rect 33811 40902 33869 40908
rect 33811 40899 33823 40902
rect 33386 40871 33823 40899
rect 33386 40859 33392 40871
rect 33811 40868 33823 40871
rect 33857 40868 33869 40902
rect 49747 40902 49805 40908
rect 49747 40899 49759 40902
rect 33811 40862 33869 40868
rect 37426 40871 49759 40899
rect 18832 40785 18838 40837
rect 18890 40825 18896 40837
rect 37426 40825 37454 40871
rect 49747 40868 49759 40871
rect 49793 40899 49805 40902
rect 49939 40902 49997 40908
rect 49939 40899 49951 40902
rect 49793 40871 49951 40899
rect 49793 40868 49805 40871
rect 49747 40862 49805 40868
rect 49939 40868 49951 40871
rect 49985 40868 49997 40902
rect 49939 40862 49997 40868
rect 18890 40797 37454 40825
rect 47506 40797 57614 40825
rect 18890 40785 18896 40797
rect 33328 40711 33334 40763
rect 33386 40751 33392 40763
rect 33619 40754 33677 40760
rect 33619 40751 33631 40754
rect 33386 40723 33631 40751
rect 33386 40711 33392 40723
rect 33619 40720 33631 40723
rect 33665 40720 33677 40754
rect 33619 40714 33677 40720
rect 40240 40711 40246 40763
rect 40298 40751 40304 40763
rect 47506 40751 47534 40797
rect 40298 40723 47534 40751
rect 57586 40751 57614 40797
rect 57715 40754 57773 40760
rect 57715 40751 57727 40754
rect 57586 40723 57727 40751
rect 40298 40711 40304 40723
rect 57715 40720 57727 40723
rect 57761 40720 57773 40754
rect 57715 40714 57773 40720
rect 1152 40652 58848 40674
rect 1152 40600 19654 40652
rect 19706 40600 19718 40652
rect 19770 40600 19782 40652
rect 19834 40600 19846 40652
rect 19898 40600 50374 40652
rect 50426 40600 50438 40652
rect 50490 40600 50502 40652
rect 50554 40600 50566 40652
rect 50618 40600 58848 40652
rect 1152 40578 58848 40600
rect 15184 40489 15190 40541
rect 15242 40529 15248 40541
rect 16531 40532 16589 40538
rect 16531 40529 16543 40532
rect 15242 40501 16543 40529
rect 15242 40489 15248 40501
rect 16531 40498 16543 40501
rect 16577 40498 16589 40532
rect 16531 40492 16589 40498
rect 15952 40045 15958 40097
rect 16010 40085 16016 40097
rect 17011 40088 17069 40094
rect 17011 40085 17023 40088
rect 16010 40057 17023 40085
rect 16010 40045 16016 40057
rect 17011 40054 17023 40057
rect 17057 40085 17069 40088
rect 17203 40088 17261 40094
rect 17203 40085 17215 40088
rect 17057 40057 17215 40085
rect 17057 40054 17069 40057
rect 17011 40048 17069 40054
rect 17203 40054 17215 40057
rect 17249 40054 17261 40088
rect 23344 40085 23350 40097
rect 23305 40057 23350 40085
rect 17203 40048 17261 40054
rect 23344 40045 23350 40057
rect 23402 40085 23408 40097
rect 23539 40088 23597 40094
rect 23539 40085 23551 40088
rect 23402 40057 23551 40085
rect 23402 40045 23408 40057
rect 23539 40054 23551 40057
rect 23585 40054 23597 40088
rect 47248 40085 47254 40097
rect 47209 40057 47254 40085
rect 23539 40048 23597 40054
rect 47248 40045 47254 40057
rect 47306 40085 47312 40097
rect 47443 40088 47501 40094
rect 47443 40085 47455 40088
rect 47306 40057 47455 40085
rect 47306 40045 47312 40057
rect 47443 40054 47455 40057
rect 47489 40054 47501 40088
rect 47443 40048 47501 40054
rect 1152 39986 58848 40008
rect 1152 39934 4294 39986
rect 4346 39934 4358 39986
rect 4410 39934 4422 39986
rect 4474 39934 4486 39986
rect 4538 39934 35014 39986
rect 35066 39934 35078 39986
rect 35130 39934 35142 39986
rect 35194 39934 35206 39986
rect 35258 39934 58848 39986
rect 1152 39912 58848 39934
rect 15856 39823 15862 39875
rect 15914 39863 15920 39875
rect 47248 39863 47254 39875
rect 15914 39835 47254 39863
rect 15914 39823 15920 39835
rect 47248 39823 47254 39835
rect 47306 39823 47312 39875
rect 47923 39570 47981 39576
rect 47923 39536 47935 39570
rect 47969 39567 47981 39570
rect 48211 39570 48269 39576
rect 48211 39567 48223 39570
rect 47969 39539 48223 39567
rect 47969 39536 47981 39539
rect 47923 39530 47981 39536
rect 48211 39536 48223 39539
rect 48257 39567 48269 39570
rect 49456 39567 49462 39579
rect 48257 39539 49462 39567
rect 48257 39536 48269 39539
rect 48211 39530 48269 39536
rect 49456 39527 49462 39539
rect 49514 39527 49520 39579
rect 51283 39570 51341 39576
rect 51283 39536 51295 39570
rect 51329 39567 51341 39570
rect 51571 39570 51629 39576
rect 51571 39567 51583 39570
rect 51329 39539 51583 39567
rect 51329 39536 51341 39539
rect 51283 39530 51341 39536
rect 51571 39536 51583 39539
rect 51617 39567 51629 39570
rect 52912 39567 52918 39579
rect 51617 39539 52918 39567
rect 51617 39536 51629 39539
rect 51571 39530 51629 39536
rect 52912 39527 52918 39539
rect 52970 39527 52976 39579
rect 1152 39320 58848 39342
rect 1152 39268 19654 39320
rect 19706 39268 19718 39320
rect 19770 39268 19782 39320
rect 19834 39268 19846 39320
rect 19898 39268 50374 39320
rect 50426 39268 50438 39320
rect 50490 39268 50502 39320
rect 50554 39268 50566 39320
rect 50618 39268 58848 39320
rect 1152 39246 58848 39268
rect 34291 38904 34349 38910
rect 34291 38870 34303 38904
rect 34337 38901 34349 38904
rect 34337 38873 34622 38901
rect 34337 38870 34349 38873
rect 34291 38864 34349 38870
rect 22960 38713 22966 38765
rect 23018 38753 23024 38765
rect 34594 38762 34622 38873
rect 32083 38756 32141 38762
rect 32083 38753 32095 38756
rect 23018 38725 32095 38753
rect 23018 38713 23024 38725
rect 32083 38722 32095 38725
rect 32129 38722 32141 38756
rect 32083 38716 32141 38722
rect 34579 38756 34637 38762
rect 34579 38722 34591 38756
rect 34625 38753 34637 38756
rect 38704 38753 38710 38765
rect 34625 38725 38710 38753
rect 34625 38722 34637 38725
rect 34579 38716 34637 38722
rect 38704 38713 38710 38725
rect 38762 38713 38768 38765
rect 1152 38654 58848 38676
rect 1152 38602 4294 38654
rect 4346 38602 4358 38654
rect 4410 38602 4422 38654
rect 4474 38602 4486 38654
rect 4538 38602 35014 38654
rect 35066 38602 35078 38654
rect 35130 38602 35142 38654
rect 35194 38602 35206 38654
rect 35258 38602 58848 38654
rect 1152 38580 58848 38602
rect 6352 38195 6358 38247
rect 6410 38235 6416 38247
rect 17683 38238 17741 38244
rect 17683 38235 17695 38238
rect 6410 38207 17695 38235
rect 6410 38195 6416 38207
rect 17683 38204 17695 38207
rect 17729 38204 17741 38238
rect 17683 38198 17741 38204
rect 20464 38195 20470 38247
rect 20522 38235 20528 38247
rect 36883 38238 36941 38244
rect 36883 38235 36895 38238
rect 20522 38207 36895 38235
rect 20522 38195 20528 38207
rect 36883 38204 36895 38207
rect 36929 38204 36941 38238
rect 36883 38198 36941 38204
rect 1152 37988 58848 38010
rect 1152 37936 19654 37988
rect 19706 37936 19718 37988
rect 19770 37936 19782 37988
rect 19834 37936 19846 37988
rect 19898 37936 50374 37988
rect 50426 37936 50438 37988
rect 50490 37936 50502 37988
rect 50554 37936 50566 37988
rect 50618 37936 58848 37988
rect 1152 37914 58848 37936
rect 51184 37455 51190 37507
rect 51242 37495 51248 37507
rect 51667 37498 51725 37504
rect 51667 37495 51679 37498
rect 51242 37467 51679 37495
rect 51242 37455 51248 37467
rect 51667 37464 51679 37467
rect 51713 37464 51725 37498
rect 51667 37458 51725 37464
rect 1843 37424 1901 37430
rect 1843 37390 1855 37424
rect 1889 37421 1901 37424
rect 2035 37424 2093 37430
rect 2035 37421 2047 37424
rect 1889 37393 2047 37421
rect 1889 37390 1901 37393
rect 1843 37384 1901 37390
rect 2035 37390 2047 37393
rect 2081 37421 2093 37424
rect 2416 37421 2422 37433
rect 2081 37393 2422 37421
rect 2081 37390 2093 37393
rect 2035 37384 2093 37390
rect 2416 37381 2422 37393
rect 2474 37381 2480 37433
rect 5491 37424 5549 37430
rect 5491 37390 5503 37424
rect 5537 37421 5549 37424
rect 6448 37421 6454 37433
rect 5537 37393 6454 37421
rect 5537 37390 5549 37393
rect 5491 37384 5549 37390
rect 6448 37381 6454 37393
rect 6506 37381 6512 37433
rect 47344 37381 47350 37433
rect 47402 37421 47408 37433
rect 47443 37424 47501 37430
rect 47443 37421 47455 37424
rect 47402 37393 47455 37421
rect 47402 37381 47408 37393
rect 47443 37390 47455 37393
rect 47489 37390 47501 37424
rect 51682 37421 51710 37458
rect 51859 37424 51917 37430
rect 51859 37421 51871 37424
rect 51682 37393 51871 37421
rect 47443 37384 47501 37390
rect 51859 37390 51871 37393
rect 51905 37390 51917 37424
rect 51859 37384 51917 37390
rect 1152 37322 58848 37344
rect 1152 37270 4294 37322
rect 4346 37270 4358 37322
rect 4410 37270 4422 37322
rect 4474 37270 4486 37322
rect 4538 37270 35014 37322
rect 35066 37270 35078 37322
rect 35130 37270 35142 37322
rect 35194 37270 35206 37322
rect 35258 37270 58848 37322
rect 1152 37248 58848 37270
rect 24979 37128 25037 37134
rect 24979 37094 24991 37128
rect 25025 37125 25037 37128
rect 25025 37097 37454 37125
rect 25025 37094 25037 37097
rect 24979 37088 25037 37094
rect 2512 37011 2518 37063
rect 2570 37051 2576 37063
rect 6931 37054 6989 37060
rect 6931 37051 6943 37054
rect 2570 37023 6943 37051
rect 2570 37011 2576 37023
rect 6931 37020 6943 37023
rect 6977 37020 6989 37054
rect 6931 37014 6989 37020
rect 23728 37011 23734 37063
rect 23786 37051 23792 37063
rect 23786 37023 31070 37051
rect 23786 37011 23792 37023
rect 27955 36906 28013 36912
rect 27955 36872 27967 36906
rect 28001 36903 28013 36906
rect 28240 36903 28246 36915
rect 28001 36875 28246 36903
rect 28001 36872 28013 36875
rect 27955 36866 28013 36872
rect 28240 36863 28246 36875
rect 28298 36863 28304 36915
rect 31042 36903 31070 37023
rect 37426 36977 37454 37097
rect 51568 36977 51574 36989
rect 37426 36949 51574 36977
rect 51568 36937 51574 36949
rect 51626 36937 51632 36989
rect 56371 36906 56429 36912
rect 56371 36903 56383 36906
rect 31042 36875 56383 36903
rect 56371 36872 56383 36875
rect 56417 36872 56429 36906
rect 56371 36866 56429 36872
rect 24115 36832 24173 36838
rect 24115 36798 24127 36832
rect 24161 36829 24173 36832
rect 24161 36801 37454 36829
rect 24161 36798 24173 36801
rect 24115 36792 24173 36798
rect 37426 36755 37454 36801
rect 49840 36755 49846 36767
rect 37426 36727 49846 36755
rect 49840 36715 49846 36727
rect 49898 36715 49904 36767
rect 1152 36656 58848 36678
rect 1152 36604 19654 36656
rect 19706 36604 19718 36656
rect 19770 36604 19782 36656
rect 19834 36604 19846 36656
rect 19898 36604 50374 36656
rect 50426 36604 50438 36656
rect 50490 36604 50502 36656
rect 50554 36604 50566 36656
rect 50618 36604 58848 36656
rect 1152 36582 58848 36604
rect 28240 36493 28246 36545
rect 28298 36533 28304 36545
rect 45424 36533 45430 36545
rect 28298 36505 45430 36533
rect 28298 36493 28304 36505
rect 45424 36493 45430 36505
rect 45482 36493 45488 36545
rect 13936 36271 13942 36323
rect 13994 36311 14000 36323
rect 33427 36314 33485 36320
rect 33427 36311 33439 36314
rect 13994 36283 33439 36311
rect 13994 36271 14000 36283
rect 33427 36280 33439 36283
rect 33473 36311 33485 36314
rect 33619 36314 33677 36320
rect 33619 36311 33631 36314
rect 33473 36283 33631 36311
rect 33473 36280 33485 36283
rect 33427 36274 33485 36280
rect 33619 36280 33631 36283
rect 33665 36280 33677 36314
rect 37168 36311 37174 36323
rect 33619 36274 33677 36280
rect 33730 36283 37174 36311
rect 5584 36197 5590 36249
rect 5642 36237 5648 36249
rect 22003 36240 22061 36246
rect 22003 36237 22015 36240
rect 5642 36209 22015 36237
rect 5642 36197 5648 36209
rect 22003 36206 22015 36209
rect 22049 36206 22061 36240
rect 22003 36200 22061 36206
rect 31024 36197 31030 36249
rect 31082 36237 31088 36249
rect 33730 36237 33758 36283
rect 37168 36271 37174 36283
rect 37226 36271 37232 36323
rect 31082 36209 33758 36237
rect 37075 36240 37133 36246
rect 31082 36197 31088 36209
rect 37075 36206 37087 36240
rect 37121 36237 37133 36240
rect 51280 36237 51286 36249
rect 37121 36209 51286 36237
rect 37121 36206 37133 36209
rect 37075 36200 37133 36206
rect 51280 36197 51286 36209
rect 51338 36197 51344 36249
rect 25555 36166 25613 36172
rect 25555 36132 25567 36166
rect 25601 36163 25613 36166
rect 25843 36166 25901 36172
rect 25843 36163 25855 36166
rect 25601 36135 25855 36163
rect 25601 36132 25613 36135
rect 25555 36126 25613 36132
rect 25843 36132 25855 36135
rect 25889 36163 25901 36166
rect 43888 36163 43894 36175
rect 25889 36135 43894 36163
rect 25889 36132 25901 36135
rect 25843 36126 25901 36132
rect 43888 36123 43894 36135
rect 43946 36123 43952 36175
rect 21235 36092 21293 36098
rect 21235 36058 21247 36092
rect 21281 36089 21293 36092
rect 21523 36092 21581 36098
rect 21523 36089 21535 36092
rect 21281 36061 21535 36089
rect 21281 36058 21293 36061
rect 21235 36052 21293 36058
rect 21523 36058 21535 36061
rect 21569 36089 21581 36092
rect 24112 36089 24118 36101
rect 21569 36061 24118 36089
rect 21569 36058 21581 36061
rect 21523 36052 21581 36058
rect 24112 36049 24118 36061
rect 24170 36049 24176 36101
rect 36691 36092 36749 36098
rect 36691 36058 36703 36092
rect 36737 36089 36749 36092
rect 36979 36092 37037 36098
rect 36979 36089 36991 36092
rect 36737 36061 36991 36089
rect 36737 36058 36749 36061
rect 36691 36052 36749 36058
rect 36979 36058 36991 36061
rect 37025 36089 37037 36092
rect 37075 36092 37133 36098
rect 37075 36089 37087 36092
rect 37025 36061 37087 36089
rect 37025 36058 37037 36061
rect 36979 36052 37037 36058
rect 37075 36058 37087 36061
rect 37121 36058 37133 36092
rect 37075 36052 37133 36058
rect 37168 36049 37174 36101
rect 37226 36089 37232 36101
rect 50611 36092 50669 36098
rect 50611 36089 50623 36092
rect 37226 36061 50623 36089
rect 37226 36049 37232 36061
rect 50611 36058 50623 36061
rect 50657 36058 50669 36092
rect 50611 36052 50669 36058
rect 1152 35990 58848 36012
rect 1152 35938 4294 35990
rect 4346 35938 4358 35990
rect 4410 35938 4422 35990
rect 4474 35938 4486 35990
rect 4538 35938 35014 35990
rect 35066 35938 35078 35990
rect 35130 35938 35142 35990
rect 35194 35938 35206 35990
rect 35258 35938 58848 35990
rect 1152 35916 58848 35938
rect 41491 35722 41549 35728
rect 41491 35688 41503 35722
rect 41537 35719 41549 35722
rect 49936 35719 49942 35731
rect 41537 35691 49942 35719
rect 41537 35688 41549 35691
rect 41491 35682 41549 35688
rect 49936 35679 49942 35691
rect 49994 35679 50000 35731
rect 46387 35574 46445 35580
rect 46387 35540 46399 35574
rect 46433 35571 46445 35574
rect 46675 35574 46733 35580
rect 46675 35571 46687 35574
rect 46433 35543 46687 35571
rect 46433 35540 46445 35543
rect 46387 35534 46445 35540
rect 46675 35540 46687 35543
rect 46721 35571 46733 35574
rect 48592 35571 48598 35583
rect 46721 35543 48598 35571
rect 46721 35540 46733 35543
rect 46675 35534 46733 35540
rect 48592 35531 48598 35543
rect 48650 35531 48656 35583
rect 1152 35324 58848 35346
rect 1152 35272 19654 35324
rect 19706 35272 19718 35324
rect 19770 35272 19782 35324
rect 19834 35272 19846 35324
rect 19898 35272 50374 35324
rect 50426 35272 50438 35324
rect 50490 35272 50502 35324
rect 50554 35272 50566 35324
rect 50618 35272 58848 35324
rect 1152 35250 58848 35272
rect 12595 34834 12653 34840
rect 12595 34800 12607 34834
rect 12641 34831 12653 34834
rect 12883 34834 12941 34840
rect 12883 34831 12895 34834
rect 12641 34803 12895 34831
rect 12641 34800 12653 34803
rect 12595 34794 12653 34800
rect 12883 34800 12895 34803
rect 12929 34831 12941 34834
rect 33712 34831 33718 34843
rect 12929 34803 33718 34831
rect 12929 34800 12941 34803
rect 12883 34794 12941 34800
rect 33712 34791 33718 34803
rect 33770 34791 33776 34843
rect 11344 34717 11350 34769
rect 11402 34757 11408 34769
rect 41491 34760 41549 34766
rect 41491 34757 41503 34760
rect 11402 34729 41503 34757
rect 11402 34717 11408 34729
rect 41491 34726 41503 34729
rect 41537 34757 41549 34760
rect 41683 34760 41741 34766
rect 41683 34757 41695 34760
rect 41537 34729 41695 34757
rect 41537 34726 41549 34729
rect 41491 34720 41549 34726
rect 41683 34726 41695 34729
rect 41729 34726 41741 34760
rect 41683 34720 41741 34726
rect 1152 34658 58848 34680
rect 1152 34606 4294 34658
rect 4346 34606 4358 34658
rect 4410 34606 4422 34658
rect 4474 34606 4486 34658
rect 4538 34606 35014 34658
rect 35066 34606 35078 34658
rect 35130 34606 35142 34658
rect 35194 34606 35206 34658
rect 35258 34606 58848 34658
rect 1152 34584 58848 34606
rect 17875 34390 17933 34396
rect 17875 34356 17887 34390
rect 17921 34387 17933 34390
rect 26992 34387 26998 34399
rect 17921 34359 26998 34387
rect 17921 34356 17933 34359
rect 17875 34350 17933 34356
rect 26992 34347 26998 34359
rect 27050 34347 27056 34399
rect 13843 34316 13901 34322
rect 13843 34282 13855 34316
rect 13889 34313 13901 34316
rect 14131 34316 14189 34322
rect 14131 34313 14143 34316
rect 13889 34285 14143 34313
rect 13889 34282 13901 34285
rect 13843 34276 13901 34282
rect 14131 34282 14143 34285
rect 14177 34313 14189 34316
rect 14177 34285 27374 34313
rect 14177 34282 14189 34285
rect 14131 34276 14189 34282
rect 9904 34239 9910 34251
rect 9865 34211 9910 34239
rect 9904 34199 9910 34211
rect 9962 34199 9968 34251
rect 21427 34242 21485 34248
rect 21427 34208 21439 34242
rect 21473 34208 21485 34242
rect 27346 34239 27374 34285
rect 49936 34239 49942 34251
rect 27346 34211 49942 34239
rect 21427 34202 21485 34208
rect 21139 34168 21197 34174
rect 21139 34134 21151 34168
rect 21185 34165 21197 34168
rect 21442 34165 21470 34202
rect 49936 34199 49942 34211
rect 49994 34199 50000 34251
rect 21185 34137 27374 34165
rect 21185 34134 21197 34137
rect 21139 34128 21197 34134
rect 27346 34091 27374 34137
rect 48784 34091 48790 34103
rect 27346 34063 48790 34091
rect 48784 34051 48790 34063
rect 48842 34051 48848 34103
rect 1152 33992 58848 34014
rect 1152 33940 19654 33992
rect 19706 33940 19718 33992
rect 19770 33940 19782 33992
rect 19834 33940 19846 33992
rect 19898 33940 50374 33992
rect 50426 33940 50438 33992
rect 50490 33940 50502 33992
rect 50554 33940 50566 33992
rect 50618 33940 58848 33992
rect 1152 33918 58848 33940
rect 42064 33681 42070 33733
rect 42122 33721 42128 33733
rect 56179 33724 56237 33730
rect 56179 33721 56191 33724
rect 42122 33693 56191 33721
rect 42122 33681 42128 33693
rect 56179 33690 56191 33693
rect 56225 33690 56237 33724
rect 56179 33684 56237 33690
rect 31696 33607 31702 33659
rect 31754 33647 31760 33659
rect 42163 33650 42221 33656
rect 42163 33647 42175 33650
rect 31754 33619 42175 33647
rect 31754 33607 31760 33619
rect 42163 33616 42175 33619
rect 42209 33647 42221 33650
rect 42355 33650 42413 33656
rect 42355 33647 42367 33650
rect 42209 33619 42367 33647
rect 42209 33616 42221 33619
rect 42163 33610 42221 33616
rect 42355 33616 42367 33619
rect 42401 33616 42413 33650
rect 42355 33610 42413 33616
rect 34768 33533 34774 33585
rect 34826 33573 34832 33585
rect 44944 33573 44950 33585
rect 34826 33545 44950 33573
rect 34826 33533 34832 33545
rect 44944 33533 44950 33545
rect 45002 33533 45008 33585
rect 35344 33459 35350 33511
rect 35402 33499 35408 33511
rect 35402 33471 42494 33499
rect 35402 33459 35408 33471
rect 27856 33385 27862 33437
rect 27914 33425 27920 33437
rect 29299 33428 29357 33434
rect 29299 33425 29311 33428
rect 27914 33397 29311 33425
rect 27914 33385 27920 33397
rect 29299 33394 29311 33397
rect 29345 33425 29357 33428
rect 29491 33428 29549 33434
rect 29491 33425 29503 33428
rect 29345 33397 29503 33425
rect 29345 33394 29357 33397
rect 29299 33388 29357 33394
rect 29491 33394 29503 33397
rect 29537 33394 29549 33428
rect 34672 33425 34678 33437
rect 34633 33397 34678 33425
rect 29491 33388 29549 33394
rect 34672 33385 34678 33397
rect 34730 33385 34736 33437
rect 37939 33428 37997 33434
rect 37939 33394 37951 33428
rect 37985 33425 37997 33428
rect 38224 33425 38230 33437
rect 37985 33397 38230 33425
rect 37985 33394 37997 33397
rect 37939 33388 37997 33394
rect 38224 33385 38230 33397
rect 38282 33385 38288 33437
rect 42466 33425 42494 33471
rect 55507 33428 55565 33434
rect 55507 33425 55519 33428
rect 42466 33397 55519 33425
rect 55507 33394 55519 33397
rect 55553 33394 55565 33428
rect 55507 33388 55565 33394
rect 1152 33326 58848 33348
rect 1152 33274 4294 33326
rect 4346 33274 4358 33326
rect 4410 33274 4422 33326
rect 4474 33274 4486 33326
rect 4538 33274 35014 33326
rect 35066 33274 35078 33326
rect 35130 33274 35142 33326
rect 35194 33274 35206 33326
rect 35258 33274 58848 33326
rect 1152 33252 58848 33274
rect 37651 33206 37709 33212
rect 37651 33172 37663 33206
rect 37697 33203 37709 33206
rect 49648 33203 49654 33215
rect 37697 33175 49654 33203
rect 37697 33172 37709 33175
rect 37651 33166 37709 33172
rect 49648 33163 49654 33175
rect 49706 33163 49712 33215
rect 44944 33129 44950 33141
rect 44905 33101 44950 33129
rect 44944 33089 44950 33101
rect 45002 33089 45008 33141
rect 29395 32910 29453 32916
rect 29395 32907 29407 32910
rect 29218 32879 29407 32907
rect 22576 32719 22582 32771
rect 22634 32759 22640 32771
rect 29218 32768 29246 32879
rect 29395 32876 29407 32879
rect 29441 32876 29453 32910
rect 29395 32870 29453 32876
rect 29203 32762 29261 32768
rect 29203 32759 29215 32762
rect 22634 32731 29215 32759
rect 22634 32719 22640 32731
rect 29203 32728 29215 32731
rect 29249 32728 29261 32762
rect 29203 32722 29261 32728
rect 1152 32660 58848 32682
rect 1152 32608 19654 32660
rect 19706 32608 19718 32660
rect 19770 32608 19782 32660
rect 19834 32608 19846 32660
rect 19898 32608 50374 32660
rect 50426 32608 50438 32660
rect 50490 32608 50502 32660
rect 50554 32608 50566 32660
rect 50618 32608 58848 32660
rect 1152 32586 58848 32608
rect 2320 32093 2326 32105
rect 2281 32065 2326 32093
rect 2320 32053 2326 32065
rect 2378 32053 2384 32105
rect 6643 32096 6701 32102
rect 6643 32062 6655 32096
rect 6689 32093 6701 32096
rect 6736 32093 6742 32105
rect 6689 32065 6742 32093
rect 6689 32062 6701 32065
rect 6643 32056 6701 32062
rect 6736 32053 6742 32065
rect 6794 32053 6800 32105
rect 1152 31994 58848 32016
rect 1152 31942 4294 31994
rect 4346 31942 4358 31994
rect 4410 31942 4422 31994
rect 4474 31942 4486 31994
rect 4538 31942 35014 31994
rect 35066 31942 35078 31994
rect 35130 31942 35142 31994
rect 35194 31942 35206 31994
rect 35258 31942 58848 31994
rect 1152 31920 58848 31942
rect 1152 31328 58848 31350
rect 1152 31276 19654 31328
rect 19706 31276 19718 31328
rect 19770 31276 19782 31328
rect 19834 31276 19846 31328
rect 19898 31276 50374 31328
rect 50426 31276 50438 31328
rect 50490 31276 50502 31328
rect 50554 31276 50566 31328
rect 50618 31276 58848 31328
rect 1152 31254 58848 31276
rect 7312 30943 7318 30995
rect 7370 30983 7376 30995
rect 43408 30983 43414 30995
rect 7370 30955 43414 30983
rect 7370 30943 7376 30955
rect 43408 30943 43414 30955
rect 43466 30943 43472 30995
rect 41299 30912 41357 30918
rect 41299 30878 41311 30912
rect 41345 30909 41357 30912
rect 53008 30909 53014 30921
rect 41345 30881 53014 30909
rect 41345 30878 41357 30881
rect 41299 30872 41357 30878
rect 53008 30869 53014 30881
rect 53066 30869 53072 30921
rect 11731 30838 11789 30844
rect 11731 30804 11743 30838
rect 11777 30835 11789 30838
rect 11777 30807 37454 30835
rect 11777 30804 11789 30807
rect 11731 30798 11789 30804
rect 6640 30761 6646 30773
rect 6601 30733 6646 30761
rect 6640 30721 6646 30733
rect 6698 30721 6704 30773
rect 28147 30764 28205 30770
rect 28147 30730 28159 30764
rect 28193 30761 28205 30764
rect 34768 30761 34774 30773
rect 28193 30733 34774 30761
rect 28193 30730 28205 30733
rect 28147 30724 28205 30730
rect 34768 30721 34774 30733
rect 34826 30721 34832 30773
rect 37426 30761 37454 30807
rect 49840 30761 49846 30773
rect 37426 30733 49846 30761
rect 49840 30721 49846 30733
rect 49898 30721 49904 30773
rect 1152 30662 58848 30684
rect 1152 30610 4294 30662
rect 4346 30610 4358 30662
rect 4410 30610 4422 30662
rect 4474 30610 4486 30662
rect 4538 30610 35014 30662
rect 35066 30610 35078 30662
rect 35130 30610 35142 30662
rect 35194 30610 35206 30662
rect 35258 30610 58848 30662
rect 1152 30588 58848 30610
rect 28339 30394 28397 30400
rect 28339 30360 28351 30394
rect 28385 30391 28397 30394
rect 28385 30363 37454 30391
rect 28385 30360 28397 30363
rect 28339 30354 28397 30360
rect 7027 30320 7085 30326
rect 7027 30286 7039 30320
rect 7073 30317 7085 30320
rect 32176 30317 32182 30329
rect 7073 30289 7358 30317
rect 32137 30289 32182 30317
rect 7073 30286 7085 30289
rect 7027 30280 7085 30286
rect 7330 30255 7358 30289
rect 32176 30277 32182 30289
rect 32234 30277 32240 30329
rect 37426 30317 37454 30363
rect 45136 30317 45142 30329
rect 37426 30289 45142 30317
rect 45136 30277 45142 30289
rect 45194 30277 45200 30329
rect 7312 30243 7318 30255
rect 7273 30215 7318 30243
rect 7312 30203 7318 30215
rect 7370 30203 7376 30255
rect 1152 29996 58848 30018
rect 1152 29944 19654 29996
rect 19706 29944 19718 29996
rect 19770 29944 19782 29996
rect 19834 29944 19846 29996
rect 19898 29944 50374 29996
rect 50426 29944 50438 29996
rect 50490 29944 50502 29996
rect 50554 29944 50566 29996
rect 50618 29944 58848 29996
rect 1152 29922 58848 29944
rect 14803 29580 14861 29586
rect 14803 29546 14815 29580
rect 14849 29577 14861 29580
rect 15091 29580 15149 29586
rect 15091 29577 15103 29580
rect 14849 29549 15103 29577
rect 14849 29546 14861 29549
rect 14803 29540 14861 29546
rect 15091 29546 15103 29549
rect 15137 29577 15149 29580
rect 15137 29549 17294 29577
rect 15137 29546 15149 29549
rect 15091 29540 15149 29546
rect 12979 29506 13037 29512
rect 12979 29472 12991 29506
rect 13025 29503 13037 29506
rect 17266 29503 17294 29549
rect 28144 29503 28150 29515
rect 13025 29475 15230 29503
rect 17266 29475 28150 29503
rect 13025 29472 13037 29475
rect 12979 29466 13037 29472
rect 9136 29389 9142 29441
rect 9194 29429 9200 29441
rect 11152 29429 11158 29441
rect 9194 29401 11158 29429
rect 9194 29389 9200 29401
rect 11152 29389 11158 29401
rect 11210 29389 11216 29441
rect 15202 29429 15230 29475
rect 28144 29463 28150 29475
rect 28202 29463 28208 29515
rect 45040 29429 45046 29441
rect 15202 29401 45046 29429
rect 45040 29389 45046 29401
rect 45098 29389 45104 29441
rect 1152 29330 58848 29352
rect 1152 29278 4294 29330
rect 4346 29278 4358 29330
rect 4410 29278 4422 29330
rect 4474 29278 4486 29330
rect 4538 29278 35014 29330
rect 35066 29278 35078 29330
rect 35130 29278 35142 29330
rect 35194 29278 35206 29330
rect 35258 29278 58848 29330
rect 1152 29256 58848 29278
rect 24304 29207 24310 29219
rect 2050 29179 24310 29207
rect 2050 29068 2078 29179
rect 24304 29167 24310 29179
rect 24362 29167 24368 29219
rect 9136 29133 9142 29145
rect 8640 29105 9142 29133
rect 9136 29093 9142 29105
rect 9194 29093 9200 29145
rect 9250 29105 11102 29133
rect 1747 29062 1805 29068
rect 1747 29028 1759 29062
rect 1793 29059 1805 29062
rect 2035 29062 2093 29068
rect 2035 29059 2047 29062
rect 1793 29031 2047 29059
rect 1793 29028 1805 29031
rect 1747 29022 1805 29028
rect 2035 29028 2047 29031
rect 2081 29028 2093 29062
rect 2035 29022 2093 29028
rect 8098 28911 8126 29008
rect 9250 28911 9278 29105
rect 11074 29059 11102 29105
rect 11152 29093 11158 29145
rect 11210 29133 11216 29145
rect 20944 29133 20950 29145
rect 11210 29105 20950 29133
rect 11210 29093 11216 29105
rect 20944 29093 20950 29105
rect 21002 29093 21008 29145
rect 15280 29059 15286 29071
rect 11074 29031 15286 29059
rect 15280 29019 15286 29031
rect 15338 29019 15344 29071
rect 8098 28883 9278 28911
rect 41296 28871 41302 28923
rect 41354 28911 41360 28923
rect 44947 28914 45005 28920
rect 44947 28911 44959 28914
rect 41354 28883 44959 28911
rect 41354 28871 41360 28883
rect 44947 28880 44959 28883
rect 44993 28880 45005 28914
rect 50323 28914 50381 28920
rect 50323 28911 50335 28914
rect 44947 28874 45005 28880
rect 47506 28883 50335 28911
rect 32656 28797 32662 28849
rect 32714 28837 32720 28849
rect 47506 28837 47534 28883
rect 50323 28880 50335 28883
rect 50369 28880 50381 28914
rect 50323 28874 50381 28880
rect 32714 28809 47534 28837
rect 32714 28797 32720 28809
rect 9136 28723 9142 28775
rect 9194 28723 9200 28775
rect 1152 28664 58848 28686
rect 1152 28612 19654 28664
rect 19706 28612 19718 28664
rect 19770 28612 19782 28664
rect 19834 28612 19846 28664
rect 19898 28612 50374 28664
rect 50426 28612 50438 28664
rect 50490 28612 50502 28664
rect 50554 28612 50566 28664
rect 50618 28612 58848 28664
rect 1152 28590 58848 28612
rect 9136 28501 9142 28553
rect 9194 28541 9200 28553
rect 10864 28541 10870 28553
rect 9194 28513 10870 28541
rect 9194 28501 9200 28513
rect 10864 28501 10870 28513
rect 10922 28501 10928 28553
rect 1840 28057 1846 28109
rect 1898 28097 1904 28109
rect 22387 28100 22445 28106
rect 22387 28097 22399 28100
rect 1898 28069 22399 28097
rect 1898 28057 1904 28069
rect 22387 28066 22399 28069
rect 22433 28097 22445 28100
rect 22579 28100 22637 28106
rect 22579 28097 22591 28100
rect 22433 28069 22591 28097
rect 22433 28066 22445 28069
rect 22387 28060 22445 28066
rect 22579 28066 22591 28069
rect 22625 28066 22637 28100
rect 22579 28060 22637 28066
rect 1152 27998 58848 28020
rect 1152 27946 4294 27998
rect 4346 27946 4358 27998
rect 4410 27946 4422 27998
rect 4474 27946 4486 27998
rect 4538 27946 35014 27998
rect 35066 27946 35078 27998
rect 35130 27946 35142 27998
rect 35194 27946 35206 27998
rect 35258 27946 58848 27998
rect 1152 27924 58848 27946
rect 17584 27875 17590 27887
rect 8242 27847 17590 27875
rect 8242 27713 8270 27847
rect 17584 27835 17590 27847
rect 17642 27835 17648 27887
rect 15376 27653 15382 27665
rect 12946 27625 15382 27653
rect 8755 27582 8813 27588
rect 8755 27548 8767 27582
rect 8801 27579 8813 27582
rect 12946 27579 12974 27625
rect 15376 27613 15382 27625
rect 15434 27613 15440 27665
rect 8801 27551 12974 27579
rect 16243 27582 16301 27588
rect 8801 27548 8813 27551
rect 8755 27542 8813 27548
rect 16243 27548 16255 27582
rect 16289 27579 16301 27582
rect 22960 27579 22966 27591
rect 16289 27551 17294 27579
rect 22921 27551 22966 27579
rect 16289 27548 16301 27551
rect 16243 27542 16301 27548
rect 8467 27508 8525 27514
rect 8467 27505 8479 27508
rect 7968 27477 8479 27505
rect 8467 27474 8479 27477
rect 8513 27474 8525 27508
rect 17266 27505 17294 27551
rect 22960 27539 22966 27551
rect 23018 27539 23024 27591
rect 49648 27579 49654 27591
rect 27346 27551 49654 27579
rect 27346 27505 27374 27551
rect 49648 27539 49654 27551
rect 49706 27539 49712 27591
rect 17266 27477 27374 27505
rect 8467 27468 8525 27474
rect 20368 27431 20374 27443
rect 8640 27403 20374 27431
rect 20368 27391 20374 27403
rect 20426 27391 20432 27443
rect 1152 27332 58848 27354
rect 1152 27280 19654 27332
rect 19706 27280 19718 27332
rect 19770 27280 19782 27332
rect 19834 27280 19846 27332
rect 19898 27280 50374 27332
rect 50426 27280 50438 27332
rect 50490 27280 50502 27332
rect 50554 27280 50566 27332
rect 50618 27280 58848 27332
rect 1152 27258 58848 27280
rect 8560 26725 8566 26777
rect 8618 26765 8624 26777
rect 18160 26765 18166 26777
rect 8618 26737 18166 26765
rect 8618 26725 8624 26737
rect 18160 26725 18166 26737
rect 18218 26725 18224 26777
rect 1152 26666 58848 26688
rect 1152 26614 4294 26666
rect 4346 26614 4358 26666
rect 4410 26614 4422 26666
rect 4474 26614 4486 26666
rect 4538 26614 35014 26666
rect 35066 26614 35078 26666
rect 35130 26614 35142 26666
rect 35194 26614 35206 26666
rect 35258 26614 58848 26666
rect 1152 26592 58848 26614
rect 8224 26503 8230 26555
rect 8282 26543 8288 26555
rect 18544 26543 18550 26555
rect 8282 26515 18550 26543
rect 8282 26503 8288 26515
rect 18544 26503 18550 26515
rect 18602 26503 18608 26555
rect 18928 26469 18934 26481
rect 8770 26441 18934 26469
rect 8770 26434 8798 26441
rect 18928 26429 18934 26441
rect 18986 26429 18992 26481
rect 8230 26370 8282 26376
rect 8230 26312 8282 26318
rect 8518 26370 8570 26376
rect 8518 26312 8570 26318
rect 33520 26247 33526 26259
rect 33481 26219 33526 26247
rect 33520 26207 33526 26219
rect 33578 26207 33584 26259
rect 17392 26173 17398 26185
rect 7954 26099 7982 26159
rect 8832 26145 17398 26173
rect 17392 26133 17398 26145
rect 17450 26133 17456 26185
rect 17872 26099 17878 26111
rect 7954 26071 17878 26099
rect 17872 26059 17878 26071
rect 17930 26059 17936 26111
rect 36499 26102 36557 26108
rect 36499 26068 36511 26102
rect 36545 26099 36557 26102
rect 36787 26102 36845 26108
rect 36787 26099 36799 26102
rect 36545 26071 36799 26099
rect 36545 26068 36557 26071
rect 36499 26062 36557 26068
rect 36787 26068 36799 26071
rect 36833 26099 36845 26102
rect 40432 26099 40438 26111
rect 36833 26071 40438 26099
rect 36833 26068 36845 26071
rect 36787 26062 36845 26068
rect 40432 26059 40438 26071
rect 40490 26059 40496 26111
rect 1152 26000 58848 26022
rect 1152 25948 19654 26000
rect 19706 25948 19718 26000
rect 19770 25948 19782 26000
rect 19834 25948 19846 26000
rect 19898 25948 50374 26000
rect 50426 25948 50438 26000
rect 50490 25948 50502 26000
rect 50554 25948 50566 26000
rect 50618 25948 58848 26000
rect 1152 25926 58848 25948
rect 1152 25334 58848 25356
rect 1152 25282 4294 25334
rect 4346 25282 4358 25334
rect 4410 25282 4422 25334
rect 4474 25282 4486 25334
rect 4538 25282 35014 25334
rect 35066 25282 35078 25334
rect 35130 25282 35142 25334
rect 35194 25282 35206 25334
rect 35258 25282 58848 25334
rect 1152 25260 58848 25282
rect 16816 25137 16822 25149
rect 7824 25109 16822 25137
rect 16816 25097 16822 25109
rect 16874 25097 16880 25149
rect 8080 24841 8086 24853
rect 7968 24813 8086 24841
rect 8080 24801 8086 24813
rect 8138 24801 8144 24853
rect 11440 24841 11446 24853
rect 8242 24767 8270 24827
rect 8544 24813 11446 24841
rect 11440 24801 11446 24813
rect 11498 24801 11504 24853
rect 10768 24767 10774 24779
rect 8242 24739 10774 24767
rect 10768 24727 10774 24739
rect 10826 24727 10832 24779
rect 1152 24668 58848 24690
rect 1152 24616 19654 24668
rect 19706 24616 19718 24668
rect 19770 24616 19782 24668
rect 19834 24616 19846 24668
rect 19898 24616 50374 24668
rect 50426 24616 50438 24668
rect 50490 24616 50502 24668
rect 50554 24616 50566 24668
rect 50618 24616 58848 24668
rect 1152 24594 58848 24616
rect 8080 24505 8086 24557
rect 8138 24545 8144 24557
rect 11152 24545 11158 24557
rect 8138 24517 11158 24545
rect 8138 24505 8144 24517
rect 11152 24505 11158 24517
rect 11210 24505 11216 24557
rect 18736 24249 18742 24261
rect 2866 24221 18742 24249
rect 2227 24178 2285 24184
rect 2227 24144 2239 24178
rect 2273 24175 2285 24178
rect 2515 24178 2573 24184
rect 2515 24175 2527 24178
rect 2273 24147 2527 24175
rect 2273 24144 2285 24147
rect 2227 24138 2285 24144
rect 2515 24144 2527 24147
rect 2561 24175 2573 24178
rect 2866 24175 2894 24221
rect 18736 24209 18742 24221
rect 18794 24209 18800 24261
rect 2561 24147 2894 24175
rect 2561 24144 2573 24147
rect 2515 24138 2573 24144
rect 10960 24135 10966 24187
rect 11018 24175 11024 24187
rect 11018 24147 17294 24175
rect 11018 24135 11024 24147
rect 13360 24101 13366 24113
rect 13321 24073 13366 24101
rect 13360 24061 13366 24073
rect 13418 24061 13424 24113
rect 17266 24101 17294 24147
rect 36691 24104 36749 24110
rect 36691 24101 36703 24104
rect 17266 24073 36703 24101
rect 36691 24070 36703 24073
rect 36737 24101 36749 24104
rect 36883 24104 36941 24110
rect 36883 24101 36895 24104
rect 36737 24073 36895 24101
rect 36737 24070 36749 24073
rect 36691 24064 36749 24070
rect 36883 24070 36895 24073
rect 36929 24070 36941 24104
rect 36883 24064 36941 24070
rect 1152 24002 58848 24024
rect 1152 23950 4294 24002
rect 4346 23950 4358 24002
rect 4410 23950 4422 24002
rect 4474 23950 4486 24002
rect 4538 23950 35014 24002
rect 35066 23950 35078 24002
rect 35130 23950 35142 24002
rect 35194 23950 35206 24002
rect 35258 23950 58848 24002
rect 1152 23928 58848 23950
rect 12976 23879 12982 23891
rect 7954 23851 12982 23879
rect 7954 23717 7982 23851
rect 12976 23839 12982 23851
rect 13034 23839 13040 23891
rect 13360 23839 13366 23891
rect 13418 23879 13424 23891
rect 22672 23879 22678 23891
rect 13418 23851 22678 23879
rect 13418 23839 13424 23851
rect 22672 23839 22678 23851
rect 22730 23839 22736 23891
rect 44080 23583 44086 23595
rect 44041 23555 44086 23583
rect 44080 23543 44086 23555
rect 44138 23543 44144 23595
rect 8080 23469 8086 23521
rect 8138 23509 8144 23521
rect 8138 23481 8256 23509
rect 8138 23469 8144 23481
rect 16048 23435 16054 23447
rect 8352 23407 16054 23435
rect 16048 23395 16054 23407
rect 16106 23395 16112 23447
rect 1152 23336 58848 23358
rect 1152 23284 19654 23336
rect 19706 23284 19718 23336
rect 19770 23284 19782 23336
rect 19834 23284 19846 23336
rect 19898 23284 50374 23336
rect 50426 23284 50438 23336
rect 50490 23284 50502 23336
rect 50554 23284 50566 23336
rect 50618 23284 58848 23336
rect 1152 23262 58848 23284
rect 8080 23173 8086 23225
rect 8138 23213 8144 23225
rect 14128 23213 14134 23225
rect 8138 23185 14134 23213
rect 8138 23173 8144 23185
rect 14128 23173 14134 23185
rect 14186 23173 14192 23225
rect 7888 22729 7894 22781
rect 7946 22769 7952 22781
rect 8083 22772 8141 22778
rect 8083 22769 8095 22772
rect 7946 22741 8095 22769
rect 7946 22729 7952 22741
rect 8083 22738 8095 22741
rect 8129 22738 8141 22772
rect 8083 22732 8141 22738
rect 28531 22772 28589 22778
rect 28531 22738 28543 22772
rect 28577 22769 28589 22772
rect 44944 22769 44950 22781
rect 28577 22741 44950 22769
rect 28577 22738 28589 22741
rect 28531 22732 28589 22738
rect 44944 22729 44950 22741
rect 45002 22729 45008 22781
rect 1152 22670 58848 22692
rect 1152 22618 4294 22670
rect 4346 22618 4358 22670
rect 4410 22618 4422 22670
rect 4474 22618 4486 22670
rect 4538 22618 35014 22670
rect 35066 22618 35078 22670
rect 35130 22618 35142 22670
rect 35194 22618 35206 22670
rect 35258 22618 58848 22670
rect 1152 22596 58848 22618
rect 15472 22473 15478 22485
rect 7824 22445 15478 22473
rect 15472 22433 15478 22445
rect 15530 22433 15536 22485
rect 2608 22251 2614 22263
rect 2569 22223 2614 22251
rect 2608 22211 2614 22223
rect 2666 22211 2672 22263
rect 8080 22177 8086 22189
rect 7968 22149 8086 22177
rect 8080 22137 8086 22149
rect 8138 22137 8144 22189
rect 13168 22177 13174 22189
rect 8242 22103 8270 22163
rect 8544 22149 13174 22177
rect 13168 22137 13174 22149
rect 13226 22137 13232 22189
rect 13456 22103 13462 22115
rect 8242 22075 13462 22103
rect 13456 22063 13462 22075
rect 13514 22063 13520 22115
rect 1152 22004 58848 22026
rect 1152 21952 19654 22004
rect 19706 21952 19718 22004
rect 19770 21952 19782 22004
rect 19834 21952 19846 22004
rect 19898 21952 50374 22004
rect 50426 21952 50438 22004
rect 50490 21952 50502 22004
rect 50554 21952 50566 22004
rect 50618 21952 58848 22004
rect 1152 21930 58848 21952
rect 8080 21841 8086 21893
rect 8138 21881 8144 21893
rect 13264 21881 13270 21893
rect 8138 21853 13270 21881
rect 8138 21841 8144 21853
rect 13264 21841 13270 21853
rect 13322 21841 13328 21893
rect 31123 21884 31181 21890
rect 31123 21850 31135 21884
rect 31169 21881 31181 21884
rect 31411 21884 31469 21890
rect 31411 21881 31423 21884
rect 31169 21853 31423 21881
rect 31169 21850 31181 21853
rect 31123 21844 31181 21850
rect 31411 21850 31423 21853
rect 31457 21881 31469 21884
rect 32560 21881 32566 21893
rect 31457 21853 32566 21881
rect 31457 21850 31469 21853
rect 31411 21844 31469 21850
rect 32560 21841 32566 21853
rect 32618 21841 32624 21893
rect 2608 21693 2614 21745
rect 2666 21733 2672 21745
rect 36496 21733 36502 21745
rect 2666 21705 36502 21733
rect 2666 21693 2672 21705
rect 36496 21693 36502 21705
rect 36554 21693 36560 21745
rect 8080 21471 8086 21523
rect 8138 21511 8144 21523
rect 55408 21511 55414 21523
rect 8138 21483 55414 21511
rect 8138 21471 8144 21483
rect 55408 21471 55414 21483
rect 55466 21471 55472 21523
rect 32272 21437 32278 21449
rect 32233 21409 32278 21437
rect 32272 21397 32278 21409
rect 32330 21397 32336 21449
rect 43024 21397 43030 21449
rect 43082 21437 43088 21449
rect 58003 21440 58061 21446
rect 58003 21437 58015 21440
rect 43082 21409 58015 21437
rect 43082 21397 43088 21409
rect 58003 21406 58015 21409
rect 58049 21406 58061 21440
rect 58003 21400 58061 21406
rect 1152 21338 58848 21360
rect 1152 21286 4294 21338
rect 4346 21286 4358 21338
rect 4410 21286 4422 21338
rect 4474 21286 4486 21338
rect 4538 21286 35014 21338
rect 35066 21286 35078 21338
rect 35130 21286 35142 21338
rect 35194 21286 35206 21338
rect 35258 21286 58848 21338
rect 1152 21264 58848 21286
rect 32272 21175 32278 21227
rect 32330 21215 32336 21227
rect 44752 21215 44758 21227
rect 32330 21187 44758 21215
rect 32330 21175 32336 21187
rect 44752 21175 44758 21187
rect 44810 21175 44816 21227
rect 26416 21027 26422 21079
rect 26474 21067 26480 21079
rect 43699 21070 43757 21076
rect 43699 21067 43711 21070
rect 26474 21039 43711 21067
rect 26474 21027 26480 21039
rect 43699 21036 43711 21039
rect 43745 21067 43757 21070
rect 43891 21070 43949 21076
rect 43891 21067 43903 21070
rect 43745 21039 43903 21067
rect 43745 21036 43757 21039
rect 43699 21030 43757 21036
rect 43891 21036 43903 21039
rect 43937 21036 43949 21070
rect 43891 21030 43949 21036
rect 30928 20953 30934 21005
rect 30986 20993 30992 21005
rect 41395 20996 41453 21002
rect 41395 20993 41407 20996
rect 30986 20965 41407 20993
rect 30986 20953 30992 20965
rect 41395 20962 41407 20965
rect 41441 20962 41453 20996
rect 41395 20956 41453 20962
rect 7120 20919 7126 20931
rect 7081 20891 7126 20919
rect 7120 20879 7126 20891
rect 7178 20879 7184 20931
rect 29200 20879 29206 20931
rect 29258 20919 29264 20931
rect 34387 20922 34445 20928
rect 34387 20919 34399 20922
rect 29258 20891 34399 20919
rect 29258 20879 29264 20891
rect 34387 20888 34399 20891
rect 34433 20888 34445 20922
rect 34387 20882 34445 20888
rect 44848 20879 44854 20931
rect 44906 20919 44912 20931
rect 53392 20919 53398 20931
rect 44906 20891 53398 20919
rect 44906 20879 44912 20891
rect 53392 20879 53398 20891
rect 53450 20879 53456 20931
rect 8080 20845 8086 20857
rect 7968 20817 8086 20845
rect 8080 20805 8086 20817
rect 8138 20805 8144 20857
rect 16528 20845 16534 20857
rect 8256 20817 16534 20845
rect 16528 20805 16534 20817
rect 16586 20805 16592 20857
rect 27346 20817 47534 20845
rect 7603 20774 7661 20780
rect 7603 20740 7615 20774
rect 7649 20771 7661 20774
rect 27346 20771 27374 20817
rect 7649 20743 27374 20771
rect 47506 20771 47534 20817
rect 57712 20771 57718 20783
rect 47506 20743 57718 20771
rect 7649 20740 7661 20743
rect 7603 20734 7661 20740
rect 57712 20731 57718 20743
rect 57770 20731 57776 20783
rect 1152 20672 58848 20694
rect 1152 20620 19654 20672
rect 19706 20620 19718 20672
rect 19770 20620 19782 20672
rect 19834 20620 19846 20672
rect 19898 20620 50374 20672
rect 50426 20620 50438 20672
rect 50490 20620 50502 20672
rect 50554 20620 50566 20672
rect 50618 20620 58848 20672
rect 1152 20598 58848 20620
rect 3376 20509 3382 20561
rect 3434 20549 3440 20561
rect 9427 20552 9485 20558
rect 9427 20549 9439 20552
rect 3434 20521 9439 20549
rect 3434 20509 3440 20521
rect 9427 20518 9439 20521
rect 9473 20549 9485 20552
rect 9616 20549 9622 20561
rect 9473 20521 9622 20549
rect 9473 20518 9485 20521
rect 9427 20512 9485 20518
rect 9616 20509 9622 20521
rect 9674 20509 9680 20561
rect 12688 20509 12694 20561
rect 12746 20549 12752 20561
rect 16243 20552 16301 20558
rect 16243 20549 16255 20552
rect 12746 20521 16255 20549
rect 12746 20509 12752 20521
rect 16243 20518 16255 20521
rect 16289 20549 16301 20552
rect 16289 20521 16478 20549
rect 16289 20518 16301 20521
rect 16243 20512 16301 20518
rect 7120 20361 7126 20413
rect 7178 20401 7184 20413
rect 16240 20401 16246 20413
rect 7178 20373 16246 20401
rect 7178 20361 7184 20373
rect 16240 20361 16246 20373
rect 16298 20361 16304 20413
rect 16450 20410 16478 20521
rect 16435 20404 16493 20410
rect 16435 20370 16447 20404
rect 16481 20370 16493 20404
rect 16435 20364 16493 20370
rect 44563 20404 44621 20410
rect 44563 20370 44575 20404
rect 44609 20401 44621 20404
rect 44848 20401 44854 20413
rect 44609 20373 44854 20401
rect 44609 20370 44621 20373
rect 44563 20364 44621 20370
rect 44848 20361 44854 20373
rect 44906 20361 44912 20413
rect 9616 20327 9622 20339
rect 9577 20299 9622 20327
rect 9616 20287 9622 20299
rect 9674 20287 9680 20339
rect 10576 20105 10582 20117
rect 10537 20077 10582 20105
rect 10576 20065 10582 20077
rect 10634 20065 10640 20117
rect 13648 20065 13654 20117
rect 13706 20105 13712 20117
rect 18835 20108 18893 20114
rect 18835 20105 18847 20108
rect 13706 20077 18847 20105
rect 13706 20065 13712 20077
rect 18835 20074 18847 20077
rect 18881 20074 18893 20108
rect 42736 20105 42742 20117
rect 42697 20077 42742 20105
rect 18835 20068 18893 20074
rect 42736 20065 42742 20077
rect 42794 20065 42800 20117
rect 43792 20065 43798 20117
rect 43850 20105 43856 20117
rect 47155 20108 47213 20114
rect 47155 20105 47167 20108
rect 43850 20077 47167 20105
rect 43850 20065 43856 20077
rect 47155 20074 47167 20077
rect 47201 20074 47213 20108
rect 47155 20068 47213 20074
rect 1152 20006 58848 20028
rect 1152 19954 4294 20006
rect 4346 19954 4358 20006
rect 4410 19954 4422 20006
rect 4474 19954 4486 20006
rect 4538 19954 35014 20006
rect 35066 19954 35078 20006
rect 35130 19954 35142 20006
rect 35194 19954 35206 20006
rect 35258 19954 58848 20006
rect 1152 19932 58848 19954
rect 52816 19883 52822 19895
rect 8242 19855 52822 19883
rect 8242 19610 8270 19855
rect 52816 19843 52822 19855
rect 52874 19843 52880 19895
rect 8371 19812 8429 19818
rect 8371 19778 8383 19812
rect 8417 19809 8429 19812
rect 8417 19781 10094 19809
rect 8417 19778 8429 19781
rect 8371 19772 8429 19778
rect 10066 19661 10094 19781
rect 10576 19769 10582 19821
rect 10634 19809 10640 19821
rect 30640 19809 30646 19821
rect 10634 19781 30646 19809
rect 10634 19769 10640 19781
rect 30640 19769 30646 19781
rect 30698 19769 30704 19821
rect 55504 19661 55510 19673
rect 10066 19633 55510 19661
rect 55504 19621 55510 19633
rect 55562 19621 55568 19673
rect 45904 19587 45910 19599
rect 45865 19559 45910 19587
rect 45904 19547 45910 19559
rect 45962 19547 45968 19599
rect 52048 19547 52054 19599
rect 52106 19587 52112 19599
rect 52915 19590 52973 19596
rect 52915 19587 52927 19590
rect 52106 19559 52927 19587
rect 52106 19547 52112 19559
rect 52915 19556 52927 19559
rect 52961 19556 52973 19590
rect 54736 19587 54742 19599
rect 54697 19559 54742 19587
rect 52915 19550 52973 19556
rect 54736 19547 54742 19559
rect 54794 19547 54800 19599
rect 50800 19513 50806 19525
rect 9120 19485 50806 19513
rect 50800 19473 50806 19485
rect 50858 19473 50864 19525
rect 7603 19442 7661 19448
rect 7603 19408 7615 19442
rect 7649 19439 7661 19442
rect 8371 19442 8429 19448
rect 8371 19439 8383 19442
rect 7649 19411 8383 19439
rect 7649 19408 7661 19411
rect 7603 19402 7661 19408
rect 8371 19408 8383 19411
rect 8417 19408 8429 19442
rect 8371 19402 8429 19408
rect 8752 19399 8758 19451
rect 8810 19399 8816 19451
rect 9328 19399 9334 19451
rect 9386 19439 9392 19451
rect 48688 19439 48694 19451
rect 9386 19411 48694 19439
rect 9386 19399 9392 19411
rect 48688 19399 48694 19411
rect 48746 19399 48752 19451
rect 1152 19340 58848 19362
rect 1152 19288 19654 19340
rect 19706 19288 19718 19340
rect 19770 19288 19782 19340
rect 19834 19288 19846 19340
rect 19898 19288 50374 19340
rect 50426 19288 50438 19340
rect 50490 19288 50502 19340
rect 50554 19288 50566 19340
rect 50618 19288 58848 19340
rect 1152 19266 58848 19288
rect 8752 19177 8758 19229
rect 8810 19217 8816 19229
rect 9328 19217 9334 19229
rect 8810 19189 9334 19217
rect 8810 19177 8816 19189
rect 9328 19177 9334 19189
rect 9386 19177 9392 19229
rect 42832 19177 42838 19229
rect 42890 19217 42896 19229
rect 54736 19217 54742 19229
rect 42890 19189 54742 19217
rect 42890 19177 42896 19189
rect 54736 19177 54742 19189
rect 54794 19177 54800 19229
rect 36208 19103 36214 19155
rect 36266 19143 36272 19155
rect 45904 19143 45910 19155
rect 36266 19115 45910 19143
rect 36266 19103 36272 19115
rect 45904 19103 45910 19115
rect 45962 19103 45968 19155
rect 21040 18881 21046 18933
rect 21098 18921 21104 18933
rect 36115 18924 36173 18930
rect 36115 18921 36127 18924
rect 21098 18893 36127 18921
rect 21098 18881 21104 18893
rect 36115 18890 36127 18893
rect 36161 18921 36173 18924
rect 36307 18924 36365 18930
rect 36307 18921 36319 18924
rect 36161 18893 36319 18921
rect 36161 18890 36173 18893
rect 36115 18884 36173 18890
rect 36307 18890 36319 18893
rect 36353 18890 36365 18924
rect 36307 18884 36365 18890
rect 4531 18850 4589 18856
rect 4531 18816 4543 18850
rect 4577 18847 4589 18850
rect 21904 18847 21910 18859
rect 4577 18819 21910 18847
rect 4577 18816 4589 18819
rect 4531 18810 4589 18816
rect 21904 18807 21910 18819
rect 21962 18807 21968 18859
rect 57331 18850 57389 18856
rect 57331 18847 57343 18850
rect 36130 18819 57343 18847
rect 36130 18785 36158 18819
rect 57331 18816 57343 18819
rect 57377 18816 57389 18850
rect 57331 18810 57389 18816
rect 15091 18776 15149 18782
rect 15091 18742 15103 18776
rect 15137 18773 15149 18776
rect 25456 18773 25462 18785
rect 15137 18745 25462 18773
rect 15137 18742 15149 18745
rect 15091 18736 15149 18742
rect 25456 18733 25462 18745
rect 25514 18733 25520 18785
rect 36112 18733 36118 18785
rect 36170 18733 36176 18785
rect 39952 18773 39958 18785
rect 39913 18745 39958 18773
rect 39952 18733 39958 18745
rect 40010 18733 40016 18785
rect 1152 18674 58848 18696
rect 1152 18622 4294 18674
rect 4346 18622 4358 18674
rect 4410 18622 4422 18674
rect 4474 18622 4486 18674
rect 4538 18622 35014 18674
rect 35066 18622 35078 18674
rect 35130 18622 35142 18674
rect 35194 18622 35206 18674
rect 35258 18622 58848 18674
rect 1152 18600 58848 18622
rect 48880 18551 48886 18563
rect 7810 18523 48886 18551
rect 7603 18480 7661 18486
rect 7603 18446 7615 18480
rect 7649 18477 7661 18480
rect 7810 18477 7838 18523
rect 48880 18511 48886 18523
rect 48938 18511 48944 18563
rect 8755 18480 8813 18486
rect 8755 18477 8767 18480
rect 7649 18463 7838 18477
rect 7649 18449 7824 18463
rect 8674 18449 8767 18477
rect 7649 18446 7661 18449
rect 7603 18440 7661 18446
rect 8674 18352 8702 18449
rect 8755 18446 8767 18449
rect 8801 18446 8813 18480
rect 8755 18440 8813 18446
rect 9043 18406 9101 18412
rect 9043 18372 9055 18406
rect 9089 18403 9101 18406
rect 46096 18403 46102 18415
rect 9089 18375 46102 18403
rect 9089 18372 9101 18375
rect 9043 18366 9101 18372
rect 46096 18363 46102 18375
rect 46154 18363 46160 18415
rect 24019 18258 24077 18264
rect 24019 18224 24031 18258
rect 24065 18255 24077 18258
rect 40336 18255 40342 18267
rect 24065 18227 40342 18255
rect 24065 18224 24077 18227
rect 24019 18218 24077 18224
rect 40336 18215 40342 18227
rect 40394 18215 40400 18267
rect 44083 18258 44141 18264
rect 44083 18224 44095 18258
rect 44129 18224 44141 18258
rect 44083 18218 44141 18224
rect 44659 18258 44717 18264
rect 44659 18224 44671 18258
rect 44705 18224 44717 18258
rect 44659 18218 44717 18224
rect 9427 18184 9485 18190
rect 9427 18150 9439 18184
rect 9473 18181 9485 18184
rect 9715 18184 9773 18190
rect 9715 18181 9727 18184
rect 9473 18153 9727 18181
rect 9473 18150 9485 18153
rect 9427 18144 9485 18150
rect 9715 18150 9727 18153
rect 9761 18181 9773 18184
rect 19984 18181 19990 18193
rect 9761 18153 19990 18181
rect 9761 18150 9773 18153
rect 9715 18144 9773 18150
rect 19984 18141 19990 18153
rect 20042 18141 20048 18193
rect 34288 18141 34294 18193
rect 34346 18181 34352 18193
rect 44098 18181 44126 18218
rect 34346 18153 44126 18181
rect 34346 18141 34352 18153
rect 14032 18067 14038 18119
rect 14090 18107 14096 18119
rect 44467 18110 44525 18116
rect 44467 18107 44479 18110
rect 14090 18079 44479 18107
rect 14090 18067 14096 18079
rect 44467 18076 44479 18079
rect 44513 18107 44525 18110
rect 44674 18107 44702 18218
rect 44513 18079 44702 18107
rect 44513 18076 44525 18079
rect 44467 18070 44525 18076
rect 1152 18008 58848 18030
rect 1152 17956 19654 18008
rect 19706 17956 19718 18008
rect 19770 17956 19782 18008
rect 19834 17956 19846 18008
rect 19898 17956 50374 18008
rect 50426 17956 50438 18008
rect 50490 17956 50502 18008
rect 50554 17956 50566 18008
rect 50618 17956 58848 18008
rect 1152 17934 58848 17956
rect 32464 17549 32470 17601
rect 32522 17589 32528 17601
rect 46483 17592 46541 17598
rect 46483 17589 46495 17592
rect 32522 17561 46495 17589
rect 32522 17549 32528 17561
rect 46483 17558 46495 17561
rect 46529 17589 46541 17592
rect 46675 17592 46733 17598
rect 46675 17589 46687 17592
rect 46529 17561 46687 17589
rect 46529 17558 46541 17561
rect 46483 17552 46541 17558
rect 46675 17558 46687 17561
rect 46721 17558 46733 17592
rect 46675 17552 46733 17558
rect 57331 17518 57389 17524
rect 57331 17515 57343 17518
rect 38626 17487 57343 17515
rect 6064 17401 6070 17453
rect 6122 17441 6128 17453
rect 7411 17444 7469 17450
rect 7411 17441 7423 17444
rect 6122 17413 7423 17441
rect 6122 17401 6128 17413
rect 7411 17410 7423 17413
rect 7457 17410 7469 17444
rect 7411 17404 7469 17410
rect 18448 17401 18454 17453
rect 18506 17441 18512 17453
rect 38626 17441 38654 17487
rect 57331 17484 57343 17487
rect 57377 17484 57389 17518
rect 57331 17478 57389 17484
rect 18506 17413 38654 17441
rect 18506 17401 18512 17413
rect 1152 17342 58848 17364
rect 1152 17290 4294 17342
rect 4346 17290 4358 17342
rect 4410 17290 4422 17342
rect 4474 17290 4486 17342
rect 4538 17290 35014 17342
rect 35066 17290 35078 17342
rect 35130 17290 35142 17342
rect 35194 17290 35206 17342
rect 35258 17290 58848 17342
rect 1152 17268 58848 17290
rect 8083 17222 8141 17228
rect 8083 17188 8095 17222
rect 8129 17219 8141 17222
rect 42928 17219 42934 17231
rect 8129 17191 42934 17219
rect 8129 17188 8141 17191
rect 8083 17182 8141 17188
rect 42928 17179 42934 17191
rect 42986 17179 42992 17231
rect 8083 16926 8141 16932
rect 8083 16892 8095 16926
rect 8129 16892 8141 16926
rect 8083 16886 8141 16892
rect 8098 16835 8126 16886
rect 7603 16778 7661 16784
rect 7603 16744 7615 16778
rect 7649 16775 7661 16778
rect 45232 16775 45238 16787
rect 7649 16747 45238 16775
rect 7649 16744 7661 16747
rect 7603 16738 7661 16744
rect 45232 16735 45238 16747
rect 45290 16735 45296 16787
rect 1152 16676 58848 16698
rect 1152 16624 19654 16676
rect 19706 16624 19718 16676
rect 19770 16624 19782 16676
rect 19834 16624 19846 16676
rect 19898 16624 50374 16676
rect 50426 16624 50438 16676
rect 50490 16624 50502 16676
rect 50554 16624 50566 16676
rect 50618 16624 58848 16676
rect 1152 16602 58848 16624
rect 2323 16556 2381 16562
rect 2323 16522 2335 16556
rect 2369 16553 2381 16556
rect 2611 16556 2669 16562
rect 2611 16553 2623 16556
rect 2369 16525 2623 16553
rect 2369 16522 2381 16525
rect 2323 16516 2381 16522
rect 2611 16522 2623 16525
rect 2657 16553 2669 16556
rect 3760 16553 3766 16565
rect 2657 16525 3766 16553
rect 2657 16522 2669 16525
rect 2611 16516 2669 16522
rect 3760 16513 3766 16525
rect 3818 16513 3824 16565
rect 1744 16217 1750 16269
rect 1802 16257 1808 16269
rect 54163 16260 54221 16266
rect 54163 16257 54175 16260
rect 1802 16229 54175 16257
rect 1802 16217 1808 16229
rect 54163 16226 54175 16229
rect 54209 16226 54221 16260
rect 54163 16220 54221 16226
rect 3856 16143 3862 16195
rect 3914 16183 3920 16195
rect 14704 16183 14710 16195
rect 3914 16155 14710 16183
rect 3914 16143 3920 16155
rect 14704 16143 14710 16155
rect 14762 16143 14768 16195
rect 26800 16143 26806 16195
rect 26858 16183 26864 16195
rect 49360 16183 49366 16195
rect 26858 16155 49366 16183
rect 26858 16143 26864 16155
rect 49360 16143 49366 16155
rect 49418 16143 49424 16195
rect 16144 16069 16150 16121
rect 16202 16109 16208 16121
rect 50032 16109 50038 16121
rect 16202 16081 50038 16109
rect 16202 16069 16208 16081
rect 50032 16069 50038 16081
rect 50090 16069 50096 16121
rect 1152 16010 58848 16032
rect 1152 15958 4294 16010
rect 4346 15958 4358 16010
rect 4410 15958 4422 16010
rect 4474 15958 4486 16010
rect 4538 15958 35014 16010
rect 35066 15958 35078 16010
rect 35130 15958 35142 16010
rect 35194 15958 35206 16010
rect 35258 15958 58848 16010
rect 1152 15936 58848 15958
rect 3856 15887 3862 15899
rect 3817 15859 3862 15887
rect 3856 15847 3862 15859
rect 3914 15847 3920 15899
rect 8851 15890 8909 15896
rect 8851 15856 8863 15890
rect 8897 15887 8909 15890
rect 12976 15887 12982 15899
rect 8897 15859 12982 15887
rect 8897 15856 8909 15859
rect 8851 15850 8909 15856
rect 12976 15847 12982 15859
rect 13034 15847 13040 15899
rect 16144 15887 16150 15899
rect 16105 15859 16150 15887
rect 16144 15847 16150 15859
rect 16202 15847 16208 15899
rect 26800 15887 26806 15899
rect 26761 15859 26806 15887
rect 26800 15847 26806 15859
rect 26858 15847 26864 15899
rect 48976 15847 48982 15899
rect 49034 15887 49040 15899
rect 50131 15890 50189 15896
rect 50131 15887 50143 15890
rect 49034 15859 50143 15887
rect 49034 15847 49040 15859
rect 50131 15856 50143 15859
rect 50177 15856 50189 15890
rect 50131 15850 50189 15856
rect 39760 15517 39766 15529
rect 7968 15489 39766 15517
rect 39760 15477 39766 15489
rect 39818 15477 39824 15529
rect 7603 15446 7661 15452
rect 7603 15412 7615 15446
rect 7649 15443 7661 15446
rect 42352 15443 42358 15455
rect 7649 15415 42358 15443
rect 7649 15412 7661 15415
rect 7603 15406 7661 15412
rect 42352 15403 42358 15415
rect 42410 15403 42416 15455
rect 1152 15344 58848 15366
rect 1152 15292 19654 15344
rect 19706 15292 19718 15344
rect 19770 15292 19782 15344
rect 19834 15292 19846 15344
rect 19898 15292 50374 15344
rect 50426 15292 50438 15344
rect 50490 15292 50502 15344
rect 50554 15292 50566 15344
rect 50618 15292 58848 15344
rect 1152 15270 58848 15292
rect 2707 14928 2765 14934
rect 2707 14894 2719 14928
rect 2753 14894 2765 14928
rect 2707 14888 2765 14894
rect 2419 14854 2477 14860
rect 2419 14820 2431 14854
rect 2465 14851 2477 14854
rect 2722 14851 2750 14888
rect 9616 14885 9622 14937
rect 9674 14925 9680 14937
rect 34864 14925 34870 14937
rect 9674 14897 34870 14925
rect 9674 14885 9680 14897
rect 34864 14885 34870 14897
rect 34922 14885 34928 14937
rect 27664 14851 27670 14863
rect 2465 14823 27670 14851
rect 2465 14820 2477 14823
rect 2419 14814 2477 14820
rect 27664 14811 27670 14823
rect 27722 14811 27728 14863
rect 25651 14780 25709 14786
rect 25651 14746 25663 14780
rect 25697 14777 25709 14780
rect 27952 14777 27958 14789
rect 25697 14749 27958 14777
rect 25697 14746 25709 14749
rect 25651 14740 25709 14746
rect 27952 14737 27958 14749
rect 28010 14737 28016 14789
rect 1152 14678 58848 14700
rect 1152 14626 4294 14678
rect 4346 14626 4358 14678
rect 4410 14626 4422 14678
rect 4474 14626 4486 14678
rect 4538 14626 35014 14678
rect 35066 14626 35078 14678
rect 35130 14626 35142 14678
rect 35194 14626 35206 14678
rect 35258 14626 58848 14678
rect 1152 14604 58848 14626
rect 9616 14555 9622 14567
rect 9577 14527 9622 14555
rect 9616 14515 9622 14527
rect 9674 14515 9680 14567
rect 14611 14558 14669 14564
rect 14611 14524 14623 14558
rect 14657 14555 14669 14558
rect 41488 14555 41494 14567
rect 14657 14527 41494 14555
rect 14657 14524 14669 14527
rect 14611 14518 14669 14524
rect 41488 14515 41494 14527
rect 41546 14515 41552 14567
rect 15088 14441 15094 14493
rect 15146 14481 15152 14493
rect 49843 14484 49901 14490
rect 49843 14481 49855 14484
rect 15146 14453 49855 14481
rect 15146 14441 15152 14453
rect 49843 14450 49855 14453
rect 49889 14450 49901 14484
rect 49843 14444 49901 14450
rect 53392 14441 53398 14493
rect 53450 14481 53456 14493
rect 56371 14484 56429 14490
rect 56371 14481 56383 14484
rect 53450 14453 56383 14481
rect 53450 14441 53456 14453
rect 56371 14450 56383 14453
rect 56417 14450 56429 14484
rect 56371 14444 56429 14450
rect 27859 14410 27917 14416
rect 27859 14407 27871 14410
rect 27346 14379 27871 14407
rect 18256 14219 18262 14271
rect 18314 14259 18320 14271
rect 27346 14259 27374 14379
rect 27859 14376 27871 14379
rect 27905 14407 27917 14410
rect 28051 14410 28109 14416
rect 28051 14407 28063 14410
rect 27905 14379 28063 14407
rect 27905 14376 27917 14379
rect 27859 14370 27917 14376
rect 28051 14376 28063 14379
rect 28097 14376 28109 14410
rect 28051 14370 28109 14376
rect 36688 14333 36694 14345
rect 18314 14231 27374 14259
rect 27586 14305 36694 14333
rect 18314 14219 18320 14231
rect 27586 14185 27614 14305
rect 36688 14293 36694 14305
rect 36746 14293 36752 14345
rect 7968 14157 27614 14185
rect 27778 14157 37454 14185
rect 7603 14114 7661 14120
rect 7603 14080 7615 14114
rect 7649 14111 7661 14114
rect 27778 14111 27806 14157
rect 7649 14083 27806 14111
rect 37426 14111 37454 14157
rect 38896 14111 38902 14123
rect 37426 14083 38902 14111
rect 7649 14080 7661 14083
rect 7603 14074 7661 14080
rect 38896 14071 38902 14083
rect 38954 14071 38960 14123
rect 1152 14012 58848 14034
rect 1152 13960 19654 14012
rect 19706 13960 19718 14012
rect 19770 13960 19782 14012
rect 19834 13960 19846 14012
rect 19898 13960 50374 14012
rect 50426 13960 50438 14012
rect 50490 13960 50502 14012
rect 50554 13960 50566 14012
rect 50618 13960 58848 14012
rect 1152 13938 58848 13960
rect 21808 13849 21814 13901
rect 21866 13889 21872 13901
rect 25267 13892 25325 13898
rect 25267 13889 25279 13892
rect 21866 13861 25279 13889
rect 21866 13849 21872 13861
rect 25267 13858 25279 13861
rect 25313 13889 25325 13892
rect 25313 13861 25502 13889
rect 25313 13858 25325 13861
rect 25267 13852 25325 13858
rect 25474 13750 25502 13861
rect 25459 13744 25517 13750
rect 25459 13710 25471 13744
rect 25505 13710 25517 13744
rect 25459 13704 25517 13710
rect 53584 13479 53590 13531
rect 53642 13519 53648 13531
rect 57523 13522 57581 13528
rect 57523 13519 57535 13522
rect 53642 13491 57535 13519
rect 53642 13479 53648 13491
rect 57523 13488 57535 13491
rect 57569 13488 57581 13522
rect 57523 13482 57581 13488
rect 33232 13405 33238 13457
rect 33290 13445 33296 13457
rect 54451 13448 54509 13454
rect 54451 13445 54463 13448
rect 33290 13417 54463 13445
rect 33290 13405 33296 13417
rect 54451 13414 54463 13417
rect 54497 13414 54509 13448
rect 54451 13408 54509 13414
rect 1152 13346 58848 13368
rect 1152 13294 4294 13346
rect 4346 13294 4358 13346
rect 4410 13294 4422 13346
rect 4474 13294 4486 13346
rect 4538 13294 35014 13346
rect 35066 13294 35078 13346
rect 35130 13294 35142 13346
rect 35194 13294 35206 13346
rect 35258 13294 58848 13346
rect 1152 13272 58848 13294
rect 56656 13223 56662 13235
rect 56617 13195 56662 13223
rect 56656 13183 56662 13195
rect 56714 13223 56720 13235
rect 56755 13226 56813 13232
rect 56755 13223 56767 13226
rect 56714 13195 56767 13223
rect 56714 13183 56720 13195
rect 56755 13192 56767 13195
rect 56801 13192 56813 13226
rect 56755 13186 56813 13192
rect 7603 13152 7661 13158
rect 7603 13118 7615 13152
rect 7649 13149 7661 13152
rect 36592 13149 36598 13161
rect 7649 13121 36598 13149
rect 7649 13118 7661 13121
rect 7603 13112 7661 13118
rect 36592 13109 36598 13121
rect 36650 13109 36656 13161
rect 34096 12853 34102 12865
rect 7968 12825 34102 12853
rect 34096 12813 34102 12825
rect 34154 12813 34160 12865
rect 1152 12680 58848 12702
rect 1152 12628 19654 12680
rect 19706 12628 19718 12680
rect 19770 12628 19782 12680
rect 19834 12628 19846 12680
rect 19898 12628 50374 12680
rect 50426 12628 50438 12680
rect 50490 12628 50502 12680
rect 50554 12628 50566 12680
rect 50618 12628 58848 12680
rect 1152 12606 58848 12628
rect 57328 12557 57334 12569
rect 57289 12529 57334 12557
rect 57328 12517 57334 12529
rect 57386 12517 57392 12569
rect 16048 12483 16054 12495
rect 15970 12455 16054 12483
rect 15970 12273 15998 12455
rect 16048 12443 16054 12455
rect 16106 12443 16112 12495
rect 57346 12409 57374 12517
rect 57619 12412 57677 12418
rect 57619 12409 57631 12412
rect 57346 12381 57631 12409
rect 57619 12378 57631 12381
rect 57665 12409 57677 12412
rect 57907 12412 57965 12418
rect 57907 12409 57919 12412
rect 57665 12381 57919 12409
rect 57665 12378 57677 12381
rect 57619 12372 57677 12378
rect 57907 12378 57919 12381
rect 57953 12378 57965 12412
rect 57907 12372 57965 12378
rect 15952 12221 15958 12273
rect 16010 12221 16016 12273
rect 57520 12221 57526 12273
rect 57578 12261 57584 12273
rect 57715 12264 57773 12270
rect 57715 12261 57727 12264
rect 57578 12233 57727 12261
rect 57578 12221 57584 12233
rect 57715 12230 57727 12233
rect 57761 12230 57773 12264
rect 57715 12224 57773 12230
rect 7792 12147 7798 12199
rect 7850 12187 7856 12199
rect 10864 12187 10870 12199
rect 7850 12159 10870 12187
rect 7850 12147 7856 12159
rect 10864 12147 10870 12159
rect 10922 12147 10928 12199
rect 9520 12073 9526 12125
rect 9578 12113 9584 12125
rect 28816 12113 28822 12125
rect 9578 12085 28822 12113
rect 9578 12073 9584 12085
rect 28816 12073 28822 12085
rect 28874 12073 28880 12125
rect 37555 12116 37613 12122
rect 37555 12082 37567 12116
rect 37601 12113 37613 12116
rect 38512 12113 38518 12125
rect 37601 12085 38518 12113
rect 37601 12082 37613 12085
rect 37555 12076 37613 12082
rect 38512 12073 38518 12085
rect 38570 12073 38576 12125
rect 1152 12014 58848 12036
rect 1152 11962 4294 12014
rect 4346 11962 4358 12014
rect 4410 11962 4422 12014
rect 4474 11962 4486 12014
rect 4538 11962 35014 12014
rect 35066 11962 35078 12014
rect 35130 11962 35142 12014
rect 35194 11962 35206 12014
rect 35258 11962 58848 12014
rect 1152 11940 58848 11962
rect 56179 11894 56237 11900
rect 56179 11891 56191 11894
rect 2866 11863 56191 11891
rect 2320 11777 2326 11829
rect 2378 11817 2384 11829
rect 2866 11817 2894 11863
rect 56179 11860 56191 11863
rect 56225 11891 56237 11894
rect 56225 11863 56510 11891
rect 56225 11860 56237 11863
rect 56179 11854 56237 11860
rect 2378 11789 2894 11817
rect 7603 11820 7661 11826
rect 2378 11777 2384 11789
rect 7603 11786 7615 11820
rect 7649 11817 7661 11820
rect 7699 11820 7757 11826
rect 7699 11817 7711 11820
rect 7649 11789 7711 11817
rect 7649 11786 7661 11789
rect 7603 11780 7661 11786
rect 7699 11786 7711 11789
rect 7745 11786 7757 11820
rect 7699 11780 7757 11786
rect 7792 11777 7798 11829
rect 7850 11777 7856 11829
rect 7891 11820 7949 11826
rect 7891 11786 7903 11820
rect 7937 11817 7949 11820
rect 10480 11817 10486 11829
rect 7937 11789 10486 11817
rect 7937 11786 7949 11789
rect 7891 11780 7949 11786
rect 10480 11777 10486 11789
rect 10538 11777 10544 11829
rect 10864 11817 10870 11829
rect 10825 11789 10870 11817
rect 10864 11777 10870 11789
rect 10922 11817 10928 11829
rect 32848 11817 32854 11829
rect 10922 11789 12974 11817
rect 10922 11777 10928 11789
rect 9520 11743 9526 11755
rect 8832 11715 9526 11743
rect 9520 11703 9526 11715
rect 9578 11703 9584 11755
rect 12946 11743 12974 11789
rect 23026 11789 32854 11817
rect 23026 11743 23054 11789
rect 32848 11777 32854 11789
rect 32906 11777 32912 11829
rect 34099 11820 34157 11826
rect 34099 11786 34111 11820
rect 34145 11817 34157 11820
rect 34387 11820 34445 11826
rect 34387 11817 34399 11820
rect 34145 11789 34399 11817
rect 34145 11786 34157 11789
rect 34099 11780 34157 11786
rect 34387 11786 34399 11789
rect 34433 11817 34445 11820
rect 35824 11817 35830 11829
rect 34433 11789 35830 11817
rect 34433 11786 34445 11789
rect 34387 11780 34445 11786
rect 35824 11777 35830 11789
rect 35882 11777 35888 11829
rect 31312 11743 31318 11755
rect 12946 11715 23054 11743
rect 24994 11715 31318 11743
rect 10630 11681 10682 11687
rect 24994 11669 25022 11715
rect 31312 11703 31318 11715
rect 31370 11703 31376 11755
rect 56482 11752 56510 11863
rect 59728 11817 59734 11829
rect 56578 11789 59734 11817
rect 56578 11752 56606 11789
rect 59728 11777 59734 11789
rect 59786 11777 59792 11829
rect 56467 11746 56525 11752
rect 56467 11712 56479 11746
rect 56513 11712 56525 11746
rect 56467 11706 56525 11712
rect 56563 11746 56621 11752
rect 56563 11712 56575 11746
rect 56609 11712 56621 11746
rect 56563 11706 56621 11712
rect 57136 11703 57142 11755
rect 57194 11743 57200 11755
rect 57235 11746 57293 11752
rect 57235 11743 57247 11746
rect 57194 11715 57247 11743
rect 57194 11703 57200 11715
rect 57235 11712 57247 11715
rect 57281 11712 57293 11746
rect 57235 11706 57293 11712
rect 10682 11641 25022 11669
rect 25075 11672 25133 11678
rect 25075 11638 25087 11672
rect 25121 11669 25133 11672
rect 44080 11669 44086 11681
rect 25121 11641 44086 11669
rect 25121 11638 25133 11641
rect 25075 11632 25133 11638
rect 44080 11629 44086 11641
rect 44138 11629 44144 11681
rect 44176 11629 44182 11681
rect 44234 11669 44240 11681
rect 57331 11672 57389 11678
rect 57331 11669 57343 11672
rect 44234 11641 57343 11669
rect 44234 11629 44240 11641
rect 57331 11638 57343 11641
rect 57377 11638 57389 11672
rect 57331 11632 57389 11638
rect 10630 11623 10682 11629
rect 44272 11595 44278 11607
rect 44233 11567 44278 11595
rect 44272 11555 44278 11567
rect 44330 11555 44336 11607
rect 9520 11407 9526 11459
rect 9578 11407 9584 11459
rect 1152 11348 58848 11370
rect 1152 11296 19654 11348
rect 19706 11296 19718 11348
rect 19770 11296 19782 11348
rect 19834 11296 19846 11348
rect 19898 11296 50374 11348
rect 50426 11296 50438 11348
rect 50490 11296 50502 11348
rect 50554 11296 50566 11348
rect 50618 11296 58848 11348
rect 1152 11274 58848 11296
rect 5200 11225 5206 11237
rect 5161 11197 5206 11225
rect 5200 11185 5206 11197
rect 5258 11185 5264 11237
rect 9520 11185 9526 11237
rect 9578 11225 9584 11237
rect 27184 11225 27190 11237
rect 9578 11197 27190 11225
rect 9578 11185 9584 11197
rect 27184 11185 27190 11197
rect 27242 11185 27248 11237
rect 56944 11225 56950 11237
rect 56905 11197 56950 11225
rect 56944 11185 56950 11197
rect 57002 11185 57008 11237
rect 5218 11077 5246 11185
rect 5395 11080 5453 11086
rect 5395 11077 5407 11080
rect 5218 11049 5407 11077
rect 5395 11046 5407 11049
rect 5441 11046 5453 11080
rect 56962 11077 56990 11185
rect 57235 11080 57293 11086
rect 57235 11077 57247 11080
rect 56962 11049 57247 11077
rect 5395 11040 5453 11046
rect 57235 11046 57247 11049
rect 57281 11077 57293 11080
rect 57523 11080 57581 11086
rect 57523 11077 57535 11080
rect 57281 11049 57535 11077
rect 57281 11046 57293 11049
rect 57235 11040 57293 11046
rect 57523 11046 57535 11049
rect 57569 11046 57581 11080
rect 57523 11040 57581 11046
rect 8080 10963 8086 11015
rect 8138 11003 8144 11015
rect 24016 11003 24022 11015
rect 8138 10975 24022 11003
rect 8138 10963 8144 10975
rect 24016 10963 24022 10975
rect 24074 10963 24080 11015
rect 48403 11006 48461 11012
rect 48403 10972 48415 11006
rect 48449 11003 48461 11006
rect 56083 11006 56141 11012
rect 56083 11003 56095 11006
rect 48449 10975 56095 11003
rect 48449 10972 48461 10975
rect 48403 10966 48461 10972
rect 56083 10972 56095 10975
rect 56129 10972 56141 11006
rect 56083 10966 56141 10972
rect 34579 10932 34637 10938
rect 34579 10898 34591 10932
rect 34625 10929 34637 10932
rect 34867 10932 34925 10938
rect 34867 10929 34879 10932
rect 34625 10901 34879 10929
rect 34625 10898 34637 10901
rect 34579 10892 34637 10898
rect 34867 10898 34879 10901
rect 34913 10929 34925 10932
rect 55987 10932 56045 10938
rect 34913 10901 37454 10929
rect 34913 10898 34925 10901
rect 34867 10892 34925 10898
rect 8272 10815 8278 10867
rect 8330 10855 8336 10867
rect 15760 10855 15766 10867
rect 8330 10827 15766 10855
rect 8330 10815 8336 10827
rect 15760 10815 15766 10827
rect 15818 10815 15824 10867
rect 37426 10855 37454 10901
rect 55987 10898 55999 10932
rect 56033 10929 56045 10932
rect 56368 10929 56374 10941
rect 56033 10901 56374 10929
rect 56033 10898 56045 10901
rect 55987 10892 56045 10898
rect 56368 10889 56374 10901
rect 56426 10889 56432 10941
rect 56752 10889 56758 10941
rect 56810 10929 56816 10941
rect 57331 10932 57389 10938
rect 57331 10929 57343 10932
rect 56810 10901 57343 10929
rect 56810 10889 56816 10901
rect 57331 10898 57343 10901
rect 57377 10898 57389 10932
rect 57331 10892 57389 10898
rect 54448 10855 54454 10867
rect 23026 10827 35006 10855
rect 37426 10827 54454 10855
rect 6736 10741 6742 10793
rect 6794 10781 6800 10793
rect 10672 10781 10678 10793
rect 6794 10753 10678 10781
rect 6794 10741 6800 10753
rect 10672 10741 10678 10753
rect 10730 10741 10736 10793
rect 15088 10741 15094 10793
rect 15146 10781 15152 10793
rect 23026 10781 23054 10827
rect 15146 10753 23054 10781
rect 34978 10781 35006 10827
rect 54448 10815 54454 10827
rect 54506 10815 54512 10867
rect 42643 10784 42701 10790
rect 42643 10781 42655 10784
rect 34978 10753 42655 10781
rect 15146 10741 15152 10753
rect 42643 10750 42655 10753
rect 42689 10750 42701 10784
rect 42643 10744 42701 10750
rect 1152 10682 58848 10704
rect 1152 10630 4294 10682
rect 4346 10630 4358 10682
rect 4410 10630 4422 10682
rect 4474 10630 4486 10682
rect 4538 10630 35014 10682
rect 35066 10630 35078 10682
rect 35130 10630 35142 10682
rect 35194 10630 35206 10682
rect 35258 10630 58848 10682
rect 1152 10608 58848 10630
rect 4627 10562 4685 10568
rect 4627 10528 4639 10562
rect 4673 10559 4685 10562
rect 10192 10559 10198 10571
rect 4673 10531 10198 10559
rect 4673 10528 4685 10531
rect 4627 10522 4685 10528
rect 10192 10519 10198 10531
rect 10250 10519 10256 10571
rect 10672 10519 10678 10571
rect 10730 10559 10736 10571
rect 55603 10562 55661 10568
rect 10730 10531 43214 10559
rect 10730 10519 10736 10531
rect 43186 10485 43214 10531
rect 55603 10528 55615 10562
rect 55649 10559 55661 10562
rect 56080 10559 56086 10571
rect 55649 10531 56086 10559
rect 55649 10528 55661 10531
rect 55603 10522 55661 10528
rect 43186 10457 55454 10485
rect 25648 10371 25654 10423
rect 25706 10411 25712 10423
rect 25706 10383 55358 10411
rect 25706 10371 25712 10383
rect 8080 10337 8086 10349
rect 7954 10309 8086 10337
rect 7954 10286 7982 10309
rect 8080 10297 8086 10309
rect 8138 10297 8144 10349
rect 24688 10297 24694 10349
rect 24746 10337 24752 10349
rect 46099 10340 46157 10346
rect 46099 10337 46111 10340
rect 24746 10309 46111 10337
rect 24746 10297 24752 10309
rect 46099 10306 46111 10309
rect 46145 10306 46157 10340
rect 46099 10300 46157 10306
rect 38800 10263 38806 10275
rect 38761 10235 38806 10263
rect 38800 10223 38806 10235
rect 38858 10223 38864 10275
rect 55027 10266 55085 10272
rect 55027 10232 55039 10266
rect 55073 10232 55085 10266
rect 55330 10263 55358 10383
rect 55426 10337 55454 10457
rect 55810 10420 55838 10531
rect 56080 10519 56086 10531
rect 56138 10519 56144 10571
rect 55795 10414 55853 10420
rect 55795 10380 55807 10414
rect 55841 10380 55853 10414
rect 55795 10374 55853 10380
rect 56464 10371 56470 10423
rect 56522 10411 56528 10423
rect 57427 10414 57485 10420
rect 57427 10411 57439 10414
rect 56522 10383 57439 10411
rect 56522 10371 56528 10383
rect 57427 10380 57439 10383
rect 57473 10380 57485 10414
rect 57427 10374 57485 10380
rect 56275 10340 56333 10346
rect 56275 10337 56287 10340
rect 55426 10309 56287 10337
rect 56275 10306 56287 10309
rect 56321 10337 56333 10340
rect 56563 10340 56621 10346
rect 56563 10337 56575 10340
rect 56321 10309 56575 10337
rect 56321 10306 56333 10309
rect 56275 10300 56333 10306
rect 56563 10306 56575 10309
rect 56609 10306 56621 10340
rect 56563 10300 56621 10306
rect 57043 10266 57101 10272
rect 57043 10263 57055 10266
rect 55330 10235 57055 10263
rect 55027 10226 55085 10232
rect 57043 10232 57055 10235
rect 57089 10263 57101 10266
rect 57331 10266 57389 10272
rect 57331 10263 57343 10266
rect 57089 10235 57343 10263
rect 57089 10232 57101 10235
rect 57043 10226 57101 10232
rect 57331 10232 57343 10235
rect 57377 10232 57389 10266
rect 57331 10226 57389 10232
rect 29776 10149 29782 10201
rect 29834 10189 29840 10201
rect 54739 10192 54797 10198
rect 54739 10189 54751 10192
rect 29834 10161 54751 10189
rect 29834 10149 29840 10161
rect 54739 10158 54751 10161
rect 54785 10189 54797 10192
rect 55042 10189 55070 10226
rect 58576 10189 58582 10201
rect 54785 10161 55070 10189
rect 55138 10161 58582 10189
rect 54785 10158 54797 10161
rect 54739 10152 54797 10158
rect 7603 10118 7661 10124
rect 7603 10084 7615 10118
rect 7649 10115 7661 10118
rect 26512 10115 26518 10127
rect 7649 10087 26518 10115
rect 7649 10084 7661 10087
rect 7603 10078 7661 10084
rect 26512 10075 26518 10087
rect 26570 10075 26576 10127
rect 55138 10124 55166 10161
rect 58576 10149 58582 10161
rect 58634 10149 58640 10201
rect 55123 10118 55181 10124
rect 55123 10084 55135 10118
rect 55169 10084 55181 10118
rect 55123 10078 55181 10084
rect 55696 10075 55702 10127
rect 55754 10115 55760 10127
rect 55891 10118 55949 10124
rect 55891 10115 55903 10118
rect 55754 10087 55903 10115
rect 55754 10075 55760 10087
rect 55891 10084 55903 10087
rect 55937 10084 55949 10118
rect 55891 10078 55949 10084
rect 56080 10075 56086 10127
rect 56138 10115 56144 10127
rect 56659 10118 56717 10124
rect 56659 10115 56671 10118
rect 56138 10087 56671 10115
rect 56138 10075 56144 10087
rect 56659 10084 56671 10087
rect 56705 10084 56717 10118
rect 56659 10078 56717 10084
rect 1152 10016 58848 10038
rect 1152 9964 19654 10016
rect 19706 9964 19718 10016
rect 19770 9964 19782 10016
rect 19834 9964 19846 10016
rect 19898 9964 50374 10016
rect 50426 9964 50438 10016
rect 50490 9964 50502 10016
rect 50554 9964 50566 10016
rect 50618 9964 58848 10016
rect 1152 9942 58848 9964
rect 8176 9853 8182 9905
rect 8234 9893 8240 9905
rect 23440 9893 23446 9905
rect 8234 9865 23446 9893
rect 8234 9853 8240 9865
rect 23440 9853 23446 9865
rect 23498 9853 23504 9905
rect 54163 9896 54221 9902
rect 54163 9862 54175 9896
rect 54209 9893 54221 9896
rect 54640 9893 54646 9905
rect 54209 9865 54646 9893
rect 54209 9862 54221 9865
rect 54163 9856 54221 9862
rect 8368 9705 8374 9757
rect 8426 9745 8432 9757
rect 20848 9745 20854 9757
rect 8426 9717 20854 9745
rect 8426 9705 8432 9717
rect 20848 9705 20854 9717
rect 20906 9705 20912 9757
rect 54370 9754 54398 9865
rect 54640 9853 54646 9865
rect 54698 9853 54704 9905
rect 55600 9893 55606 9905
rect 55561 9865 55606 9893
rect 55600 9853 55606 9865
rect 55658 9853 55664 9905
rect 54355 9748 54413 9754
rect 54355 9714 54367 9748
rect 54401 9714 54413 9748
rect 55618 9745 55646 9853
rect 55987 9748 56045 9754
rect 55987 9745 55999 9748
rect 55618 9717 55999 9745
rect 54355 9708 54413 9714
rect 55987 9714 55999 9717
rect 56033 9714 56045 9748
rect 55987 9708 56045 9714
rect 8080 9631 8086 9683
rect 8138 9671 8144 9683
rect 19312 9671 19318 9683
rect 8138 9643 19318 9671
rect 8138 9631 8144 9643
rect 19312 9631 19318 9643
rect 19370 9631 19376 9683
rect 57616 9671 57622 9683
rect 57577 9643 57622 9671
rect 57616 9631 57622 9643
rect 57674 9631 57680 9683
rect 8656 9557 8662 9609
rect 8714 9597 8720 9609
rect 13360 9597 13366 9609
rect 8714 9569 13366 9597
rect 8714 9557 8720 9569
rect 13360 9557 13366 9569
rect 13418 9557 13424 9609
rect 17296 9557 17302 9609
rect 17354 9597 17360 9609
rect 36784 9597 36790 9609
rect 17354 9569 36790 9597
rect 17354 9557 17360 9569
rect 36784 9557 36790 9569
rect 36842 9557 36848 9609
rect 54256 9557 54262 9609
rect 54314 9597 54320 9609
rect 54451 9600 54509 9606
rect 54451 9597 54463 9600
rect 54314 9569 54463 9597
rect 54314 9557 54320 9569
rect 54451 9566 54463 9569
rect 54497 9566 54509 9600
rect 55123 9600 55181 9606
rect 55123 9597 55135 9600
rect 54451 9560 54509 9566
rect 54850 9569 55135 9597
rect 5683 9526 5741 9532
rect 5683 9492 5695 9526
rect 5729 9523 5741 9526
rect 11536 9523 11542 9535
rect 5729 9495 11542 9523
rect 5729 9492 5741 9495
rect 5683 9486 5741 9492
rect 11536 9483 11542 9495
rect 11594 9483 11600 9535
rect 24304 9483 24310 9535
rect 24362 9523 24368 9535
rect 50704 9523 50710 9535
rect 24362 9495 50710 9523
rect 24362 9483 24368 9495
rect 50704 9483 50710 9495
rect 50762 9483 50768 9535
rect 10672 9409 10678 9461
rect 10730 9449 10736 9461
rect 17968 9449 17974 9461
rect 10730 9421 17974 9449
rect 10730 9409 10736 9421
rect 17968 9409 17974 9421
rect 18026 9409 18032 9461
rect 25360 9409 25366 9461
rect 25418 9449 25424 9461
rect 28627 9452 28685 9458
rect 28627 9449 28639 9452
rect 25418 9421 28639 9449
rect 25418 9409 25424 9421
rect 28627 9418 28639 9421
rect 28673 9418 28685 9452
rect 28627 9412 28685 9418
rect 36787 9452 36845 9458
rect 36787 9418 36799 9452
rect 36833 9449 36845 9452
rect 37264 9449 37270 9461
rect 36833 9421 37270 9449
rect 36833 9418 36845 9421
rect 36787 9412 36845 9418
rect 37264 9409 37270 9421
rect 37322 9409 37328 9461
rect 48208 9409 48214 9461
rect 48266 9449 48272 9461
rect 54850 9458 54878 9569
rect 55123 9566 55135 9569
rect 55169 9566 55181 9600
rect 55123 9560 55181 9566
rect 55219 9600 55277 9606
rect 55219 9566 55231 9600
rect 55265 9566 55277 9600
rect 55219 9560 55277 9566
rect 54928 9483 54934 9535
rect 54986 9523 54992 9535
rect 55234 9523 55262 9560
rect 55504 9557 55510 9609
rect 55562 9597 55568 9609
rect 55891 9600 55949 9606
rect 55891 9597 55903 9600
rect 55562 9569 55903 9597
rect 55562 9557 55568 9569
rect 55891 9566 55903 9569
rect 55937 9566 55949 9600
rect 55891 9560 55949 9566
rect 54986 9495 55262 9523
rect 54986 9483 54992 9495
rect 54835 9452 54893 9458
rect 54835 9449 54847 9452
rect 48266 9421 54847 9449
rect 48266 9409 48272 9421
rect 54835 9418 54847 9421
rect 54881 9418 54893 9452
rect 54835 9412 54893 9418
rect 1152 9350 58848 9372
rect 1152 9298 4294 9350
rect 4346 9298 4358 9350
rect 4410 9298 4422 9350
rect 4474 9298 4486 9350
rect 4538 9298 35014 9350
rect 35066 9298 35078 9350
rect 35130 9298 35142 9350
rect 35194 9298 35206 9350
rect 35258 9298 58848 9350
rect 1152 9276 58848 9298
rect 10672 9227 10678 9239
rect 8530 9199 10678 9227
rect 7603 9156 7661 9162
rect 7603 9122 7615 9156
rect 7649 9153 7661 9156
rect 8176 9153 8182 9165
rect 7649 9125 8182 9153
rect 7649 9122 7661 9125
rect 7603 9116 7661 9122
rect 8176 9113 8182 9125
rect 8234 9113 8240 9165
rect 8080 9079 8086 9091
rect 7968 9051 8086 9079
rect 8080 9039 8086 9051
rect 8138 9039 8144 9091
rect 8368 9079 8374 9091
rect 8256 9051 8374 9079
rect 8368 9039 8374 9051
rect 8426 9039 8432 9091
rect 8530 9065 8558 9199
rect 10672 9187 10678 9199
rect 10730 9187 10736 9239
rect 12016 9227 12022 9239
rect 11977 9199 12022 9227
rect 12016 9187 12022 9199
rect 12074 9227 12080 9239
rect 12403 9230 12461 9236
rect 12403 9227 12415 9230
rect 12074 9199 12415 9227
rect 12074 9187 12080 9199
rect 12403 9196 12415 9199
rect 12449 9196 12461 9230
rect 12403 9190 12461 9196
rect 9619 9156 9677 9162
rect 9619 9122 9631 9156
rect 9665 9153 9677 9156
rect 9907 9156 9965 9162
rect 9907 9153 9919 9156
rect 9665 9125 9919 9153
rect 9665 9122 9677 9125
rect 9619 9116 9677 9122
rect 9907 9122 9919 9125
rect 9953 9153 9965 9156
rect 48208 9153 48214 9165
rect 9953 9125 48214 9153
rect 9953 9122 9965 9125
rect 9907 9116 9965 9122
rect 48208 9113 48214 9125
rect 48266 9113 48272 9165
rect 55027 9156 55085 9162
rect 55027 9153 55039 9156
rect 53266 9125 55039 9153
rect 16336 9079 16342 9091
rect 8832 9051 16342 9079
rect 16336 9039 16342 9051
rect 16394 9039 16400 9091
rect 22960 9039 22966 9091
rect 23018 9079 23024 9091
rect 53266 9079 53294 9125
rect 55027 9122 55039 9125
rect 55073 9153 55085 9156
rect 55073 9125 55358 9153
rect 55073 9122 55085 9125
rect 55027 9116 55085 9122
rect 53392 9079 53398 9091
rect 23018 9051 53294 9079
rect 53353 9051 53398 9079
rect 23018 9039 23024 9051
rect 53392 9039 53398 9051
rect 53450 9039 53456 9091
rect 55330 9088 55358 9125
rect 55315 9082 55373 9088
rect 55315 9048 55327 9082
rect 55361 9048 55373 9082
rect 55315 9042 55373 9048
rect 12976 8965 12982 9017
rect 13034 9005 13040 9017
rect 54259 9008 54317 9014
rect 54259 9005 54271 9008
rect 13034 8977 54271 9005
rect 13034 8965 13040 8977
rect 54259 8974 54271 8977
rect 54305 9005 54317 9008
rect 54547 9008 54605 9014
rect 54547 9005 54559 9008
rect 54305 8977 54559 9005
rect 54305 8974 54317 8977
rect 54259 8968 54317 8974
rect 54547 8974 54559 8977
rect 54593 8974 54605 9008
rect 54547 8968 54605 8974
rect 56563 9008 56621 9014
rect 56563 8974 56575 9008
rect 56609 9005 56621 9008
rect 56848 9005 56854 9017
rect 56609 8977 56854 9005
rect 56609 8974 56621 8977
rect 56563 8968 56621 8974
rect 56848 8965 56854 8977
rect 56906 8965 56912 9017
rect 57232 9005 57238 9017
rect 57193 8977 57238 9005
rect 57232 8965 57238 8977
rect 57290 8965 57296 9017
rect 13744 8891 13750 8943
rect 13802 8931 13808 8943
rect 46288 8931 46294 8943
rect 13802 8903 23054 8931
rect 46249 8903 46294 8931
rect 13802 8891 13808 8903
rect 16720 8817 16726 8869
rect 16778 8857 16784 8869
rect 18064 8857 18070 8869
rect 16778 8829 18070 8857
rect 16778 8817 16784 8829
rect 18064 8817 18070 8829
rect 18122 8817 18128 8869
rect 8080 8743 8086 8795
rect 8138 8743 8144 8795
rect 16816 8743 16822 8795
rect 16874 8783 16880 8795
rect 17680 8783 17686 8795
rect 16874 8755 17686 8783
rect 16874 8743 16880 8755
rect 17680 8743 17686 8755
rect 17738 8743 17744 8795
rect 23026 8783 23054 8903
rect 46288 8891 46294 8903
rect 46346 8891 46352 8943
rect 55984 8931 55990 8943
rect 53314 8903 55990 8931
rect 49744 8817 49750 8869
rect 49802 8857 49808 8869
rect 50224 8857 50230 8869
rect 49802 8829 50230 8857
rect 49802 8817 49808 8829
rect 50224 8817 50230 8829
rect 50282 8817 50288 8869
rect 53314 8792 53342 8903
rect 55984 8891 55990 8903
rect 56042 8891 56048 8943
rect 54544 8817 54550 8869
rect 54602 8857 54608 8869
rect 54602 8829 55454 8857
rect 54602 8817 54608 8829
rect 51283 8786 51341 8792
rect 51283 8783 51295 8786
rect 23026 8755 51295 8783
rect 51283 8752 51295 8755
rect 51329 8783 51341 8786
rect 51475 8786 51533 8792
rect 51475 8783 51487 8786
rect 51329 8755 51487 8783
rect 51329 8752 51341 8755
rect 51283 8746 51341 8752
rect 51475 8752 51487 8755
rect 51521 8752 51533 8786
rect 51475 8746 51533 8752
rect 53299 8786 53357 8792
rect 53299 8752 53311 8786
rect 53345 8752 53357 8786
rect 53299 8746 53357 8752
rect 53872 8743 53878 8795
rect 53930 8783 53936 8795
rect 55426 8792 55454 8829
rect 54643 8786 54701 8792
rect 54643 8783 54655 8786
rect 53930 8755 54655 8783
rect 53930 8743 53936 8755
rect 54643 8752 54655 8755
rect 54689 8752 54701 8786
rect 54643 8746 54701 8752
rect 55411 8786 55469 8792
rect 55411 8752 55423 8786
rect 55457 8752 55469 8786
rect 55411 8746 55469 8752
rect 1152 8684 58848 8706
rect 1152 8632 19654 8684
rect 19706 8632 19718 8684
rect 19770 8632 19782 8684
rect 19834 8632 19846 8684
rect 19898 8632 50374 8684
rect 50426 8632 50438 8684
rect 50490 8632 50502 8684
rect 50554 8632 50566 8684
rect 50618 8632 58848 8684
rect 1152 8610 58848 8632
rect 9904 8521 9910 8573
rect 9962 8561 9968 8573
rect 9962 8533 11870 8561
rect 9962 8521 9968 8533
rect 11728 8487 11734 8499
rect 4546 8459 11734 8487
rect 1744 8413 1750 8425
rect 1705 8385 1750 8413
rect 1744 8373 1750 8385
rect 1802 8373 1808 8425
rect 2227 8416 2285 8422
rect 2227 8382 2239 8416
rect 2273 8413 2285 8416
rect 2416 8413 2422 8425
rect 2273 8385 2422 8413
rect 2273 8382 2285 8385
rect 2227 8376 2285 8382
rect 2416 8373 2422 8385
rect 2474 8373 2480 8425
rect 2995 8416 3053 8422
rect 2995 8382 3007 8416
rect 3041 8413 3053 8416
rect 3280 8413 3286 8425
rect 3041 8385 3286 8413
rect 3041 8382 3053 8385
rect 2995 8376 3053 8382
rect 3280 8373 3286 8385
rect 3338 8373 3344 8425
rect 4546 8422 4574 8459
rect 11728 8447 11734 8459
rect 11786 8447 11792 8499
rect 4531 8416 4589 8422
rect 4531 8382 4543 8416
rect 4577 8382 4589 8416
rect 4531 8376 4589 8382
rect 7792 8373 7798 8425
rect 7850 8413 7856 8425
rect 7891 8416 7949 8422
rect 7891 8413 7903 8416
rect 7850 8385 7903 8413
rect 7850 8373 7856 8385
rect 7891 8382 7903 8385
rect 7937 8382 7949 8416
rect 7891 8376 7949 8382
rect 10288 8373 10294 8425
rect 10346 8413 10352 8425
rect 10499 8416 10557 8422
rect 10499 8413 10511 8416
rect 10346 8385 10511 8413
rect 10346 8373 10352 8385
rect 10499 8382 10511 8385
rect 10545 8382 10557 8416
rect 10499 8376 10557 8382
rect 11059 8416 11117 8422
rect 11059 8382 11071 8416
rect 11105 8413 11117 8416
rect 11344 8413 11350 8425
rect 11105 8385 11350 8413
rect 11105 8382 11117 8385
rect 11059 8376 11117 8382
rect 11344 8373 11350 8385
rect 11402 8373 11408 8425
rect 11842 8413 11870 8533
rect 12208 8521 12214 8573
rect 12266 8561 12272 8573
rect 12883 8564 12941 8570
rect 12883 8561 12895 8564
rect 12266 8533 12895 8561
rect 12266 8521 12272 8533
rect 12883 8530 12895 8533
rect 12929 8530 12941 8564
rect 12883 8524 12941 8530
rect 15955 8564 16013 8570
rect 15955 8530 15967 8564
rect 16001 8561 16013 8564
rect 16048 8561 16054 8573
rect 16001 8533 16054 8561
rect 16001 8530 16013 8533
rect 15955 8524 16013 8530
rect 16048 8521 16054 8533
rect 16106 8521 16112 8573
rect 34672 8561 34678 8573
rect 23026 8533 34678 8561
rect 11920 8447 11926 8499
rect 11978 8487 11984 8499
rect 23026 8487 23054 8533
rect 34672 8521 34678 8533
rect 34730 8521 34736 8573
rect 48592 8561 48598 8573
rect 48553 8533 48598 8561
rect 48592 8521 48598 8533
rect 48650 8521 48656 8573
rect 50128 8521 50134 8573
rect 50186 8561 50192 8573
rect 52147 8564 52205 8570
rect 52147 8561 52159 8564
rect 50186 8533 52159 8561
rect 50186 8521 50192 8533
rect 52147 8530 52159 8533
rect 52193 8530 52205 8564
rect 52912 8561 52918 8573
rect 52873 8533 52918 8561
rect 52147 8524 52205 8530
rect 11978 8459 23054 8487
rect 32578 8459 43214 8487
rect 11978 8447 11984 8459
rect 12115 8416 12173 8422
rect 12115 8413 12127 8416
rect 11842 8385 12127 8413
rect 12115 8382 12127 8385
rect 12161 8382 12173 8416
rect 13648 8413 13654 8425
rect 13609 8385 13654 8413
rect 12115 8376 12173 8382
rect 13648 8373 13654 8385
rect 13706 8373 13712 8425
rect 16048 8373 16054 8425
rect 16106 8413 16112 8425
rect 16243 8416 16301 8422
rect 16243 8413 16255 8416
rect 16106 8385 16255 8413
rect 16106 8373 16112 8385
rect 16243 8382 16255 8385
rect 16289 8382 16301 8416
rect 20080 8413 20086 8425
rect 16243 8376 16301 8382
rect 16354 8385 20086 8413
rect 7600 8299 7606 8351
rect 7658 8339 7664 8351
rect 8272 8339 8278 8351
rect 7658 8311 8278 8339
rect 7658 8299 7664 8311
rect 8272 8299 8278 8311
rect 8330 8299 8336 8351
rect 9427 8342 9485 8348
rect 9427 8308 9439 8342
rect 9473 8339 9485 8342
rect 9811 8342 9869 8348
rect 9811 8339 9823 8342
rect 9473 8311 9823 8339
rect 9473 8308 9485 8311
rect 9427 8302 9485 8308
rect 9811 8308 9823 8311
rect 9857 8339 9869 8342
rect 16354 8339 16382 8385
rect 20080 8373 20086 8385
rect 20138 8373 20144 8425
rect 25648 8413 25654 8425
rect 25609 8385 25654 8413
rect 25648 8373 25654 8385
rect 25706 8373 25712 8425
rect 32578 8422 32606 8459
rect 32563 8416 32621 8422
rect 32563 8382 32575 8416
rect 32609 8382 32621 8416
rect 32563 8376 32621 8382
rect 9857 8311 16382 8339
rect 9857 8308 9869 8311
rect 9811 8302 9869 8308
rect 16816 8299 16822 8351
rect 16874 8339 16880 8351
rect 17011 8342 17069 8348
rect 17011 8339 17023 8342
rect 16874 8311 17023 8339
rect 16874 8299 16880 8311
rect 17011 8308 17023 8311
rect 17057 8308 17069 8342
rect 23536 8339 23542 8351
rect 17011 8302 17069 8308
rect 17266 8311 23542 8339
rect 1648 8265 1654 8277
rect 1609 8237 1654 8265
rect 1648 8225 1654 8237
rect 1706 8225 1712 8277
rect 2515 8268 2573 8274
rect 2515 8234 2527 8268
rect 2561 8234 2573 8268
rect 2515 8228 2573 8234
rect 3187 8268 3245 8274
rect 3187 8234 3199 8268
rect 3233 8265 3245 8268
rect 3280 8265 3286 8277
rect 3233 8237 3286 8265
rect 3233 8234 3245 8237
rect 3187 8228 3245 8234
rect 2224 8151 2230 8203
rect 2282 8191 2288 8203
rect 2530 8191 2558 8228
rect 3280 8225 3286 8237
rect 3338 8225 3344 8277
rect 4435 8268 4493 8274
rect 4435 8234 4447 8268
rect 4481 8234 4493 8268
rect 4435 8228 4493 8234
rect 2282 8163 2558 8191
rect 4450 8191 4478 8228
rect 7696 8225 7702 8277
rect 7754 8265 7760 8277
rect 7795 8268 7853 8274
rect 7795 8265 7807 8268
rect 7754 8237 7807 8265
rect 7754 8225 7760 8237
rect 7795 8234 7807 8237
rect 7841 8234 7853 8268
rect 7795 8228 7853 8234
rect 9520 8225 9526 8277
rect 9578 8265 9584 8277
rect 9715 8268 9773 8274
rect 9715 8265 9727 8268
rect 9578 8237 9727 8265
rect 9578 8225 9584 8237
rect 9715 8234 9727 8237
rect 9761 8234 9773 8268
rect 10576 8265 10582 8277
rect 10537 8237 10582 8265
rect 9715 8228 9773 8234
rect 10576 8225 10582 8237
rect 10634 8225 10640 8277
rect 10672 8225 10678 8277
rect 10730 8265 10736 8277
rect 11251 8268 11309 8274
rect 11251 8265 11263 8268
rect 10730 8237 11263 8265
rect 10730 8225 10736 8237
rect 11251 8234 11263 8237
rect 11297 8234 11309 8268
rect 11251 8228 11309 8234
rect 11344 8225 11350 8277
rect 11402 8265 11408 8277
rect 12019 8268 12077 8274
rect 12019 8265 12031 8268
rect 11402 8237 12031 8265
rect 11402 8225 11408 8237
rect 12019 8234 12031 8237
rect 12065 8234 12077 8268
rect 12019 8228 12077 8234
rect 12304 8225 12310 8277
rect 12362 8265 12368 8277
rect 12499 8268 12557 8274
rect 12499 8265 12511 8268
rect 12362 8237 12511 8265
rect 12362 8225 12368 8237
rect 12499 8234 12511 8237
rect 12545 8265 12557 8268
rect 12787 8268 12845 8274
rect 12787 8265 12799 8268
rect 12545 8237 12799 8265
rect 12545 8234 12557 8237
rect 12499 8228 12557 8234
rect 12787 8234 12799 8237
rect 12833 8234 12845 8268
rect 12787 8228 12845 8234
rect 12880 8225 12886 8277
rect 12938 8265 12944 8277
rect 13555 8268 13613 8274
rect 13555 8265 13567 8268
rect 12938 8237 13567 8265
rect 12938 8225 12944 8237
rect 13555 8234 13567 8237
rect 13601 8234 13613 8268
rect 13555 8228 13613 8234
rect 16048 8225 16054 8277
rect 16106 8265 16112 8277
rect 16147 8268 16205 8274
rect 16147 8265 16159 8268
rect 16106 8237 16159 8265
rect 16106 8225 16112 8237
rect 16147 8234 16159 8237
rect 16193 8234 16205 8268
rect 16147 8228 16205 8234
rect 16336 8225 16342 8277
rect 16394 8265 16400 8277
rect 16915 8268 16973 8274
rect 16915 8265 16927 8268
rect 16394 8237 16927 8265
rect 16394 8225 16400 8237
rect 16915 8234 16927 8237
rect 16961 8234 16973 8268
rect 17266 8265 17294 8311
rect 23536 8299 23542 8311
rect 23594 8299 23600 8351
rect 43186 8339 43214 8459
rect 48610 8413 48638 8521
rect 48883 8416 48941 8422
rect 48883 8413 48895 8416
rect 48610 8385 48895 8413
rect 48883 8382 48895 8385
rect 48929 8382 48941 8416
rect 52162 8413 52190 8524
rect 52912 8521 52918 8533
rect 52970 8521 52976 8573
rect 52435 8416 52493 8422
rect 52435 8413 52447 8416
rect 52162 8385 52447 8413
rect 48883 8376 48941 8382
rect 52435 8382 52447 8385
rect 52481 8413 52493 8416
rect 52723 8416 52781 8422
rect 52723 8413 52735 8416
rect 52481 8385 52735 8413
rect 52481 8382 52493 8385
rect 52435 8376 52493 8382
rect 52723 8382 52735 8385
rect 52769 8382 52781 8416
rect 52930 8413 52958 8521
rect 53203 8416 53261 8422
rect 53203 8413 53215 8416
rect 52930 8385 53215 8413
rect 52723 8376 52781 8382
rect 53203 8382 53215 8385
rect 53249 8382 53261 8416
rect 53203 8376 53261 8382
rect 49747 8342 49805 8348
rect 49747 8339 49759 8342
rect 43186 8311 49759 8339
rect 49747 8308 49759 8311
rect 49793 8308 49805 8342
rect 49747 8302 49805 8308
rect 49840 8299 49846 8351
rect 49898 8339 49904 8351
rect 54067 8342 54125 8348
rect 54067 8339 54079 8342
rect 49898 8311 54079 8339
rect 49898 8299 49904 8311
rect 54067 8308 54079 8311
rect 54113 8308 54125 8342
rect 54067 8302 54125 8308
rect 55219 8342 55277 8348
rect 55219 8308 55231 8342
rect 55265 8308 55277 8342
rect 55219 8302 55277 8308
rect 55987 8342 56045 8348
rect 55987 8308 55999 8342
rect 56033 8308 56045 8342
rect 55987 8302 56045 8308
rect 16915 8228 16973 8234
rect 17026 8237 17294 8265
rect 4816 8191 4822 8203
rect 4450 8163 4822 8191
rect 2282 8151 2288 8163
rect 4816 8151 4822 8163
rect 4874 8151 4880 8203
rect 5299 8194 5357 8200
rect 5299 8160 5311 8194
rect 5345 8191 5357 8194
rect 13744 8191 13750 8203
rect 5345 8163 13750 8191
rect 5345 8160 5357 8163
rect 5299 8154 5357 8160
rect 13744 8151 13750 8163
rect 13802 8151 13808 8203
rect 8080 8077 8086 8129
rect 8138 8117 8144 8129
rect 9808 8117 9814 8129
rect 8138 8089 9814 8117
rect 8138 8077 8144 8089
rect 9808 8077 9814 8089
rect 9866 8077 9872 8129
rect 10291 8120 10349 8126
rect 10291 8086 10303 8120
rect 10337 8117 10349 8120
rect 10576 8117 10582 8129
rect 10337 8089 10582 8117
rect 10337 8086 10349 8089
rect 10291 8080 10349 8086
rect 10576 8077 10582 8089
rect 10634 8117 10640 8129
rect 17026 8117 17054 8237
rect 48016 8225 48022 8277
rect 48074 8265 48080 8277
rect 48115 8268 48173 8274
rect 48115 8265 48127 8268
rect 48074 8237 48127 8265
rect 48074 8225 48080 8237
rect 48115 8234 48127 8237
rect 48161 8234 48173 8268
rect 48115 8228 48173 8234
rect 48211 8268 48269 8274
rect 48211 8234 48223 8268
rect 48257 8265 48269 8268
rect 48880 8265 48886 8277
rect 48257 8237 48886 8265
rect 48257 8234 48269 8237
rect 48211 8228 48269 8234
rect 48880 8225 48886 8237
rect 48938 8225 48944 8277
rect 48979 8268 49037 8274
rect 48979 8234 48991 8268
rect 49025 8234 49037 8268
rect 48979 8228 49037 8234
rect 17104 8151 17110 8203
rect 17162 8191 17168 8203
rect 17162 8163 47678 8191
rect 17162 8151 17168 8163
rect 10634 8089 17054 8117
rect 10634 8077 10640 8089
rect 28048 8077 28054 8129
rect 28106 8117 28112 8129
rect 33520 8117 33526 8129
rect 28106 8089 33526 8117
rect 28106 8077 28112 8089
rect 33520 8077 33526 8089
rect 33578 8077 33584 8129
rect 44368 8077 44374 8129
rect 44426 8117 44432 8129
rect 45523 8120 45581 8126
rect 45523 8117 45535 8120
rect 44426 8089 45535 8117
rect 44426 8077 44432 8089
rect 45523 8086 45535 8089
rect 45569 8086 45581 8120
rect 47650 8117 47678 8163
rect 48688 8151 48694 8203
rect 48746 8191 48752 8203
rect 48994 8191 49022 8228
rect 49456 8225 49462 8277
rect 49514 8265 49520 8277
rect 49651 8268 49709 8274
rect 49651 8265 49663 8268
rect 49514 8237 49663 8265
rect 49514 8225 49520 8237
rect 49651 8234 49663 8237
rect 49697 8234 49709 8268
rect 49651 8228 49709 8234
rect 52531 8268 52589 8274
rect 52531 8234 52543 8268
rect 52577 8234 52589 8268
rect 52531 8228 52589 8234
rect 52144 8191 52150 8203
rect 48746 8163 49022 8191
rect 49090 8163 52150 8191
rect 48746 8151 48752 8163
rect 49090 8117 49118 8163
rect 52144 8151 52150 8163
rect 52202 8151 52208 8203
rect 52546 8191 52574 8228
rect 53104 8225 53110 8277
rect 53162 8265 53168 8277
rect 53299 8268 53357 8274
rect 53299 8265 53311 8268
rect 53162 8237 53311 8265
rect 53162 8225 53168 8237
rect 53299 8234 53311 8237
rect 53345 8234 53357 8268
rect 53299 8228 53357 8234
rect 53488 8225 53494 8277
rect 53546 8265 53552 8277
rect 53971 8268 54029 8274
rect 53971 8265 53983 8268
rect 53546 8237 53983 8265
rect 53546 8225 53552 8237
rect 53971 8234 53983 8237
rect 54017 8234 54029 8268
rect 53971 8228 54029 8234
rect 55234 8191 55262 8302
rect 56002 8265 56030 8302
rect 56944 8299 56950 8351
rect 57002 8339 57008 8351
rect 57139 8342 57197 8348
rect 57139 8339 57151 8342
rect 57002 8311 57151 8339
rect 57002 8299 57008 8311
rect 57139 8308 57151 8311
rect 57185 8308 57197 8342
rect 57139 8302 57197 8308
rect 58384 8265 58390 8277
rect 56002 8237 58390 8265
rect 58384 8225 58390 8237
rect 58442 8225 58448 8277
rect 59824 8191 59830 8203
rect 52546 8163 53294 8191
rect 55234 8163 59830 8191
rect 47650 8089 49118 8117
rect 50515 8120 50573 8126
rect 45523 8080 45581 8086
rect 50515 8086 50527 8120
rect 50561 8117 50573 8120
rect 50800 8117 50806 8129
rect 50561 8089 50806 8117
rect 50561 8086 50573 8089
rect 50515 8080 50573 8086
rect 50800 8077 50806 8089
rect 50858 8077 50864 8129
rect 53266 8117 53294 8163
rect 59824 8151 59830 8163
rect 59882 8151 59888 8203
rect 58960 8117 58966 8129
rect 53266 8089 58966 8117
rect 58960 8077 58966 8089
rect 59018 8077 59024 8129
rect 1152 8018 58848 8040
rect 1152 7966 4294 8018
rect 4346 7966 4358 8018
rect 4410 7966 4422 8018
rect 4474 7966 4486 8018
rect 4538 7966 35014 8018
rect 35066 7966 35078 8018
rect 35130 7966 35142 8018
rect 35194 7966 35206 8018
rect 35258 7966 58848 8018
rect 1152 7944 58848 7966
rect 2128 7895 2134 7907
rect 2089 7867 2134 7895
rect 2128 7855 2134 7867
rect 2186 7855 2192 7907
rect 3664 7895 3670 7907
rect 3625 7867 3670 7895
rect 3664 7855 3670 7867
rect 3722 7895 3728 7907
rect 7600 7895 7606 7907
rect 3722 7867 4094 7895
rect 7561 7867 7606 7895
rect 3722 7855 3728 7867
rect 2146 7747 2174 7855
rect 4066 7756 4094 7867
rect 7600 7855 7606 7867
rect 7658 7855 7664 7907
rect 9040 7895 9046 7907
rect 7714 7867 8126 7895
rect 9001 7867 9046 7895
rect 2515 7750 2573 7756
rect 2515 7747 2527 7750
rect 2146 7719 2527 7747
rect 2515 7716 2527 7719
rect 2561 7716 2573 7750
rect 2515 7710 2573 7716
rect 4051 7750 4109 7756
rect 4051 7716 4063 7750
rect 4097 7716 4109 7750
rect 4051 7710 4109 7716
rect 4819 7750 4877 7756
rect 4819 7716 4831 7750
rect 4865 7747 4877 7750
rect 5680 7747 5686 7759
rect 4865 7719 5686 7747
rect 4865 7716 4877 7719
rect 4819 7710 4877 7716
rect 5680 7707 5686 7719
rect 5738 7707 5744 7759
rect 1456 7633 1462 7685
rect 1514 7673 1520 7685
rect 1555 7676 1613 7682
rect 1555 7673 1567 7676
rect 1514 7645 1567 7673
rect 1514 7633 1520 7645
rect 1555 7642 1567 7645
rect 1601 7642 1613 7676
rect 1555 7636 1613 7642
rect 3283 7676 3341 7682
rect 3283 7642 3295 7676
rect 3329 7673 3341 7676
rect 7714 7673 7742 7867
rect 8098 7821 8126 7867
rect 9040 7855 9046 7867
rect 9098 7855 9104 7907
rect 28048 7895 28054 7907
rect 9538 7867 28054 7895
rect 9538 7821 9566 7867
rect 28048 7855 28054 7867
rect 28106 7855 28112 7907
rect 29008 7895 29014 7907
rect 28969 7867 29014 7895
rect 29008 7855 29014 7867
rect 29066 7895 29072 7907
rect 36496 7895 36502 7907
rect 29066 7867 29342 7895
rect 36457 7867 36502 7895
rect 29066 7855 29072 7867
rect 8098 7793 9566 7821
rect 9616 7781 9622 7833
rect 9674 7821 9680 7833
rect 10675 7824 10733 7830
rect 9674 7793 10622 7821
rect 9674 7781 9680 7793
rect 8080 7747 8086 7759
rect 7968 7719 8086 7747
rect 8080 7707 8086 7719
rect 8138 7707 8144 7759
rect 8368 7747 8374 7759
rect 8256 7719 8374 7747
rect 8368 7707 8374 7719
rect 8426 7707 8432 7759
rect 9040 7707 9046 7759
rect 9098 7747 9104 7759
rect 9427 7750 9485 7756
rect 9427 7747 9439 7750
rect 9098 7719 9439 7747
rect 9098 7707 9104 7719
rect 9427 7716 9439 7719
rect 9473 7716 9485 7750
rect 10099 7750 10157 7756
rect 10099 7747 10111 7750
rect 9427 7710 9485 7716
rect 9538 7719 10111 7747
rect 3329 7645 7742 7673
rect 3329 7642 3341 7645
rect 3283 7636 3341 7642
rect 9136 7633 9142 7685
rect 9194 7673 9200 7685
rect 9538 7673 9566 7719
rect 10099 7716 10111 7719
rect 10145 7716 10157 7750
rect 10099 7710 10157 7716
rect 10192 7673 10198 7685
rect 9194 7645 9566 7673
rect 10153 7645 10198 7673
rect 9194 7633 9200 7645
rect 10192 7633 10198 7645
rect 10250 7633 10256 7685
rect 10594 7673 10622 7793
rect 10675 7790 10687 7824
rect 10721 7821 10733 7824
rect 10721 7793 11006 7821
rect 10721 7790 10733 7793
rect 10675 7784 10733 7790
rect 10978 7756 11006 7793
rect 13744 7781 13750 7833
rect 13802 7821 13808 7833
rect 25072 7821 25078 7833
rect 13802 7793 13982 7821
rect 25033 7793 25078 7821
rect 13802 7781 13808 7793
rect 10963 7750 11021 7756
rect 10963 7716 10975 7750
rect 11009 7747 11021 7750
rect 12592 7747 12598 7759
rect 11009 7719 12598 7747
rect 11009 7716 11021 7719
rect 10963 7710 11021 7716
rect 12592 7707 12598 7719
rect 12650 7707 12656 7759
rect 12688 7707 12694 7759
rect 12746 7747 12752 7759
rect 13954 7756 13982 7793
rect 25072 7781 25078 7793
rect 25130 7821 25136 7833
rect 25130 7793 25502 7821
rect 25130 7781 25136 7793
rect 13843 7750 13901 7756
rect 13843 7747 13855 7750
rect 12746 7719 13855 7747
rect 12746 7707 12752 7719
rect 13843 7716 13855 7719
rect 13889 7716 13901 7750
rect 13843 7710 13901 7716
rect 13939 7750 13997 7756
rect 13939 7716 13951 7750
rect 13985 7716 13997 7750
rect 13939 7710 13997 7716
rect 15571 7750 15629 7756
rect 15571 7716 15583 7750
rect 15617 7747 15629 7750
rect 15856 7747 15862 7759
rect 15617 7719 15862 7747
rect 15617 7716 15629 7719
rect 15571 7710 15629 7716
rect 15856 7707 15862 7719
rect 15914 7707 15920 7759
rect 20944 7747 20950 7759
rect 20905 7719 20950 7747
rect 20944 7707 20950 7719
rect 21002 7707 21008 7759
rect 23635 7750 23693 7756
rect 23635 7716 23647 7750
rect 23681 7747 23693 7750
rect 23920 7747 23926 7759
rect 23681 7719 23926 7747
rect 23681 7716 23693 7719
rect 23635 7710 23693 7716
rect 23920 7707 23926 7719
rect 23978 7707 23984 7759
rect 24688 7747 24694 7759
rect 24649 7719 24694 7747
rect 24688 7707 24694 7719
rect 24746 7707 24752 7759
rect 25474 7756 25502 7793
rect 27760 7781 27766 7833
rect 27818 7821 27824 7833
rect 27955 7824 28013 7830
rect 27955 7821 27967 7824
rect 27818 7793 27967 7821
rect 27818 7781 27824 7793
rect 27955 7790 27967 7793
rect 28001 7821 28013 7824
rect 28001 7793 28286 7821
rect 28001 7790 28013 7793
rect 27955 7784 28013 7790
rect 25459 7750 25517 7756
rect 25459 7716 25471 7750
rect 25505 7716 25517 7750
rect 25459 7710 25517 7716
rect 25939 7750 25997 7756
rect 25939 7716 25951 7750
rect 25985 7747 25997 7750
rect 26128 7747 26134 7759
rect 25985 7719 26134 7747
rect 25985 7716 25997 7719
rect 25939 7710 25997 7716
rect 26128 7707 26134 7719
rect 26186 7707 26192 7759
rect 26992 7747 26998 7759
rect 26953 7719 26998 7747
rect 26992 7707 26998 7719
rect 27050 7707 27056 7759
rect 28258 7756 28286 7793
rect 29314 7756 29342 7867
rect 36496 7855 36502 7867
rect 36554 7895 36560 7907
rect 41488 7895 41494 7907
rect 36554 7867 36830 7895
rect 41449 7867 41494 7895
rect 36554 7855 36560 7867
rect 28243 7750 28301 7756
rect 28243 7716 28255 7750
rect 28289 7716 28301 7750
rect 28243 7710 28301 7716
rect 29299 7750 29357 7756
rect 29299 7716 29311 7750
rect 29345 7716 29357 7750
rect 29299 7710 29357 7716
rect 29875 7750 29933 7756
rect 29875 7716 29887 7750
rect 29921 7747 29933 7750
rect 30160 7747 30166 7759
rect 29921 7719 30166 7747
rect 29921 7716 29933 7719
rect 29875 7710 29933 7716
rect 30160 7707 30166 7719
rect 30218 7707 30224 7759
rect 33328 7747 33334 7759
rect 30274 7719 33334 7747
rect 12304 7673 12310 7685
rect 10594 7645 12310 7673
rect 12304 7633 12310 7645
rect 12362 7633 12368 7685
rect 13171 7676 13229 7682
rect 13171 7642 13183 7676
rect 13217 7673 13229 7676
rect 28915 7676 28973 7682
rect 28915 7673 28927 7676
rect 13217 7645 28927 7673
rect 13217 7642 13229 7645
rect 13171 7636 13229 7642
rect 28915 7642 28927 7645
rect 28961 7642 28973 7676
rect 28915 7636 28973 7642
rect 5299 7602 5357 7608
rect 5299 7568 5311 7602
rect 5345 7599 5357 7602
rect 5584 7599 5590 7611
rect 5345 7571 5590 7599
rect 5345 7568 5357 7571
rect 5299 7562 5357 7568
rect 5584 7559 5590 7571
rect 5642 7559 5648 7611
rect 11248 7599 11254 7611
rect 9058 7571 11254 7599
rect 9058 7525 9086 7571
rect 11248 7559 11254 7571
rect 11306 7559 11312 7611
rect 12115 7602 12173 7608
rect 12115 7568 12127 7602
rect 12161 7599 12173 7602
rect 12403 7602 12461 7608
rect 12403 7599 12415 7602
rect 12161 7571 12415 7599
rect 12161 7568 12173 7571
rect 12115 7562 12173 7568
rect 12403 7568 12415 7571
rect 12449 7568 12461 7602
rect 12403 7562 12461 7568
rect 8544 7497 9086 7525
rect 12418 7525 12446 7562
rect 12496 7559 12502 7611
rect 12554 7599 12560 7611
rect 17104 7599 17110 7611
rect 12554 7571 17110 7599
rect 12554 7559 12560 7571
rect 17104 7559 17110 7571
rect 17162 7559 17168 7611
rect 30274 7599 30302 7719
rect 33328 7707 33334 7719
rect 33386 7707 33392 7759
rect 33523 7750 33581 7756
rect 33523 7716 33535 7750
rect 33569 7747 33581 7750
rect 33715 7750 33773 7756
rect 33715 7747 33727 7750
rect 33569 7719 33727 7747
rect 33569 7716 33581 7719
rect 33523 7710 33581 7716
rect 33715 7716 33727 7719
rect 33761 7747 33773 7750
rect 33808 7747 33814 7759
rect 33761 7719 33814 7747
rect 33761 7716 33773 7719
rect 33715 7710 33773 7716
rect 33808 7707 33814 7719
rect 33866 7707 33872 7759
rect 34291 7750 34349 7756
rect 34291 7716 34303 7750
rect 34337 7747 34349 7750
rect 34576 7747 34582 7759
rect 34337 7719 34582 7747
rect 34337 7716 34349 7719
rect 34291 7710 34349 7716
rect 34576 7707 34582 7719
rect 34634 7707 34640 7759
rect 35344 7747 35350 7759
rect 35305 7719 35350 7747
rect 35344 7707 35350 7719
rect 35402 7707 35408 7759
rect 36112 7747 36118 7759
rect 36073 7719 36118 7747
rect 36112 7707 36118 7719
rect 36170 7707 36176 7759
rect 36802 7756 36830 7867
rect 41488 7855 41494 7867
rect 41546 7855 41552 7907
rect 42256 7895 42262 7907
rect 42217 7867 42262 7895
rect 42256 7855 42262 7867
rect 42314 7895 42320 7907
rect 42314 7867 42686 7895
rect 42314 7855 42320 7867
rect 38800 7821 38806 7833
rect 37426 7793 38806 7821
rect 36787 7750 36845 7756
rect 36787 7716 36799 7750
rect 36833 7716 36845 7750
rect 36787 7710 36845 7716
rect 31219 7676 31277 7682
rect 31219 7642 31231 7676
rect 31265 7673 31277 7676
rect 37426 7673 37454 7793
rect 38800 7781 38806 7793
rect 38858 7781 38864 7833
rect 39682 7793 41150 7821
rect 38515 7750 38573 7756
rect 38515 7716 38527 7750
rect 38561 7747 38573 7750
rect 38704 7747 38710 7759
rect 38561 7719 38710 7747
rect 38561 7716 38573 7719
rect 38515 7710 38573 7716
rect 38704 7707 38710 7719
rect 38762 7707 38768 7759
rect 39283 7750 39341 7756
rect 39283 7716 39295 7750
rect 39329 7747 39341 7750
rect 39472 7747 39478 7759
rect 39329 7719 39478 7747
rect 39329 7716 39341 7719
rect 39283 7710 39341 7716
rect 39472 7707 39478 7719
rect 39530 7707 39536 7759
rect 39571 7750 39629 7756
rect 39571 7716 39583 7750
rect 39617 7716 39629 7750
rect 39571 7710 39629 7716
rect 31265 7645 37454 7673
rect 31265 7642 31277 7645
rect 31219 7636 31277 7642
rect 38800 7633 38806 7685
rect 38858 7673 38864 7685
rect 39586 7673 39614 7710
rect 38858 7645 39614 7673
rect 38858 7633 38864 7645
rect 27970 7571 30302 7599
rect 31987 7602 32045 7608
rect 27970 7525 27998 7571
rect 31987 7568 31999 7602
rect 32033 7599 32045 7602
rect 34480 7599 34486 7611
rect 32033 7571 34486 7599
rect 32033 7568 32045 7571
rect 31987 7562 32045 7568
rect 34480 7559 34486 7571
rect 34538 7559 34544 7611
rect 39682 7599 39710 7793
rect 40336 7747 40342 7759
rect 40297 7719 40342 7747
rect 40336 7707 40342 7719
rect 40394 7707 40400 7759
rect 41011 7750 41069 7756
rect 41011 7716 41023 7750
rect 41057 7716 41069 7750
rect 41011 7710 41069 7716
rect 40240 7633 40246 7685
rect 40298 7673 40304 7685
rect 41026 7673 41054 7710
rect 40298 7645 41054 7673
rect 41122 7673 41150 7793
rect 41392 7707 41398 7759
rect 41450 7747 41456 7759
rect 42658 7756 42686 7867
rect 45040 7855 45046 7907
rect 45098 7895 45104 7907
rect 45235 7898 45293 7904
rect 45235 7895 45247 7898
rect 45098 7867 45247 7895
rect 45098 7855 45104 7867
rect 45235 7864 45247 7867
rect 45281 7895 45293 7898
rect 47536 7895 47542 7907
rect 45281 7867 45566 7895
rect 47497 7867 47542 7895
rect 45281 7864 45293 7867
rect 45235 7858 45293 7864
rect 41875 7750 41933 7756
rect 41875 7747 41887 7750
rect 41450 7719 41887 7747
rect 41450 7707 41456 7719
rect 41875 7716 41887 7719
rect 41921 7716 41933 7750
rect 41875 7710 41933 7716
rect 42643 7750 42701 7756
rect 42643 7716 42655 7750
rect 42689 7716 42701 7750
rect 42643 7710 42701 7716
rect 44752 7707 44758 7759
rect 44810 7747 44816 7759
rect 45538 7756 45566 7867
rect 47536 7855 47542 7867
rect 47594 7895 47600 7907
rect 48115 7898 48173 7904
rect 48115 7895 48127 7898
rect 47594 7867 48127 7895
rect 47594 7855 47600 7867
rect 44851 7750 44909 7756
rect 44851 7747 44863 7750
rect 44810 7719 44863 7747
rect 44810 7707 44816 7719
rect 44851 7716 44863 7719
rect 44897 7716 44909 7750
rect 44851 7710 44909 7716
rect 45523 7750 45581 7756
rect 45523 7716 45535 7750
rect 45569 7716 45581 7750
rect 45523 7710 45581 7716
rect 46288 7707 46294 7759
rect 46346 7747 46352 7759
rect 47842 7756 47870 7867
rect 48115 7864 48127 7867
rect 48161 7864 48173 7898
rect 48115 7858 48173 7864
rect 49552 7855 49558 7907
rect 49610 7895 49616 7907
rect 50707 7898 50765 7904
rect 50707 7895 50719 7898
rect 49610 7867 50719 7895
rect 49610 7855 49616 7867
rect 50707 7864 50719 7867
rect 50753 7895 50765 7898
rect 50753 7867 51038 7895
rect 50753 7864 50765 7867
rect 50707 7858 50765 7864
rect 46387 7750 46445 7756
rect 46387 7747 46399 7750
rect 46346 7719 46399 7747
rect 46346 7707 46352 7719
rect 46387 7716 46399 7719
rect 46433 7716 46445 7750
rect 46387 7710 46445 7716
rect 47827 7750 47885 7756
rect 47827 7716 47839 7750
rect 47873 7716 47885 7750
rect 49360 7747 49366 7759
rect 49321 7719 49366 7747
rect 47827 7710 47885 7716
rect 49360 7707 49366 7719
rect 49418 7707 49424 7759
rect 50032 7707 50038 7759
rect 50090 7747 50096 7759
rect 51010 7756 51038 7867
rect 59344 7821 59350 7833
rect 53266 7793 59350 7821
rect 50131 7750 50189 7756
rect 50131 7747 50143 7750
rect 50090 7719 50143 7747
rect 50090 7707 50096 7719
rect 50131 7716 50143 7719
rect 50177 7716 50189 7750
rect 50131 7710 50189 7716
rect 50995 7750 51053 7756
rect 50995 7716 51007 7750
rect 51041 7716 51053 7750
rect 50995 7710 51053 7716
rect 51091 7750 51149 7756
rect 51091 7716 51103 7750
rect 51137 7747 51149 7750
rect 53266 7747 53294 7793
rect 59344 7781 59350 7793
rect 59402 7781 59408 7833
rect 51137 7719 53294 7747
rect 53395 7750 53453 7756
rect 51137 7716 51149 7719
rect 51091 7710 51149 7716
rect 53395 7716 53407 7750
rect 53441 7747 53453 7750
rect 53584 7747 53590 7759
rect 53441 7719 53590 7747
rect 53441 7716 53453 7719
rect 53395 7710 53453 7716
rect 53584 7707 53590 7719
rect 53642 7707 53648 7759
rect 44272 7673 44278 7685
rect 41122 7645 44278 7673
rect 40298 7633 40304 7645
rect 44272 7633 44278 7645
rect 44330 7633 44336 7685
rect 45424 7633 45430 7685
rect 45482 7673 45488 7685
rect 46771 7676 46829 7682
rect 46771 7673 46783 7676
rect 45482 7645 46783 7673
rect 45482 7633 45488 7645
rect 46771 7642 46783 7645
rect 46817 7673 46829 7676
rect 47059 7676 47117 7682
rect 47059 7673 47071 7676
rect 46817 7645 47071 7673
rect 46817 7642 46829 7645
rect 46771 7636 46829 7642
rect 47059 7642 47071 7645
rect 47105 7642 47117 7676
rect 47059 7636 47117 7642
rect 49744 7633 49750 7685
rect 49802 7673 49808 7685
rect 51475 7676 51533 7682
rect 51475 7673 51487 7676
rect 49802 7645 51487 7673
rect 49802 7633 49808 7645
rect 51475 7642 51487 7645
rect 51521 7673 51533 7676
rect 51763 7676 51821 7682
rect 51763 7673 51775 7676
rect 51521 7645 51775 7673
rect 51521 7642 51533 7645
rect 51475 7636 51533 7642
rect 51763 7642 51775 7645
rect 51809 7642 51821 7676
rect 51763 7636 51821 7642
rect 55123 7676 55181 7682
rect 55123 7642 55135 7676
rect 55169 7642 55181 7676
rect 55792 7673 55798 7685
rect 55753 7645 55798 7673
rect 55123 7636 55181 7642
rect 37426 7571 39710 7599
rect 12418 7497 27998 7525
rect 28915 7528 28973 7534
rect 28915 7494 28927 7528
rect 28961 7525 28973 7528
rect 37426 7525 37454 7571
rect 39952 7559 39958 7611
rect 40010 7599 40016 7611
rect 41107 7602 41165 7608
rect 41107 7599 41119 7602
rect 40010 7571 41119 7599
rect 40010 7559 40016 7571
rect 41107 7568 41119 7571
rect 41153 7568 41165 7602
rect 41107 7562 41165 7568
rect 41488 7559 41494 7611
rect 41546 7599 41552 7611
rect 41779 7602 41837 7608
rect 41779 7599 41791 7602
rect 41546 7571 41791 7599
rect 41546 7559 41552 7571
rect 41779 7568 41791 7571
rect 41825 7568 41837 7602
rect 41779 7562 41837 7568
rect 43795 7602 43853 7608
rect 43795 7568 43807 7602
rect 43841 7599 43853 7602
rect 44083 7602 44141 7608
rect 44083 7599 44095 7602
rect 43841 7571 44095 7599
rect 43841 7568 43853 7571
rect 43795 7562 43853 7568
rect 44083 7568 44095 7571
rect 44129 7599 44141 7602
rect 45328 7599 45334 7611
rect 44129 7571 45334 7599
rect 44129 7568 44141 7571
rect 44083 7562 44141 7568
rect 45328 7559 45334 7571
rect 45386 7559 45392 7611
rect 52627 7602 52685 7608
rect 52627 7568 52639 7602
rect 52673 7599 52685 7602
rect 52816 7599 52822 7611
rect 52673 7571 52822 7599
rect 52673 7568 52685 7571
rect 52627 7562 52685 7568
rect 52816 7559 52822 7571
rect 52874 7559 52880 7611
rect 55138 7599 55166 7636
rect 55792 7633 55798 7645
rect 55850 7633 55856 7685
rect 56176 7633 56182 7685
rect 56234 7673 56240 7685
rect 56563 7676 56621 7682
rect 56563 7673 56575 7676
rect 56234 7645 56575 7673
rect 56234 7633 56240 7645
rect 56563 7642 56575 7645
rect 56609 7642 56621 7676
rect 56563 7636 56621 7642
rect 56656 7633 56662 7685
rect 56714 7673 56720 7685
rect 57331 7676 57389 7682
rect 57331 7673 57343 7676
rect 56714 7645 57343 7673
rect 56714 7633 56720 7645
rect 57331 7642 57343 7645
rect 57377 7642 57389 7676
rect 57331 7636 57389 7642
rect 58768 7599 58774 7611
rect 55138 7571 58774 7599
rect 58768 7559 58774 7571
rect 58826 7559 58832 7611
rect 28961 7497 37454 7525
rect 28961 7494 28973 7497
rect 28915 7488 28973 7494
rect 39472 7485 39478 7537
rect 39530 7525 39536 7537
rect 39530 7497 40286 7525
rect 39530 7485 39536 7497
rect 2320 7411 2326 7463
rect 2378 7451 2384 7463
rect 2419 7454 2477 7460
rect 2419 7451 2431 7454
rect 2378 7423 2431 7451
rect 2378 7411 2384 7423
rect 2419 7420 2431 7423
rect 2465 7420 2477 7454
rect 2419 7414 2477 7420
rect 2992 7411 2998 7463
rect 3050 7451 3056 7463
rect 3187 7454 3245 7460
rect 3187 7451 3199 7454
rect 3050 7423 3199 7451
rect 3050 7411 3056 7423
rect 3187 7420 3199 7423
rect 3233 7420 3245 7454
rect 3952 7451 3958 7463
rect 3913 7423 3958 7451
rect 3187 7414 3245 7420
rect 3952 7411 3958 7423
rect 4010 7411 4016 7463
rect 4048 7411 4054 7463
rect 4106 7451 4112 7463
rect 4723 7454 4781 7460
rect 4723 7451 4735 7454
rect 4106 7423 4735 7451
rect 4106 7411 4112 7423
rect 4723 7420 4735 7423
rect 4769 7420 4781 7454
rect 4723 7414 4781 7420
rect 5296 7411 5302 7463
rect 5354 7451 5360 7463
rect 5491 7454 5549 7460
rect 5491 7451 5503 7454
rect 5354 7423 5503 7451
rect 5354 7411 5360 7423
rect 5491 7420 5503 7423
rect 5537 7420 5549 7454
rect 5491 7414 5549 7420
rect 8368 7411 8374 7463
rect 8426 7411 8432 7463
rect 8752 7411 8758 7463
rect 8810 7451 8816 7463
rect 9331 7454 9389 7460
rect 9331 7451 9343 7454
rect 8810 7423 9343 7451
rect 8810 7411 8816 7423
rect 9331 7420 9343 7423
rect 9377 7420 9389 7454
rect 9331 7414 9389 7420
rect 9904 7411 9910 7463
rect 9962 7451 9968 7463
rect 10867 7454 10925 7460
rect 10867 7451 10879 7454
rect 9962 7423 10879 7451
rect 9962 7411 9968 7423
rect 10867 7420 10879 7423
rect 10913 7420 10925 7454
rect 10867 7414 10925 7420
rect 10960 7411 10966 7463
rect 11018 7451 11024 7463
rect 12307 7454 12365 7460
rect 12307 7451 12319 7454
rect 11018 7423 12319 7451
rect 11018 7411 11024 7423
rect 12307 7420 12319 7423
rect 12353 7420 12365 7454
rect 12307 7414 12365 7420
rect 12400 7411 12406 7463
rect 12458 7451 12464 7463
rect 13075 7454 13133 7460
rect 13075 7451 13087 7454
rect 12458 7423 13087 7451
rect 12458 7411 12464 7423
rect 13075 7420 13087 7423
rect 13121 7420 13133 7454
rect 13075 7414 13133 7420
rect 15664 7411 15670 7463
rect 15722 7451 15728 7463
rect 15763 7454 15821 7460
rect 15763 7451 15775 7454
rect 15722 7423 15775 7451
rect 15722 7411 15728 7423
rect 15763 7420 15775 7423
rect 15809 7420 15821 7454
rect 15763 7414 15821 7420
rect 20752 7411 20758 7463
rect 20810 7451 20816 7463
rect 20851 7454 20909 7460
rect 20851 7451 20863 7454
rect 20810 7423 20863 7451
rect 20810 7411 20816 7423
rect 20851 7420 20863 7423
rect 20897 7420 20909 7454
rect 23824 7451 23830 7463
rect 23785 7423 23830 7451
rect 20851 7414 20909 7420
rect 23824 7411 23830 7423
rect 23882 7411 23888 7463
rect 24208 7411 24214 7463
rect 24266 7451 24272 7463
rect 24595 7454 24653 7460
rect 24595 7451 24607 7454
rect 24266 7423 24607 7451
rect 24266 7411 24272 7423
rect 24595 7420 24607 7423
rect 24641 7420 24653 7454
rect 24595 7414 24653 7420
rect 24784 7411 24790 7463
rect 24842 7451 24848 7463
rect 25363 7454 25421 7460
rect 25363 7451 25375 7454
rect 24842 7423 25375 7451
rect 24842 7411 24848 7423
rect 25363 7420 25375 7423
rect 25409 7420 25421 7454
rect 25363 7414 25421 7420
rect 25552 7411 25558 7463
rect 25610 7451 25616 7463
rect 26227 7454 26285 7460
rect 26227 7451 26239 7454
rect 25610 7423 26239 7451
rect 25610 7411 25616 7423
rect 26227 7420 26239 7423
rect 26273 7420 26285 7454
rect 26227 7414 26285 7420
rect 26704 7411 26710 7463
rect 26762 7451 26768 7463
rect 26899 7454 26957 7460
rect 26899 7451 26911 7454
rect 26762 7423 26911 7451
rect 26762 7411 26768 7423
rect 26899 7420 26911 7423
rect 26945 7420 26957 7454
rect 26899 7414 26957 7420
rect 28144 7411 28150 7463
rect 28202 7451 28208 7463
rect 28339 7454 28397 7460
rect 28339 7451 28351 7454
rect 28202 7423 28351 7451
rect 28202 7411 28208 7423
rect 28339 7420 28351 7423
rect 28385 7420 28397 7454
rect 28339 7414 28397 7420
rect 29200 7411 29206 7463
rect 29258 7451 29264 7463
rect 29395 7454 29453 7460
rect 29395 7451 29407 7454
rect 29258 7423 29407 7451
rect 29258 7411 29264 7423
rect 29395 7420 29407 7423
rect 29441 7420 29453 7454
rect 29395 7414 29453 7420
rect 29584 7411 29590 7463
rect 29642 7451 29648 7463
rect 30067 7454 30125 7460
rect 30067 7451 30079 7454
rect 29642 7423 30079 7451
rect 29642 7411 29648 7423
rect 30067 7420 30079 7423
rect 30113 7420 30125 7454
rect 31120 7451 31126 7463
rect 31081 7423 31126 7451
rect 30067 7414 30125 7420
rect 31120 7411 31126 7423
rect 31178 7411 31184 7463
rect 33616 7411 33622 7463
rect 33674 7451 33680 7463
rect 33811 7454 33869 7460
rect 33811 7451 33823 7454
rect 33674 7423 33823 7451
rect 33674 7411 33680 7423
rect 33811 7420 33823 7423
rect 33857 7420 33869 7454
rect 33811 7414 33869 7420
rect 34384 7411 34390 7463
rect 34442 7451 34448 7463
rect 34483 7454 34541 7460
rect 34483 7451 34495 7454
rect 34442 7423 34495 7451
rect 34442 7411 34448 7423
rect 34483 7420 34495 7423
rect 34529 7420 34541 7454
rect 34483 7414 34541 7420
rect 34672 7411 34678 7463
rect 34730 7451 34736 7463
rect 35251 7454 35309 7460
rect 35251 7451 35263 7454
rect 34730 7423 35263 7451
rect 34730 7411 34736 7423
rect 35251 7420 35263 7423
rect 35297 7420 35309 7454
rect 36016 7451 36022 7463
rect 35977 7423 36022 7451
rect 35251 7414 35309 7420
rect 36016 7411 36022 7423
rect 36074 7411 36080 7463
rect 36592 7411 36598 7463
rect 36650 7451 36656 7463
rect 36883 7454 36941 7460
rect 36883 7451 36895 7454
rect 36650 7423 36895 7451
rect 36650 7411 36656 7423
rect 36883 7420 36895 7423
rect 36929 7420 36941 7454
rect 36883 7414 36941 7420
rect 38032 7411 38038 7463
rect 38090 7451 38096 7463
rect 40258 7460 40286 7497
rect 38803 7454 38861 7460
rect 38803 7451 38815 7454
rect 38090 7423 38815 7451
rect 38090 7411 38096 7423
rect 38803 7420 38815 7423
rect 38849 7420 38861 7454
rect 38803 7414 38861 7420
rect 40243 7454 40301 7460
rect 40243 7420 40255 7454
rect 40289 7420 40301 7454
rect 40243 7414 40301 7420
rect 42448 7411 42454 7463
rect 42506 7451 42512 7463
rect 42547 7454 42605 7460
rect 42547 7451 42559 7454
rect 42506 7423 42559 7451
rect 42506 7411 42512 7423
rect 42547 7420 42559 7423
rect 42593 7420 42605 7454
rect 42547 7414 42605 7420
rect 43888 7411 43894 7463
rect 43946 7451 43952 7463
rect 43987 7454 44045 7460
rect 43987 7451 43999 7454
rect 43946 7423 43999 7451
rect 43946 7411 43952 7423
rect 43987 7420 43999 7423
rect 44033 7420 44045 7454
rect 43987 7414 44045 7420
rect 44656 7411 44662 7463
rect 44714 7451 44720 7463
rect 44755 7454 44813 7460
rect 44755 7451 44767 7454
rect 44714 7423 44767 7451
rect 44714 7411 44720 7423
rect 44755 7420 44767 7423
rect 44801 7420 44813 7454
rect 44755 7414 44813 7420
rect 45040 7411 45046 7463
rect 45098 7451 45104 7463
rect 45619 7454 45677 7460
rect 45619 7451 45631 7454
rect 45098 7423 45631 7451
rect 45098 7411 45104 7423
rect 45619 7420 45631 7423
rect 45665 7420 45677 7454
rect 45619 7414 45677 7420
rect 45808 7411 45814 7463
rect 45866 7451 45872 7463
rect 46291 7454 46349 7460
rect 46291 7451 46303 7454
rect 45866 7423 46303 7451
rect 45866 7411 45872 7423
rect 46291 7420 46303 7423
rect 46337 7420 46349 7454
rect 46291 7414 46349 7420
rect 46576 7411 46582 7463
rect 46634 7451 46640 7463
rect 47155 7454 47213 7460
rect 47155 7451 47167 7454
rect 46634 7423 47167 7451
rect 46634 7411 46640 7423
rect 47155 7420 47167 7423
rect 47201 7420 47213 7454
rect 47155 7414 47213 7420
rect 47248 7411 47254 7463
rect 47306 7451 47312 7463
rect 47923 7454 47981 7460
rect 47923 7451 47935 7454
rect 47306 7423 47935 7451
rect 47306 7411 47312 7423
rect 47923 7420 47935 7423
rect 47969 7420 47981 7454
rect 47923 7414 47981 7420
rect 48304 7411 48310 7463
rect 48362 7451 48368 7463
rect 49267 7454 49325 7460
rect 49267 7451 49279 7454
rect 48362 7423 49279 7451
rect 48362 7411 48368 7423
rect 49267 7420 49279 7423
rect 49313 7420 49325 7454
rect 50032 7451 50038 7463
rect 49993 7423 50038 7451
rect 49267 7414 49325 7420
rect 50032 7411 50038 7423
rect 50090 7411 50096 7463
rect 51664 7411 51670 7463
rect 51722 7451 51728 7463
rect 51859 7454 51917 7460
rect 51859 7451 51871 7454
rect 51722 7423 51871 7451
rect 51722 7411 51728 7423
rect 51859 7420 51871 7423
rect 51905 7420 51917 7454
rect 51859 7414 51917 7420
rect 52336 7411 52342 7463
rect 52394 7451 52400 7463
rect 52531 7454 52589 7460
rect 52531 7451 52543 7454
rect 52394 7423 52543 7451
rect 52394 7411 52400 7423
rect 52531 7420 52543 7423
rect 52577 7420 52589 7454
rect 52531 7414 52589 7420
rect 52720 7411 52726 7463
rect 52778 7451 52784 7463
rect 53299 7454 53357 7460
rect 53299 7451 53311 7454
rect 52778 7423 53311 7451
rect 52778 7411 52784 7423
rect 53299 7420 53311 7423
rect 53345 7420 53357 7454
rect 53299 7414 53357 7420
rect 1152 7352 58848 7374
rect 1152 7300 19654 7352
rect 19706 7300 19718 7352
rect 19770 7300 19782 7352
rect 19834 7300 19846 7352
rect 19898 7300 50374 7352
rect 50426 7300 50438 7352
rect 50490 7300 50502 7352
rect 50554 7300 50566 7352
rect 50618 7300 58848 7352
rect 1152 7278 58848 7300
rect 5584 7189 5590 7241
rect 5642 7229 5648 7241
rect 12496 7229 12502 7241
rect 5642 7201 12502 7229
rect 5642 7189 5648 7201
rect 12496 7189 12502 7201
rect 12554 7189 12560 7241
rect 12784 7189 12790 7241
rect 12842 7229 12848 7241
rect 12976 7229 12982 7241
rect 12842 7201 12982 7229
rect 12842 7189 12848 7201
rect 12976 7189 12982 7201
rect 13034 7189 13040 7241
rect 13282 7201 13502 7229
rect 8848 7115 8854 7167
rect 8906 7155 8912 7167
rect 10499 7158 10557 7164
rect 10499 7155 10511 7158
rect 8906 7127 10511 7155
rect 8906 7115 8912 7127
rect 10499 7124 10511 7127
rect 10545 7124 10557 7158
rect 10499 7118 10557 7124
rect 11536 7115 11542 7167
rect 11594 7155 11600 7167
rect 13282 7155 13310 7201
rect 11594 7127 13310 7155
rect 11594 7115 11600 7127
rect 6064 7081 6070 7093
rect 6025 7053 6070 7081
rect 6064 7041 6070 7053
rect 6122 7041 6128 7093
rect 13474 7081 13502 7201
rect 17104 7189 17110 7241
rect 17162 7229 17168 7241
rect 17203 7232 17261 7238
rect 17203 7229 17215 7232
rect 17162 7201 17215 7229
rect 17162 7189 17168 7201
rect 17203 7198 17215 7201
rect 17249 7198 17261 7232
rect 17968 7229 17974 7241
rect 17929 7201 17974 7229
rect 17203 7192 17261 7198
rect 17968 7189 17974 7201
rect 18026 7189 18032 7241
rect 18640 7189 18646 7241
rect 18698 7229 18704 7241
rect 18739 7232 18797 7238
rect 18739 7229 18751 7232
rect 18698 7201 18751 7229
rect 18698 7189 18704 7201
rect 18739 7198 18751 7201
rect 18785 7198 18797 7232
rect 44563 7232 44621 7238
rect 18739 7192 18797 7198
rect 28162 7201 29534 7229
rect 17011 7158 17069 7164
rect 17011 7124 17023 7158
rect 17057 7155 17069 7158
rect 17296 7155 17302 7167
rect 17057 7127 17302 7155
rect 17057 7124 17069 7127
rect 17011 7118 17069 7124
rect 17296 7115 17302 7127
rect 17354 7115 17360 7167
rect 17890 7127 18206 7155
rect 13651 7084 13709 7090
rect 13651 7081 13663 7084
rect 6754 7053 12974 7081
rect 13474 7053 13663 7081
rect 1648 7007 1654 7019
rect 1609 6979 1654 7007
rect 1648 6967 1654 6979
rect 1706 6967 1712 7019
rect 2512 7007 2518 7019
rect 2473 6979 2518 7007
rect 2512 6967 2518 6979
rect 2570 6967 2576 7019
rect 5011 7010 5069 7016
rect 5011 6976 5023 7010
rect 5057 7007 5069 7010
rect 5299 7010 5357 7016
rect 5299 7007 5311 7010
rect 5057 6979 5311 7007
rect 5057 6976 5069 6979
rect 5011 6970 5069 6976
rect 5299 6976 5311 6979
rect 5345 7007 5357 7010
rect 6754 7007 6782 7053
rect 5345 6979 6782 7007
rect 6835 7010 6893 7016
rect 5345 6976 5357 6979
rect 5299 6970 5357 6976
rect 6835 6976 6847 7010
rect 6881 7007 6893 7010
rect 11248 7007 11254 7019
rect 6881 6979 10046 7007
rect 11209 6979 11254 7007
rect 6881 6976 6893 6979
rect 6835 6970 6893 6976
rect 4435 6936 4493 6942
rect 4435 6902 4447 6936
rect 4481 6902 4493 6936
rect 4435 6896 4493 6902
rect 4531 6936 4589 6942
rect 4531 6902 4543 6936
rect 4577 6933 4589 6936
rect 5104 6933 5110 6945
rect 4577 6905 5110 6933
rect 4577 6902 4589 6905
rect 4531 6896 4589 6902
rect 4450 6859 4478 6896
rect 5104 6893 5110 6905
rect 5162 6893 5168 6945
rect 5203 6936 5261 6942
rect 5203 6902 5215 6936
rect 5249 6902 5261 6936
rect 5203 6896 5261 6902
rect 5008 6859 5014 6871
rect 4450 6831 5014 6859
rect 5008 6819 5014 6831
rect 5066 6819 5072 6871
rect 3664 6745 3670 6797
rect 3722 6785 3728 6797
rect 5218 6785 5246 6896
rect 5872 6893 5878 6945
rect 5930 6933 5936 6945
rect 5971 6936 6029 6942
rect 5971 6933 5983 6936
rect 5930 6905 5983 6933
rect 5930 6893 5936 6905
rect 5971 6902 5983 6905
rect 6017 6902 6029 6936
rect 5971 6896 6029 6902
rect 6544 6893 6550 6945
rect 6602 6933 6608 6945
rect 6739 6936 6797 6942
rect 6739 6933 6751 6936
rect 6602 6905 6751 6933
rect 6602 6893 6608 6905
rect 6739 6902 6751 6905
rect 6785 6902 6797 6936
rect 6739 6896 6797 6902
rect 6928 6893 6934 6945
rect 6986 6933 6992 6945
rect 7507 6936 7565 6942
rect 7507 6933 7519 6936
rect 6986 6905 7519 6933
rect 6986 6893 6992 6905
rect 7507 6902 7519 6905
rect 7553 6902 7565 6936
rect 7507 6896 7565 6902
rect 7603 6936 7661 6942
rect 7603 6902 7615 6936
rect 7649 6933 7661 6936
rect 7792 6933 7798 6945
rect 7649 6905 7798 6933
rect 7649 6902 7661 6905
rect 7603 6896 7661 6902
rect 7792 6893 7798 6905
rect 7850 6893 7856 6945
rect 8275 6936 8333 6942
rect 8275 6902 8287 6936
rect 8321 6902 8333 6936
rect 8275 6896 8333 6902
rect 8371 6936 8429 6942
rect 8371 6902 8383 6936
rect 8417 6902 8429 6936
rect 9712 6933 9718 6945
rect 9673 6905 9718 6933
rect 8371 6896 8429 6902
rect 7312 6819 7318 6871
rect 7370 6859 7376 6871
rect 8290 6859 8318 6896
rect 7370 6831 8318 6859
rect 7370 6819 7376 6831
rect 3722 6757 5246 6785
rect 8083 6788 8141 6794
rect 3722 6745 3728 6757
rect 8083 6754 8095 6788
rect 8129 6785 8141 6788
rect 8386 6785 8414 6896
rect 9712 6893 9718 6905
rect 9770 6893 9776 6945
rect 9808 6893 9814 6945
rect 9866 6933 9872 6945
rect 9866 6905 9911 6933
rect 9866 6893 9872 6905
rect 9523 6862 9581 6868
rect 9523 6828 9535 6862
rect 9569 6859 9581 6862
rect 9826 6859 9854 6893
rect 9569 6831 9854 6859
rect 10018 6859 10046 6979
rect 11248 6967 11254 6979
rect 11306 6967 11312 7019
rect 12688 7007 12694 7019
rect 12649 6979 12694 7007
rect 12688 6967 12694 6979
rect 12746 6967 12752 7019
rect 12946 7007 12974 7053
rect 13651 7050 13663 7053
rect 13697 7050 13709 7084
rect 15088 7081 15094 7093
rect 15049 7053 15094 7081
rect 13651 7044 13709 7050
rect 15088 7041 15094 7053
rect 15146 7041 15152 7093
rect 15859 7084 15917 7090
rect 15859 7050 15871 7084
rect 15905 7081 15917 7084
rect 15952 7081 15958 7093
rect 15905 7053 15958 7081
rect 15905 7050 15917 7053
rect 15859 7044 15917 7050
rect 15952 7041 15958 7053
rect 16010 7041 16016 7093
rect 17890 7081 17918 7127
rect 18064 7081 18070 7093
rect 16066 7053 17918 7081
rect 18025 7053 18070 7081
rect 16066 7007 16094 7053
rect 18064 7041 18070 7053
rect 18122 7041 18128 7093
rect 18178 7081 18206 7127
rect 18754 7127 22814 7155
rect 18754 7081 18782 7127
rect 18178 7053 18782 7081
rect 18835 7084 18893 7090
rect 18835 7050 18847 7084
rect 18881 7081 18893 7084
rect 18928 7081 18934 7093
rect 18881 7053 18934 7081
rect 18881 7050 18893 7053
rect 18835 7044 18893 7050
rect 18928 7041 18934 7053
rect 18986 7041 18992 7093
rect 20368 7081 20374 7093
rect 20329 7053 20374 7081
rect 20368 7041 20374 7053
rect 20426 7041 20432 7093
rect 20851 7084 20909 7090
rect 20851 7050 20863 7084
rect 20897 7081 20909 7084
rect 21136 7081 21142 7093
rect 20897 7053 21142 7081
rect 20897 7050 20909 7053
rect 20851 7044 20909 7050
rect 21136 7041 21142 7053
rect 21194 7041 21200 7093
rect 21904 7081 21910 7093
rect 21865 7053 21910 7081
rect 21904 7041 21910 7053
rect 21962 7041 21968 7093
rect 22672 7081 22678 7093
rect 22633 7053 22678 7081
rect 22672 7041 22678 7053
rect 22730 7041 22736 7093
rect 22786 7081 22814 7127
rect 23056 7115 23062 7167
rect 23114 7155 23120 7167
rect 28162 7155 28190 7201
rect 28336 7155 28342 7167
rect 23114 7127 23486 7155
rect 23114 7115 23120 7127
rect 23344 7081 23350 7093
rect 22786 7053 23350 7081
rect 23344 7041 23350 7053
rect 23402 7041 23408 7093
rect 23458 7090 23486 7127
rect 25090 7127 28190 7155
rect 28297 7127 28342 7155
rect 23443 7084 23501 7090
rect 23443 7050 23455 7084
rect 23489 7050 23501 7084
rect 23443 7044 23501 7050
rect 23923 7084 23981 7090
rect 23923 7050 23935 7084
rect 23969 7081 23981 7084
rect 24211 7084 24269 7090
rect 24211 7081 24223 7084
rect 23969 7053 24223 7081
rect 23969 7050 23981 7053
rect 23923 7044 23981 7050
rect 24211 7050 24223 7053
rect 24257 7081 24269 7084
rect 24304 7081 24310 7093
rect 24257 7053 24310 7081
rect 24257 7050 24269 7053
rect 24211 7044 24269 7050
rect 24304 7041 24310 7053
rect 24362 7041 24368 7093
rect 12946 6979 16094 7007
rect 16339 7010 16397 7016
rect 16339 6976 16351 7010
rect 16385 7007 16397 7010
rect 16624 7007 16630 7019
rect 16385 6979 16630 7007
rect 16385 6976 16397 6979
rect 16339 6970 16397 6976
rect 16624 6967 16630 6979
rect 16682 6967 16688 7019
rect 25090 7007 25118 7127
rect 28336 7115 28342 7127
rect 28394 7155 28400 7167
rect 28394 7127 28670 7155
rect 28394 7115 28400 7127
rect 25456 7041 25462 7093
rect 25514 7081 25520 7093
rect 25651 7084 25709 7090
rect 25651 7081 25663 7084
rect 25514 7053 25663 7081
rect 25514 7041 25520 7053
rect 25651 7050 25663 7053
rect 25697 7050 25709 7084
rect 25651 7044 25709 7050
rect 26131 7084 26189 7090
rect 26131 7050 26143 7084
rect 26177 7081 26189 7084
rect 26320 7081 26326 7093
rect 26177 7053 26326 7081
rect 26177 7050 26189 7053
rect 26131 7044 26189 7050
rect 26320 7041 26326 7053
rect 26378 7041 26384 7093
rect 26899 7084 26957 7090
rect 26899 7050 26911 7084
rect 26945 7081 26957 7084
rect 27187 7084 27245 7090
rect 27187 7081 27199 7084
rect 26945 7053 27199 7081
rect 26945 7050 26957 7053
rect 26899 7044 26957 7050
rect 27187 7050 27199 7053
rect 27233 7081 27245 7084
rect 27280 7081 27286 7093
rect 27233 7053 27286 7081
rect 27233 7050 27245 7053
rect 27187 7044 27245 7050
rect 27280 7041 27286 7053
rect 27338 7041 27344 7093
rect 27952 7081 27958 7093
rect 27913 7053 27958 7081
rect 27952 7041 27958 7053
rect 28010 7041 28016 7093
rect 28642 7090 28670 7127
rect 29008 7115 29014 7167
rect 29066 7155 29072 7167
rect 29107 7158 29165 7164
rect 29107 7155 29119 7158
rect 29066 7127 29119 7155
rect 29066 7115 29072 7127
rect 29107 7124 29119 7127
rect 29153 7155 29165 7158
rect 29506 7155 29534 7201
rect 44563 7198 44575 7232
rect 44609 7198 44621 7232
rect 44563 7192 44621 7198
rect 32176 7155 32182 7167
rect 29153 7127 29438 7155
rect 29506 7127 32182 7155
rect 29153 7124 29165 7127
rect 29107 7118 29165 7124
rect 29410 7090 29438 7127
rect 32176 7115 32182 7127
rect 32234 7115 32240 7167
rect 33712 7155 33718 7167
rect 33673 7127 33718 7155
rect 33712 7115 33718 7127
rect 33770 7115 33776 7167
rect 37648 7115 37654 7167
rect 37706 7155 37712 7167
rect 39267 7158 39325 7164
rect 39267 7155 39279 7158
rect 37706 7127 39279 7155
rect 37706 7115 37712 7127
rect 39267 7124 39279 7127
rect 39313 7124 39325 7158
rect 41104 7155 41110 7167
rect 41065 7127 41110 7155
rect 39267 7118 39325 7124
rect 41104 7115 41110 7127
rect 41162 7155 41168 7167
rect 41162 7127 41438 7155
rect 41162 7115 41168 7127
rect 28627 7084 28685 7090
rect 28627 7050 28639 7084
rect 28673 7050 28685 7084
rect 28627 7044 28685 7050
rect 29395 7084 29453 7090
rect 29395 7050 29407 7084
rect 29441 7050 29453 7084
rect 29395 7044 29453 7050
rect 30931 7084 30989 7090
rect 30931 7050 30943 7084
rect 30977 7081 30989 7084
rect 31024 7081 31030 7093
rect 30977 7053 31030 7081
rect 30977 7050 30989 7053
rect 30931 7044 30989 7050
rect 31024 7041 31030 7053
rect 31082 7041 31088 7093
rect 31411 7084 31469 7090
rect 31411 7050 31423 7084
rect 31457 7081 31469 7084
rect 31696 7081 31702 7093
rect 31457 7053 31702 7081
rect 31457 7050 31469 7053
rect 31411 7044 31469 7050
rect 31696 7041 31702 7053
rect 31754 7041 31760 7093
rect 32467 7084 32525 7090
rect 32467 7050 32479 7084
rect 32513 7081 32525 7084
rect 32656 7081 32662 7093
rect 32513 7053 32662 7081
rect 32513 7050 32525 7053
rect 32467 7044 32525 7050
rect 32656 7041 32662 7053
rect 32714 7041 32720 7093
rect 33232 7081 33238 7093
rect 33193 7053 33238 7081
rect 33232 7041 33238 7053
rect 33290 7041 33296 7093
rect 33730 7081 33758 7115
rect 33907 7084 33965 7090
rect 33907 7081 33919 7084
rect 33730 7053 33919 7081
rect 33907 7050 33919 7053
rect 33953 7050 33965 7084
rect 34768 7081 34774 7093
rect 34729 7053 34774 7081
rect 33907 7044 33965 7050
rect 34768 7041 34774 7053
rect 34826 7041 34832 7093
rect 36208 7081 36214 7093
rect 36169 7053 36214 7081
rect 36208 7041 36214 7053
rect 36266 7041 36272 7093
rect 37459 7084 37517 7090
rect 37459 7050 37471 7084
rect 37505 7081 37517 7084
rect 37744 7081 37750 7093
rect 37505 7053 37750 7081
rect 37505 7050 37517 7053
rect 37459 7044 37517 7050
rect 37744 7041 37750 7053
rect 37802 7041 37808 7093
rect 38512 7081 38518 7093
rect 38473 7053 38518 7081
rect 38512 7041 38518 7053
rect 38570 7041 38576 7093
rect 41410 7090 41438 7127
rect 41488 7115 41494 7167
rect 41546 7155 41552 7167
rect 42179 7158 42237 7164
rect 42179 7155 42191 7158
rect 41546 7127 42191 7155
rect 41546 7115 41552 7127
rect 42179 7124 42191 7127
rect 42225 7124 42237 7158
rect 42179 7118 42237 7124
rect 43600 7115 43606 7167
rect 43658 7155 43664 7167
rect 44578 7155 44606 7192
rect 48784 7155 48790 7167
rect 43658 7127 44606 7155
rect 48745 7127 48790 7155
rect 43658 7115 43664 7127
rect 48784 7115 48790 7127
rect 48842 7155 48848 7167
rect 49267 7158 49325 7164
rect 49267 7155 49279 7158
rect 48842 7127 49279 7155
rect 48842 7115 48848 7127
rect 39187 7084 39245 7090
rect 39187 7050 39199 7084
rect 39233 7081 39245 7084
rect 39475 7084 39533 7090
rect 39475 7081 39487 7084
rect 39233 7053 39487 7081
rect 39233 7050 39245 7053
rect 39187 7044 39245 7050
rect 39475 7050 39487 7053
rect 39521 7050 39533 7084
rect 39475 7044 39533 7050
rect 41395 7084 41453 7090
rect 41395 7050 41407 7084
rect 41441 7081 41453 7084
rect 41683 7084 41741 7090
rect 41683 7081 41695 7084
rect 41441 7053 41695 7081
rect 41441 7050 41453 7053
rect 41395 7044 41453 7050
rect 41683 7050 41695 7053
rect 41729 7050 41741 7084
rect 43024 7081 43030 7093
rect 42985 7053 43030 7081
rect 41683 7044 41741 7050
rect 43024 7041 43030 7053
rect 43082 7041 43088 7093
rect 43792 7081 43798 7093
rect 43753 7053 43798 7081
rect 43792 7041 43798 7053
rect 43850 7041 43856 7093
rect 44272 7041 44278 7093
rect 44330 7081 44336 7093
rect 44330 7053 44510 7081
rect 44330 7041 44336 7053
rect 16738 6979 25118 7007
rect 10576 6933 10582 6945
rect 10537 6905 10582 6933
rect 10576 6893 10582 6905
rect 10634 6893 10640 6945
rect 13456 6893 13462 6945
rect 13514 6933 13520 6945
rect 13555 6936 13613 6942
rect 13555 6933 13567 6936
rect 13514 6905 13567 6933
rect 13514 6893 13520 6905
rect 13555 6902 13567 6905
rect 13601 6902 13613 6936
rect 13555 6896 13613 6902
rect 14608 6893 14614 6945
rect 14666 6933 14672 6945
rect 14995 6936 15053 6942
rect 14995 6933 15007 6936
rect 14666 6905 15007 6933
rect 14666 6893 14672 6905
rect 14995 6902 15007 6905
rect 15041 6902 15053 6936
rect 14995 6896 15053 6902
rect 15376 6893 15382 6945
rect 15434 6933 15440 6945
rect 15763 6936 15821 6942
rect 15763 6933 15775 6936
rect 15434 6905 15775 6933
rect 15434 6893 15440 6905
rect 15763 6902 15775 6905
rect 15809 6902 15821 6936
rect 15763 6896 15821 6902
rect 16738 6859 16766 6979
rect 25168 6967 25174 7019
rect 25226 7007 25232 7019
rect 25226 6979 25694 7007
rect 25226 6967 25232 6979
rect 17296 6893 17302 6945
rect 17354 6933 17360 6945
rect 17354 6905 17399 6933
rect 17354 6893 17360 6905
rect 19504 6893 19510 6945
rect 19562 6933 19568 6945
rect 20275 6936 20333 6942
rect 20275 6933 20287 6936
rect 19562 6905 20287 6933
rect 19562 6893 19568 6905
rect 20275 6902 20287 6905
rect 20321 6902 20333 6936
rect 20275 6896 20333 6902
rect 20368 6893 20374 6945
rect 20426 6933 20432 6945
rect 21043 6936 21101 6942
rect 21043 6933 21055 6936
rect 20426 6905 21055 6933
rect 20426 6893 20432 6905
rect 21043 6902 21055 6905
rect 21089 6902 21101 6936
rect 21043 6896 21101 6902
rect 21136 6893 21142 6945
rect 21194 6933 21200 6945
rect 21811 6936 21869 6942
rect 21811 6933 21823 6936
rect 21194 6905 21823 6933
rect 21194 6893 21200 6905
rect 21811 6902 21823 6905
rect 21857 6902 21869 6936
rect 21811 6896 21869 6902
rect 21904 6893 21910 6945
rect 21962 6933 21968 6945
rect 22579 6936 22637 6942
rect 22579 6933 22591 6936
rect 21962 6905 22591 6933
rect 21962 6893 21968 6905
rect 22579 6902 22591 6905
rect 22625 6902 22637 6936
rect 22579 6896 22637 6902
rect 22672 6893 22678 6945
rect 22730 6933 22736 6945
rect 23347 6936 23405 6942
rect 23347 6933 23359 6936
rect 22730 6905 23359 6933
rect 22730 6893 22736 6905
rect 23347 6902 23359 6905
rect 23393 6902 23405 6936
rect 23347 6896 23405 6902
rect 23440 6893 23446 6945
rect 23498 6933 23504 6945
rect 24115 6936 24173 6942
rect 24115 6933 24127 6936
rect 23498 6905 24127 6933
rect 23498 6893 23504 6905
rect 24115 6902 24127 6905
rect 24161 6902 24173 6936
rect 24115 6896 24173 6902
rect 24496 6893 24502 6945
rect 24554 6933 24560 6945
rect 25555 6936 25613 6942
rect 25555 6933 25567 6936
rect 24554 6905 25567 6933
rect 24554 6893 24560 6905
rect 25555 6902 25567 6905
rect 25601 6902 25613 6936
rect 25666 6933 25694 6979
rect 25936 6967 25942 7019
rect 25994 7007 26000 7019
rect 25994 6979 26558 7007
rect 25994 6967 26000 6979
rect 26419 6936 26477 6942
rect 26419 6933 26431 6936
rect 25666 6905 26431 6933
rect 25555 6896 25613 6902
rect 26419 6902 26431 6905
rect 26465 6902 26477 6936
rect 26530 6933 26558 6979
rect 26992 6967 26998 7019
rect 27050 7007 27056 7019
rect 27050 6979 27902 7007
rect 27050 6967 27056 6979
rect 27874 6942 27902 6979
rect 28528 6967 28534 7019
rect 28586 7007 28592 7019
rect 28586 6979 29534 7007
rect 28586 6967 28592 6979
rect 27091 6936 27149 6942
rect 27091 6933 27103 6936
rect 26530 6905 27103 6933
rect 26419 6896 26477 6902
rect 27091 6902 27103 6905
rect 27137 6902 27149 6936
rect 27091 6896 27149 6902
rect 27859 6936 27917 6942
rect 27859 6902 27871 6936
rect 27905 6902 27917 6936
rect 27859 6896 27917 6902
rect 27952 6893 27958 6945
rect 28010 6933 28016 6945
rect 29506 6942 29534 6979
rect 30736 6967 30742 7019
rect 30794 7007 30800 7019
rect 30794 6979 31646 7007
rect 30794 6967 30800 6979
rect 28723 6936 28781 6942
rect 28723 6933 28735 6936
rect 28010 6905 28735 6933
rect 28010 6893 28016 6905
rect 28723 6902 28735 6905
rect 28769 6902 28781 6936
rect 28723 6896 28781 6902
rect 29491 6936 29549 6942
rect 29491 6902 29503 6936
rect 29537 6902 29549 6936
rect 29491 6896 29549 6902
rect 29968 6893 29974 6945
rect 30026 6933 30032 6945
rect 31618 6942 31646 6979
rect 32176 6967 32182 7019
rect 32234 7007 32240 7019
rect 32234 6979 32510 7007
rect 32234 6967 32240 6979
rect 30835 6936 30893 6942
rect 30835 6933 30847 6936
rect 30026 6905 30847 6933
rect 30026 6893 30032 6905
rect 30835 6902 30847 6905
rect 30881 6902 30893 6936
rect 30835 6896 30893 6902
rect 31603 6936 31661 6942
rect 31603 6902 31615 6936
rect 31649 6902 31661 6936
rect 31603 6896 31661 6902
rect 31696 6893 31702 6945
rect 31754 6933 31760 6945
rect 32371 6936 32429 6942
rect 32371 6933 32383 6936
rect 31754 6905 32383 6933
rect 31754 6893 31760 6905
rect 32371 6902 32383 6905
rect 32417 6902 32429 6936
rect 32482 6933 32510 6979
rect 34480 6967 34486 7019
rect 34538 7007 34544 7019
rect 36979 7010 37037 7016
rect 36979 7007 36991 7010
rect 34538 6979 36991 7007
rect 34538 6967 34544 6979
rect 36979 6976 36991 6979
rect 37025 6976 37037 7010
rect 36979 6970 37037 6976
rect 37360 6967 37366 7019
rect 37418 7007 37424 7019
rect 40051 7010 40109 7016
rect 37418 6979 38462 7007
rect 37418 6967 37424 6979
rect 33139 6936 33197 6942
rect 33139 6933 33151 6936
rect 32482 6905 33151 6933
rect 32371 6896 32429 6902
rect 33139 6902 33151 6905
rect 33185 6902 33197 6936
rect 33139 6896 33197 6902
rect 33712 6893 33718 6945
rect 33770 6933 33776 6945
rect 34003 6936 34061 6942
rect 34003 6933 34015 6936
rect 33770 6905 34015 6933
rect 33770 6893 33776 6905
rect 34003 6902 34015 6905
rect 34049 6902 34061 6936
rect 34003 6896 34061 6902
rect 34096 6893 34102 6945
rect 34154 6933 34160 6945
rect 34675 6936 34733 6942
rect 34675 6933 34687 6936
rect 34154 6905 34687 6933
rect 34154 6893 34160 6905
rect 34675 6902 34687 6905
rect 34721 6902 34733 6936
rect 34675 6896 34733 6902
rect 35536 6893 35542 6945
rect 35594 6933 35600 6945
rect 36115 6936 36173 6942
rect 36115 6933 36127 6936
rect 35594 6905 36127 6933
rect 35594 6893 35600 6905
rect 36115 6902 36127 6905
rect 36161 6902 36173 6936
rect 36115 6896 36173 6902
rect 36496 6893 36502 6945
rect 36554 6933 36560 6945
rect 36883 6936 36941 6942
rect 36883 6933 36895 6936
rect 36554 6905 36895 6933
rect 36554 6893 36560 6905
rect 36883 6902 36895 6905
rect 36929 6902 36941 6936
rect 36883 6896 36941 6902
rect 37072 6893 37078 6945
rect 37130 6933 37136 6945
rect 38434 6942 38462 6979
rect 38530 6979 39998 7007
rect 38530 6945 38558 6979
rect 37651 6936 37709 6942
rect 37651 6933 37663 6936
rect 37130 6905 37663 6933
rect 37130 6893 37136 6905
rect 37651 6902 37663 6905
rect 37697 6902 37709 6936
rect 37651 6896 37709 6902
rect 38419 6936 38477 6942
rect 38419 6902 38431 6936
rect 38465 6902 38477 6936
rect 38419 6896 38477 6902
rect 38512 6893 38518 6945
rect 38570 6893 38576 6945
rect 39970 6942 39998 6979
rect 40051 6976 40063 7010
rect 40097 7007 40109 7010
rect 44368 7007 44374 7019
rect 40097 6979 44374 7007
rect 40097 6976 40109 6979
rect 40051 6970 40109 6976
rect 44368 6967 44374 6979
rect 44426 6967 44432 7019
rect 44482 7007 44510 7053
rect 45136 7041 45142 7093
rect 45194 7081 45200 7093
rect 45331 7084 45389 7090
rect 45331 7081 45343 7084
rect 45194 7053 45343 7081
rect 45194 7041 45200 7053
rect 45331 7050 45343 7053
rect 45377 7050 45389 7084
rect 45331 7044 45389 7050
rect 47344 7041 47350 7093
rect 47402 7081 47408 7093
rect 48994 7090 49022 7127
rect 49267 7124 49279 7127
rect 49313 7124 49325 7158
rect 49936 7155 49942 7167
rect 49897 7127 49942 7155
rect 49267 7118 49325 7124
rect 49936 7115 49942 7127
rect 49994 7155 50000 7167
rect 50515 7158 50573 7164
rect 50515 7155 50527 7158
rect 49994 7127 50527 7155
rect 49994 7115 50000 7127
rect 50242 7090 50270 7127
rect 50515 7124 50527 7127
rect 50561 7124 50573 7158
rect 50515 7118 50573 7124
rect 48307 7084 48365 7090
rect 48307 7081 48319 7084
rect 47402 7053 48319 7081
rect 47402 7041 47408 7053
rect 48307 7050 48319 7053
rect 48353 7050 48365 7084
rect 48307 7044 48365 7050
rect 48979 7084 49037 7090
rect 48979 7050 48991 7084
rect 49025 7050 49037 7084
rect 48979 7044 49037 7050
rect 50227 7084 50285 7090
rect 50227 7050 50239 7084
rect 50273 7050 50285 7084
rect 52048 7081 52054 7093
rect 52009 7053 52054 7081
rect 50227 7044 50285 7050
rect 52048 7041 52054 7053
rect 52106 7041 52112 7093
rect 47251 7010 47309 7016
rect 44482 6979 45278 7007
rect 39955 6936 40013 6942
rect 39394 6905 39806 6933
rect 38128 6859 38134 6871
rect 10018 6831 16766 6859
rect 17266 6831 31646 6859
rect 9569 6828 9581 6831
rect 9523 6822 9581 6828
rect 8659 6788 8717 6794
rect 8659 6785 8671 6788
rect 8129 6757 8671 6785
rect 8129 6754 8141 6757
rect 8083 6748 8141 6754
rect 8659 6754 8671 6757
rect 8705 6785 8717 6788
rect 17266 6785 17294 6831
rect 8705 6757 17294 6785
rect 31618 6785 31646 6831
rect 33106 6831 38134 6859
rect 33106 6785 33134 6831
rect 38128 6819 38134 6831
rect 38186 6819 38192 6871
rect 38224 6819 38230 6871
rect 38282 6859 38288 6871
rect 39394 6859 39422 6905
rect 38282 6831 39422 6859
rect 39475 6862 39533 6868
rect 38282 6819 38288 6831
rect 39475 6828 39487 6862
rect 39521 6828 39533 6862
rect 39475 6822 39533 6828
rect 31618 6757 33134 6785
rect 8705 6754 8717 6757
rect 8659 6748 8717 6754
rect 36400 6745 36406 6797
rect 36458 6785 36464 6797
rect 38899 6788 38957 6794
rect 38899 6785 38911 6788
rect 36458 6757 38911 6785
rect 36458 6745 36464 6757
rect 38899 6754 38911 6757
rect 38945 6785 38957 6788
rect 39490 6785 39518 6822
rect 38945 6757 39518 6785
rect 39778 6785 39806 6905
rect 39955 6902 39967 6936
rect 40001 6902 40013 6936
rect 39955 6896 40013 6902
rect 41491 6936 41549 6942
rect 41491 6902 41503 6936
rect 41537 6902 41549 6936
rect 42256 6933 42262 6945
rect 42217 6905 42262 6933
rect 41491 6896 41549 6902
rect 39856 6819 39862 6871
rect 39914 6859 39920 6871
rect 41506 6859 41534 6896
rect 42256 6893 42262 6905
rect 42314 6893 42320 6945
rect 42931 6936 42989 6942
rect 42931 6902 42943 6936
rect 42977 6902 42989 6936
rect 42931 6896 42989 6902
rect 39914 6831 41534 6859
rect 39914 6819 39920 6831
rect 41584 6819 41590 6871
rect 41642 6859 41648 6871
rect 42946 6859 42974 6896
rect 43024 6893 43030 6945
rect 43082 6933 43088 6945
rect 45250 6942 45278 6979
rect 47251 6976 47263 7010
rect 47297 7007 47309 7010
rect 47539 7010 47597 7016
rect 47539 7007 47551 7010
rect 47297 6979 47551 7007
rect 47297 6976 47309 6979
rect 47251 6970 47309 6976
rect 47539 6976 47551 6979
rect 47585 7007 47597 7010
rect 52528 7007 52534 7019
rect 47585 6979 52534 7007
rect 47585 6976 47597 6979
rect 47539 6970 47597 6976
rect 52528 6967 52534 6979
rect 52586 6967 52592 7019
rect 54067 7010 54125 7016
rect 54067 6976 54079 7010
rect 54113 6976 54125 7010
rect 54736 7007 54742 7019
rect 54697 6979 54742 7007
rect 54067 6970 54125 6976
rect 43699 6936 43757 6942
rect 43699 6933 43711 6936
rect 43082 6905 43711 6933
rect 43082 6893 43088 6905
rect 43699 6902 43711 6905
rect 43745 6902 43757 6936
rect 44467 6936 44525 6942
rect 44467 6933 44479 6936
rect 43699 6896 43757 6902
rect 43906 6905 44479 6933
rect 41642 6831 42974 6859
rect 41642 6819 41648 6831
rect 43906 6785 43934 6905
rect 44467 6902 44479 6905
rect 44513 6902 44525 6936
rect 44467 6896 44525 6902
rect 45235 6936 45293 6942
rect 45235 6902 45247 6936
rect 45281 6902 45293 6936
rect 46387 6936 46445 6942
rect 46387 6933 46399 6936
rect 45235 6896 45293 6902
rect 45634 6905 46399 6933
rect 43984 6819 43990 6871
rect 44042 6859 44048 6871
rect 45634 6859 45662 6905
rect 46387 6902 46399 6905
rect 46433 6933 46445 6936
rect 46675 6936 46733 6942
rect 46675 6933 46687 6936
rect 46433 6905 46687 6933
rect 46433 6902 46445 6905
rect 46387 6896 46445 6902
rect 46675 6902 46687 6905
rect 46721 6902 46733 6936
rect 46675 6896 46733 6902
rect 46771 6936 46829 6942
rect 46771 6902 46783 6936
rect 46817 6902 46829 6936
rect 46771 6896 46829 6902
rect 44042 6831 45662 6859
rect 44042 6819 44048 6831
rect 45712 6819 45718 6871
rect 45770 6859 45776 6871
rect 46786 6859 46814 6896
rect 47056 6893 47062 6945
rect 47114 6933 47120 6945
rect 47443 6936 47501 6942
rect 47443 6933 47455 6936
rect 47114 6905 47455 6933
rect 47114 6893 47120 6905
rect 47443 6902 47455 6905
rect 47489 6902 47501 6936
rect 47443 6896 47501 6902
rect 48211 6936 48269 6942
rect 48211 6902 48223 6936
rect 48257 6902 48269 6936
rect 48211 6896 48269 6902
rect 45770 6831 46814 6859
rect 45770 6819 45776 6831
rect 46864 6819 46870 6871
rect 46922 6859 46928 6871
rect 48226 6859 48254 6896
rect 48400 6893 48406 6945
rect 48458 6933 48464 6945
rect 49075 6936 49133 6942
rect 49075 6933 49087 6936
rect 48458 6905 49087 6933
rect 48458 6893 48464 6905
rect 49075 6902 49087 6905
rect 49121 6902 49133 6936
rect 49075 6896 49133 6902
rect 50323 6936 50381 6942
rect 50323 6902 50335 6936
rect 50369 6902 50381 6936
rect 50323 6896 50381 6902
rect 46922 6831 48254 6859
rect 46922 6819 46928 6831
rect 50128 6819 50134 6871
rect 50186 6859 50192 6871
rect 50338 6859 50366 6896
rect 50416 6893 50422 6945
rect 50474 6933 50480 6945
rect 51184 6933 51190 6945
rect 50474 6905 51190 6933
rect 50474 6893 50480 6905
rect 51184 6893 51190 6905
rect 51242 6893 51248 6945
rect 51568 6893 51574 6945
rect 51626 6933 51632 6945
rect 51955 6936 52013 6942
rect 51955 6933 51967 6936
rect 51626 6905 51967 6933
rect 51626 6893 51632 6905
rect 51955 6902 51967 6905
rect 52001 6902 52013 6936
rect 52723 6936 52781 6942
rect 52723 6933 52735 6936
rect 51955 6896 52013 6902
rect 52162 6905 52735 6933
rect 50186 6831 50366 6859
rect 50186 6819 50192 6831
rect 44179 6788 44237 6794
rect 44179 6785 44191 6788
rect 39778 6757 44191 6785
rect 38945 6754 38957 6757
rect 38899 6748 38957 6754
rect 44179 6754 44191 6757
rect 44225 6754 44237 6788
rect 44179 6748 44237 6754
rect 50224 6745 50230 6797
rect 50282 6785 50288 6797
rect 52162 6785 52190 6905
rect 52723 6902 52735 6905
rect 52769 6902 52781 6936
rect 52723 6896 52781 6902
rect 52819 6936 52877 6942
rect 52819 6902 52831 6936
rect 52865 6902 52877 6936
rect 54082 6933 54110 6970
rect 54736 6967 54742 6979
rect 54794 6967 54800 7019
rect 55408 6967 55414 7019
rect 55466 7007 55472 7019
rect 55507 7010 55565 7016
rect 55507 7007 55519 7010
rect 55466 6979 55519 7007
rect 55466 6967 55472 6979
rect 55507 6976 55519 6979
rect 55553 6976 55565 7010
rect 55507 6970 55565 6976
rect 57811 7010 57869 7016
rect 57811 6976 57823 7010
rect 57857 7007 57869 7010
rect 58480 7007 58486 7019
rect 57857 6979 58486 7007
rect 57857 6976 57869 6979
rect 57811 6970 57869 6976
rect 58480 6967 58486 6979
rect 58538 6967 58544 7019
rect 57040 6933 57046 6945
rect 54082 6905 57046 6933
rect 52819 6896 52877 6902
rect 52240 6819 52246 6871
rect 52298 6859 52304 6871
rect 52834 6859 52862 6896
rect 57040 6893 57046 6905
rect 57098 6893 57104 6945
rect 52298 6831 52862 6859
rect 52298 6819 52304 6831
rect 52435 6788 52493 6794
rect 52435 6785 52447 6788
rect 50282 6757 52447 6785
rect 50282 6745 50288 6757
rect 52435 6754 52447 6757
rect 52481 6754 52493 6788
rect 52435 6748 52493 6754
rect 1152 6686 58848 6708
rect 1152 6634 4294 6686
rect 4346 6634 4358 6686
rect 4410 6634 4422 6686
rect 4474 6634 4486 6686
rect 4538 6634 35014 6686
rect 35066 6634 35078 6686
rect 35130 6634 35142 6686
rect 35194 6634 35206 6686
rect 35258 6634 58848 6686
rect 1152 6612 58848 6634
rect 5392 6563 5398 6575
rect 5353 6535 5398 6563
rect 5392 6523 5398 6535
rect 5450 6563 5456 6575
rect 5450 6535 5726 6563
rect 5450 6523 5456 6535
rect 5698 6424 5726 6535
rect 6640 6523 6646 6575
rect 6698 6563 6704 6575
rect 10576 6563 10582 6575
rect 6698 6535 10582 6563
rect 6698 6523 6704 6535
rect 10576 6523 10582 6535
rect 10634 6523 10640 6575
rect 13072 6523 13078 6575
rect 13130 6563 13136 6575
rect 14032 6563 14038 6575
rect 13130 6535 14038 6563
rect 13130 6523 13136 6535
rect 14032 6523 14038 6535
rect 14090 6523 14096 6575
rect 18832 6563 18838 6575
rect 18793 6535 18838 6563
rect 18832 6523 18838 6535
rect 18890 6523 18896 6575
rect 20467 6566 20525 6572
rect 20467 6532 20479 6566
rect 20513 6563 20525 6566
rect 20560 6563 20566 6575
rect 20513 6535 20566 6563
rect 20513 6532 20525 6535
rect 20467 6526 20525 6532
rect 20560 6523 20566 6535
rect 20618 6523 20624 6575
rect 22576 6563 22582 6575
rect 22537 6535 22582 6563
rect 22576 6523 22582 6535
rect 22634 6523 22640 6575
rect 24112 6563 24118 6575
rect 24073 6535 24118 6563
rect 24112 6523 24118 6535
rect 24170 6523 24176 6575
rect 27856 6563 27862 6575
rect 27817 6535 27862 6563
rect 27856 6523 27862 6535
rect 27914 6523 27920 6575
rect 31792 6563 31798 6575
rect 31753 6535 31798 6563
rect 31792 6523 31798 6535
rect 31850 6523 31856 6575
rect 42256 6523 42262 6575
rect 42314 6563 42320 6575
rect 45427 6566 45485 6572
rect 45427 6563 45439 6566
rect 42314 6535 45439 6563
rect 42314 6523 42320 6535
rect 45427 6532 45439 6535
rect 45473 6532 45485 6566
rect 45427 6526 45485 6532
rect 46195 6566 46253 6572
rect 46195 6532 46207 6566
rect 46241 6563 46253 6566
rect 46480 6563 46486 6575
rect 46241 6535 46486 6563
rect 46241 6532 46253 6535
rect 46195 6526 46253 6532
rect 46480 6523 46486 6535
rect 46538 6523 46544 6575
rect 49648 6523 49654 6575
rect 49706 6563 49712 6575
rect 50515 6566 50573 6572
rect 50515 6563 50527 6566
rect 49706 6535 50527 6563
rect 49706 6523 49712 6535
rect 50515 6532 50527 6535
rect 50561 6563 50573 6566
rect 51280 6563 51286 6575
rect 50561 6535 51038 6563
rect 51241 6535 51286 6563
rect 50561 6532 50573 6535
rect 50515 6526 50573 6532
rect 7603 6492 7661 6498
rect 7603 6458 7615 6492
rect 7649 6489 7661 6492
rect 9232 6489 9238 6501
rect 7649 6461 9238 6489
rect 7649 6458 7661 6461
rect 7603 6452 7661 6458
rect 9232 6449 9238 6461
rect 9290 6449 9296 6501
rect 9808 6449 9814 6501
rect 9866 6489 9872 6501
rect 50416 6489 50422 6501
rect 9866 6461 50422 6489
rect 9866 6449 9872 6461
rect 50416 6449 50422 6461
rect 50474 6449 50480 6501
rect 5683 6418 5741 6424
rect 5683 6384 5695 6418
rect 5729 6384 5741 6418
rect 5683 6378 5741 6384
rect 6256 6375 6262 6427
rect 6314 6415 6320 6427
rect 7027 6418 7085 6424
rect 7027 6415 7039 6418
rect 6314 6387 7039 6415
rect 6314 6375 6320 6387
rect 7027 6384 7039 6387
rect 7073 6384 7085 6418
rect 7027 6378 7085 6384
rect 7120 6375 7126 6427
rect 7178 6415 7184 6427
rect 13651 6418 13709 6424
rect 7178 6387 7968 6415
rect 7178 6375 7184 6387
rect 13651 6384 13663 6418
rect 13697 6415 13709 6418
rect 13936 6415 13942 6427
rect 13697 6387 13942 6415
rect 13697 6384 13709 6387
rect 13651 6378 13709 6384
rect 13936 6375 13942 6387
rect 13994 6375 14000 6427
rect 14704 6415 14710 6427
rect 14665 6387 14710 6415
rect 14704 6375 14710 6387
rect 14762 6375 14768 6427
rect 15472 6415 15478 6427
rect 15433 6387 15478 6415
rect 15472 6375 15478 6387
rect 15530 6375 15536 6427
rect 16240 6415 16246 6427
rect 16201 6387 16246 6415
rect 16240 6375 16246 6387
rect 16298 6375 16304 6427
rect 17680 6415 17686 6427
rect 17641 6387 17686 6415
rect 17680 6375 17686 6387
rect 17738 6375 17744 6427
rect 18448 6415 18454 6427
rect 18409 6387 18454 6415
rect 18448 6375 18454 6387
rect 18506 6375 18512 6427
rect 18832 6375 18838 6427
rect 18890 6415 18896 6427
rect 19219 6418 19277 6424
rect 19219 6415 19231 6418
rect 18890 6387 19231 6415
rect 18890 6375 18896 6387
rect 19219 6384 19231 6387
rect 19265 6384 19277 6418
rect 19219 6378 19277 6384
rect 20560 6375 20566 6427
rect 20618 6415 20624 6427
rect 20755 6418 20813 6424
rect 20755 6415 20767 6418
rect 20618 6387 20767 6415
rect 20618 6375 20624 6387
rect 20755 6384 20767 6387
rect 20801 6384 20813 6418
rect 20755 6378 20813 6384
rect 21427 6418 21485 6424
rect 21427 6384 21439 6418
rect 21473 6384 21485 6418
rect 21427 6378 21485 6384
rect 1552 6341 1558 6353
rect 1513 6313 1558 6341
rect 1552 6301 1558 6313
rect 1610 6301 1616 6353
rect 2032 6301 2038 6353
rect 2090 6341 2096 6353
rect 2323 6344 2381 6350
rect 2323 6341 2335 6344
rect 2090 6313 2335 6341
rect 2090 6301 2096 6313
rect 2323 6310 2335 6313
rect 2369 6310 2381 6344
rect 3184 6341 3190 6353
rect 3145 6313 3190 6341
rect 2323 6304 2381 6310
rect 3184 6301 3190 6313
rect 3242 6301 3248 6353
rect 3856 6301 3862 6353
rect 3914 6341 3920 6353
rect 3955 6344 4013 6350
rect 3955 6341 3967 6344
rect 3914 6313 3967 6341
rect 3914 6301 3920 6313
rect 3955 6310 3967 6313
rect 4001 6310 4013 6344
rect 3955 6304 4013 6310
rect 4624 6301 4630 6353
rect 4682 6341 4688 6353
rect 4723 6344 4781 6350
rect 4723 6341 4735 6344
rect 4682 6313 4735 6341
rect 4682 6301 4688 6313
rect 4723 6310 4735 6313
rect 4769 6310 4781 6344
rect 9424 6341 9430 6353
rect 9385 6313 9430 6341
rect 4723 6304 4781 6310
rect 9424 6301 9430 6313
rect 9482 6301 9488 6353
rect 10096 6301 10102 6353
rect 10154 6341 10160 6353
rect 10195 6344 10253 6350
rect 10195 6341 10207 6344
rect 10154 6313 10207 6341
rect 10154 6301 10160 6313
rect 10195 6310 10207 6313
rect 10241 6310 10253 6344
rect 10195 6304 10253 6310
rect 10864 6301 10870 6353
rect 10922 6341 10928 6353
rect 10963 6344 11021 6350
rect 10963 6341 10975 6344
rect 10922 6313 10975 6341
rect 10922 6301 10928 6313
rect 10963 6310 10975 6313
rect 11009 6310 11021 6344
rect 10963 6304 11021 6310
rect 11632 6301 11638 6353
rect 11690 6341 11696 6353
rect 12211 6344 12269 6350
rect 12211 6341 12223 6344
rect 11690 6313 12223 6341
rect 11690 6301 11696 6313
rect 12211 6310 12223 6313
rect 12257 6310 12269 6344
rect 13072 6341 13078 6353
rect 13033 6313 13078 6341
rect 12211 6304 12269 6310
rect 13072 6301 13078 6313
rect 13130 6301 13136 6353
rect 15952 6301 15958 6353
rect 16010 6341 16016 6353
rect 19987 6344 20045 6350
rect 19987 6341 19999 6344
rect 16010 6313 19999 6341
rect 16010 6301 16016 6313
rect 19987 6310 19999 6313
rect 20033 6310 20045 6344
rect 19987 6304 20045 6310
rect 20080 6301 20086 6353
rect 20138 6341 20144 6353
rect 21442 6341 21470 6378
rect 22576 6375 22582 6427
rect 22634 6415 22640 6427
rect 22963 6418 23021 6424
rect 22963 6415 22975 6418
rect 22634 6387 22975 6415
rect 22634 6375 22640 6387
rect 22963 6384 22975 6387
rect 23009 6384 23021 6418
rect 23728 6415 23734 6427
rect 23689 6387 23734 6415
rect 22963 6378 23021 6384
rect 23728 6375 23734 6387
rect 23786 6375 23792 6427
rect 24112 6375 24118 6427
rect 24170 6415 24176 6427
rect 24403 6418 24461 6424
rect 24403 6415 24415 6418
rect 24170 6387 24415 6415
rect 24170 6375 24176 6387
rect 24403 6384 24415 6387
rect 24449 6384 24461 6418
rect 24403 6378 24461 6384
rect 27856 6375 27862 6427
rect 27914 6415 27920 6427
rect 28243 6418 28301 6424
rect 28243 6415 28255 6418
rect 27914 6387 28255 6415
rect 27914 6375 27920 6387
rect 28243 6384 28255 6387
rect 28289 6384 28301 6418
rect 28243 6378 28301 6384
rect 29011 6418 29069 6424
rect 29011 6384 29023 6418
rect 29057 6415 29069 6418
rect 29104 6415 29110 6427
rect 29057 6387 29110 6415
rect 29057 6384 29069 6387
rect 29011 6378 29069 6384
rect 29104 6375 29110 6387
rect 29162 6375 29168 6427
rect 30640 6415 30646 6427
rect 30601 6387 30646 6415
rect 30640 6375 30646 6387
rect 30698 6375 30704 6427
rect 31792 6375 31798 6427
rect 31850 6415 31856 6427
rect 32179 6418 32237 6424
rect 32179 6415 32191 6418
rect 31850 6387 32191 6415
rect 31850 6375 31856 6387
rect 32179 6384 32191 6387
rect 32225 6384 32237 6418
rect 34288 6415 34294 6427
rect 34249 6387 34294 6415
rect 32179 6378 32237 6384
rect 34288 6375 34294 6387
rect 34346 6375 34352 6427
rect 34864 6375 34870 6427
rect 34922 6415 34928 6427
rect 35059 6418 35117 6424
rect 35059 6415 35071 6418
rect 34922 6387 35071 6415
rect 34922 6375 34928 6387
rect 35059 6384 35071 6387
rect 35105 6384 35117 6418
rect 37264 6415 37270 6427
rect 37225 6387 37270 6415
rect 35059 6378 35117 6384
rect 37264 6375 37270 6387
rect 37322 6375 37328 6427
rect 41296 6415 41302 6427
rect 41257 6387 41302 6415
rect 41296 6375 41302 6387
rect 41354 6375 41360 6427
rect 42832 6415 42838 6427
rect 42793 6387 42838 6415
rect 42832 6375 42838 6387
rect 42890 6375 42896 6427
rect 44080 6415 44086 6427
rect 44041 6387 44086 6415
rect 44080 6375 44086 6387
rect 44138 6375 44144 6427
rect 44851 6418 44909 6424
rect 44851 6384 44863 6418
rect 44897 6415 44909 6418
rect 44944 6415 44950 6427
rect 44897 6387 44950 6415
rect 44897 6384 44909 6387
rect 44851 6378 44909 6384
rect 44944 6375 44950 6387
rect 45002 6375 45008 6427
rect 49840 6375 49846 6427
rect 49898 6415 49904 6427
rect 50899 6418 50957 6424
rect 50899 6415 50911 6418
rect 49898 6387 50911 6415
rect 49898 6375 49904 6387
rect 50899 6384 50911 6387
rect 50945 6384 50957 6418
rect 50899 6378 50957 6384
rect 20138 6313 21470 6341
rect 21523 6344 21581 6350
rect 20138 6301 20144 6313
rect 21523 6310 21535 6344
rect 21569 6341 21581 6344
rect 25360 6341 25366 6353
rect 21569 6313 25366 6341
rect 21569 6310 21581 6313
rect 21523 6304 21581 6310
rect 25360 6301 25366 6313
rect 25418 6301 25424 6353
rect 25648 6341 25654 6353
rect 25609 6313 25654 6341
rect 25648 6301 25654 6313
rect 25706 6301 25712 6353
rect 26800 6341 26806 6353
rect 26761 6313 26806 6341
rect 26800 6301 26806 6313
rect 26858 6301 26864 6353
rect 29680 6341 29686 6353
rect 29641 6313 29686 6341
rect 29680 6301 29686 6313
rect 29738 6301 29744 6353
rect 31216 6341 31222 6353
rect 31177 6313 31222 6341
rect 31216 6301 31222 6313
rect 31274 6301 31280 6353
rect 32560 6301 32566 6353
rect 32618 6341 32624 6353
rect 34211 6344 34269 6350
rect 34211 6341 34223 6344
rect 32618 6313 34223 6341
rect 32618 6301 32624 6313
rect 34211 6310 34223 6313
rect 34257 6310 34269 6344
rect 36304 6341 36310 6353
rect 36265 6313 36310 6341
rect 34211 6304 34269 6310
rect 36304 6301 36310 6313
rect 36362 6301 36368 6353
rect 38896 6341 38902 6353
rect 38857 6313 38902 6341
rect 38896 6301 38902 6313
rect 38954 6301 38960 6353
rect 40336 6341 40342 6353
rect 40297 6313 40342 6341
rect 40336 6301 40342 6313
rect 40394 6301 40400 6353
rect 41872 6341 41878 6353
rect 41833 6313 41878 6341
rect 41872 6301 41878 6313
rect 41930 6301 41936 6353
rect 45520 6341 45526 6353
rect 45481 6313 45526 6341
rect 45520 6301 45526 6313
rect 45578 6301 45584 6353
rect 46960 6341 46966 6353
rect 46921 6313 46966 6341
rect 46960 6301 46966 6313
rect 47018 6301 47024 6353
rect 47728 6341 47734 6353
rect 47689 6313 47734 6341
rect 47728 6301 47734 6313
rect 47786 6301 47792 6353
rect 48784 6301 48790 6353
rect 48842 6341 48848 6353
rect 49171 6344 49229 6350
rect 49171 6341 49183 6344
rect 48842 6313 49183 6341
rect 48842 6301 48848 6313
rect 49171 6310 49183 6313
rect 49217 6310 49229 6344
rect 49171 6304 49229 6310
rect 49552 6301 49558 6353
rect 49610 6341 49616 6353
rect 49939 6344 49997 6350
rect 49939 6341 49951 6344
rect 49610 6313 49951 6341
rect 49610 6301 49616 6313
rect 49939 6310 49951 6313
rect 49985 6310 49997 6344
rect 49939 6304 49997 6310
rect 50803 6344 50861 6350
rect 50803 6310 50815 6344
rect 50849 6341 50861 6344
rect 51010 6341 51038 6535
rect 51280 6523 51286 6535
rect 51338 6563 51344 6575
rect 51338 6535 51614 6563
rect 51338 6523 51344 6535
rect 51586 6424 51614 6535
rect 51571 6418 51629 6424
rect 51571 6384 51583 6418
rect 51617 6384 51629 6418
rect 51571 6378 51629 6384
rect 50849 6313 51038 6341
rect 50849 6310 50861 6313
rect 50803 6304 50861 6310
rect 51088 6301 51094 6353
rect 51146 6341 51152 6353
rect 52051 6344 52109 6350
rect 52051 6341 52063 6344
rect 51146 6313 52063 6341
rect 51146 6301 51152 6313
rect 52051 6310 52063 6313
rect 52097 6341 52109 6344
rect 52339 6344 52397 6350
rect 52339 6341 52351 6344
rect 52097 6313 52351 6341
rect 52097 6310 52109 6313
rect 52051 6304 52109 6310
rect 52339 6310 52351 6313
rect 52385 6310 52397 6344
rect 52339 6304 52397 6310
rect 53299 6344 53357 6350
rect 53299 6310 53311 6344
rect 53345 6310 53357 6344
rect 53299 6304 53357 6310
rect 6835 6270 6893 6276
rect 6835 6236 6847 6270
rect 6881 6267 6893 6270
rect 7120 6267 7126 6279
rect 6881 6239 7126 6267
rect 6881 6236 6893 6239
rect 6835 6230 6893 6236
rect 7120 6227 7126 6239
rect 7178 6227 7184 6279
rect 14896 6227 14902 6279
rect 14954 6267 14960 6279
rect 14954 6239 16190 6267
rect 14954 6227 14960 6239
rect 5200 6153 5206 6205
rect 5258 6193 5264 6205
rect 5258 6165 7838 6193
rect 5258 6153 5264 6165
rect 5488 6079 5494 6131
rect 5546 6119 5552 6131
rect 5587 6122 5645 6128
rect 5587 6119 5599 6122
rect 5546 6091 5599 6119
rect 5546 6079 5552 6091
rect 5587 6088 5599 6091
rect 5633 6088 5645 6122
rect 7810 6119 7838 6165
rect 8242 6119 8270 6179
rect 14224 6153 14230 6205
rect 14282 6193 14288 6205
rect 14282 6165 15422 6193
rect 14282 6153 14288 6165
rect 7810 6091 8270 6119
rect 5587 6082 5645 6088
rect 13744 6079 13750 6131
rect 13802 6119 13808 6131
rect 13843 6122 13901 6128
rect 13843 6119 13855 6122
rect 13802 6091 13855 6119
rect 13802 6079 13808 6091
rect 13843 6088 13855 6091
rect 13889 6088 13901 6122
rect 13843 6082 13901 6088
rect 13936 6079 13942 6131
rect 13994 6119 14000 6131
rect 15394 6128 15422 6165
rect 16162 6128 16190 6239
rect 19312 6227 19318 6279
rect 19370 6267 19376 6279
rect 19370 6239 20702 6267
rect 19370 6227 19376 6239
rect 18064 6153 18070 6205
rect 18122 6193 18128 6205
rect 18122 6165 18494 6193
rect 18122 6153 18128 6165
rect 14611 6122 14669 6128
rect 14611 6119 14623 6122
rect 13994 6091 14623 6119
rect 13994 6079 14000 6091
rect 14611 6088 14623 6091
rect 14657 6088 14669 6122
rect 14611 6082 14669 6088
rect 15379 6122 15437 6128
rect 15379 6088 15391 6122
rect 15425 6088 15437 6122
rect 15379 6082 15437 6088
rect 16147 6122 16205 6128
rect 16147 6088 16159 6122
rect 16193 6088 16205 6122
rect 16147 6082 16205 6088
rect 16720 6079 16726 6131
rect 16778 6119 16784 6131
rect 17587 6122 17645 6128
rect 17587 6119 17599 6122
rect 16778 6091 17599 6119
rect 16778 6079 16784 6091
rect 17587 6088 17599 6091
rect 17633 6088 17645 6122
rect 18352 6119 18358 6131
rect 18313 6091 18358 6119
rect 17587 6082 17645 6088
rect 18352 6079 18358 6091
rect 18410 6079 18416 6131
rect 18466 6119 18494 6165
rect 18928 6153 18934 6205
rect 18986 6193 18992 6205
rect 18986 6165 19934 6193
rect 18986 6153 18992 6165
rect 19906 6128 19934 6165
rect 20674 6128 20702 6239
rect 22960 6227 22966 6279
rect 23018 6267 23024 6279
rect 33520 6267 33526 6279
rect 23018 6239 24542 6267
rect 33481 6239 33526 6267
rect 23018 6227 23024 6239
rect 22288 6153 22294 6205
rect 22346 6193 22352 6205
rect 22346 6165 23054 6193
rect 22346 6153 22352 6165
rect 19123 6122 19181 6128
rect 19123 6119 19135 6122
rect 18466 6091 19135 6119
rect 19123 6088 19135 6091
rect 19169 6088 19181 6122
rect 19123 6082 19181 6088
rect 19891 6122 19949 6128
rect 19891 6088 19903 6122
rect 19937 6088 19949 6122
rect 19891 6082 19949 6088
rect 20659 6122 20717 6128
rect 20659 6088 20671 6122
rect 20705 6088 20717 6122
rect 22864 6119 22870 6131
rect 22825 6091 22870 6119
rect 20659 6082 20717 6088
rect 22864 6079 22870 6091
rect 22922 6079 22928 6131
rect 23026 6119 23054 6165
rect 24514 6128 24542 6239
rect 33520 6227 33526 6239
rect 33578 6227 33584 6279
rect 38128 6227 38134 6279
rect 38186 6267 38192 6279
rect 46672 6267 46678 6279
rect 38186 6239 46678 6267
rect 38186 6227 38192 6239
rect 46672 6227 46678 6239
rect 46730 6227 46736 6279
rect 52432 6267 52438 6279
rect 50386 6239 52438 6267
rect 27472 6153 27478 6205
rect 27530 6193 27536 6205
rect 27530 6165 28958 6193
rect 27530 6153 27536 6165
rect 23635 6122 23693 6128
rect 23635 6119 23647 6122
rect 23026 6091 23647 6119
rect 23635 6088 23647 6091
rect 23681 6088 23693 6122
rect 23635 6082 23693 6088
rect 24499 6122 24557 6128
rect 24499 6088 24511 6122
rect 24545 6088 24557 6122
rect 24499 6082 24557 6088
rect 26320 6079 26326 6131
rect 26378 6119 26384 6131
rect 28930 6128 28958 6165
rect 31792 6153 31798 6205
rect 31850 6193 31856 6205
rect 31850 6165 33470 6193
rect 31850 6153 31856 6165
rect 28147 6122 28205 6128
rect 28147 6119 28159 6122
rect 26378 6091 28159 6119
rect 26378 6079 26384 6091
rect 28147 6088 28159 6091
rect 28193 6088 28205 6122
rect 28147 6082 28205 6088
rect 28915 6122 28973 6128
rect 28915 6088 28927 6122
rect 28961 6088 28973 6122
rect 28915 6082 28973 6088
rect 29776 6079 29782 6131
rect 29834 6119 29840 6131
rect 30547 6122 30605 6128
rect 30547 6119 30559 6122
rect 29834 6091 30559 6119
rect 29834 6079 29840 6091
rect 30547 6088 30559 6091
rect 30593 6088 30605 6122
rect 30547 6082 30605 6088
rect 31504 6079 31510 6131
rect 31562 6119 31568 6131
rect 33442 6128 33470 6165
rect 40624 6153 40630 6205
rect 40682 6193 40688 6205
rect 40682 6165 41342 6193
rect 40682 6153 40688 6165
rect 32083 6122 32141 6128
rect 32083 6119 32095 6122
rect 31562 6091 32095 6119
rect 31562 6079 31568 6091
rect 32083 6088 32095 6091
rect 32129 6088 32141 6122
rect 32083 6082 32141 6088
rect 33427 6122 33485 6128
rect 33427 6088 33439 6122
rect 33473 6088 33485 6122
rect 33427 6082 33485 6088
rect 33808 6079 33814 6131
rect 33866 6119 33872 6131
rect 34963 6122 35021 6128
rect 34963 6119 34975 6122
rect 33866 6091 34975 6119
rect 33866 6079 33872 6091
rect 34963 6088 34975 6091
rect 35009 6088 35021 6122
rect 34963 6082 35021 6088
rect 35344 6079 35350 6131
rect 35402 6119 35408 6131
rect 37171 6122 37229 6128
rect 37171 6119 37183 6122
rect 35402 6091 37183 6119
rect 35402 6079 35408 6091
rect 37171 6088 37183 6091
rect 37217 6088 37229 6122
rect 37171 6082 37229 6088
rect 39184 6079 39190 6131
rect 39242 6119 39248 6131
rect 41203 6122 41261 6128
rect 41203 6119 41215 6122
rect 39242 6091 41215 6119
rect 39242 6079 39248 6091
rect 41203 6088 41215 6091
rect 41249 6088 41261 6122
rect 41314 6119 41342 6165
rect 42160 6153 42166 6205
rect 42218 6193 42224 6205
rect 45427 6196 45485 6202
rect 42218 6165 43214 6193
rect 42218 6153 42224 6165
rect 42739 6122 42797 6128
rect 42739 6119 42751 6122
rect 41314 6091 42751 6119
rect 41203 6082 41261 6088
rect 42739 6088 42751 6091
rect 42785 6088 42797 6122
rect 43186 6119 43214 6165
rect 45427 6162 45439 6196
rect 45473 6193 45485 6196
rect 50386 6193 50414 6239
rect 52432 6227 52438 6239
rect 52490 6227 52496 6279
rect 45473 6165 50414 6193
rect 45473 6162 45485 6165
rect 45427 6156 45485 6162
rect 51472 6153 51478 6205
rect 51530 6193 51536 6205
rect 53314 6193 53342 6304
rect 53968 6301 53974 6353
rect 54026 6341 54032 6353
rect 54451 6344 54509 6350
rect 54451 6341 54463 6344
rect 54026 6313 54463 6341
rect 54026 6301 54032 6313
rect 54451 6310 54463 6313
rect 54497 6310 54509 6344
rect 54451 6304 54509 6310
rect 54640 6301 54646 6353
rect 54698 6341 54704 6353
rect 55219 6344 55277 6350
rect 55219 6341 55231 6344
rect 54698 6313 55231 6341
rect 54698 6301 54704 6313
rect 55219 6310 55231 6313
rect 55265 6310 55277 6344
rect 55219 6304 55277 6310
rect 55987 6344 56045 6350
rect 55987 6310 55999 6344
rect 56033 6310 56045 6344
rect 55987 6304 56045 6310
rect 57043 6344 57101 6350
rect 57043 6310 57055 6344
rect 57089 6310 57101 6344
rect 57043 6304 57101 6310
rect 57811 6344 57869 6350
rect 57811 6310 57823 6344
rect 57857 6341 57869 6344
rect 58096 6341 58102 6353
rect 57857 6313 58102 6341
rect 57857 6310 57869 6313
rect 57811 6304 57869 6310
rect 55024 6227 55030 6279
rect 55082 6267 55088 6279
rect 56002 6267 56030 6304
rect 55082 6239 56030 6267
rect 57058 6267 57086 6304
rect 58096 6301 58102 6313
rect 58154 6301 58160 6353
rect 58864 6267 58870 6279
rect 57058 6239 58870 6267
rect 55082 6227 55088 6239
rect 58864 6227 58870 6239
rect 58922 6227 58928 6279
rect 56272 6193 56278 6205
rect 51530 6165 52478 6193
rect 53314 6165 56278 6193
rect 51530 6153 51536 6165
rect 43987 6122 44045 6128
rect 43987 6119 43999 6122
rect 43186 6091 43999 6119
rect 42739 6082 42797 6088
rect 43987 6088 43999 6091
rect 44033 6088 44045 6122
rect 43987 6082 44045 6088
rect 44176 6079 44182 6131
rect 44234 6119 44240 6131
rect 44755 6122 44813 6128
rect 44755 6119 44767 6122
rect 44234 6091 44767 6119
rect 44234 6079 44240 6091
rect 44755 6088 44767 6091
rect 44801 6088 44813 6122
rect 44755 6082 44813 6088
rect 51088 6079 51094 6131
rect 51146 6119 51152 6131
rect 52450 6128 52478 6165
rect 56272 6153 56278 6165
rect 56330 6153 56336 6205
rect 51667 6122 51725 6128
rect 51667 6119 51679 6122
rect 51146 6091 51679 6119
rect 51146 6079 51152 6091
rect 51667 6088 51679 6091
rect 51713 6088 51725 6122
rect 51667 6082 51725 6088
rect 52435 6122 52493 6128
rect 52435 6088 52447 6122
rect 52481 6088 52493 6122
rect 52435 6082 52493 6088
rect 1152 6020 58848 6042
rect 1152 5968 19654 6020
rect 19706 5968 19718 6020
rect 19770 5968 19782 6020
rect 19834 5968 19846 6020
rect 19898 5968 50374 6020
rect 50426 5968 50438 6020
rect 50490 5968 50502 6020
rect 50554 5968 50566 6020
rect 50618 5968 58848 6020
rect 1152 5946 58848 5968
rect 5104 5783 5110 5835
rect 5162 5823 5168 5835
rect 42736 5823 42742 5835
rect 5162 5795 42742 5823
rect 5162 5783 5168 5795
rect 42736 5783 42742 5795
rect 42794 5783 42800 5835
rect 57040 5783 57046 5835
rect 57098 5823 57104 5835
rect 57712 5823 57718 5835
rect 57098 5795 57718 5823
rect 57098 5783 57104 5795
rect 57712 5783 57718 5795
rect 57770 5783 57776 5835
rect 12115 5752 12173 5758
rect 12115 5718 12127 5752
rect 12161 5749 12173 5752
rect 15952 5749 15958 5761
rect 12161 5721 15958 5749
rect 12161 5718 12173 5721
rect 12115 5712 12173 5718
rect 15952 5709 15958 5721
rect 16010 5709 16016 5761
rect 21616 5709 21622 5761
rect 21674 5749 21680 5761
rect 21674 5721 22526 5749
rect 21674 5709 21680 5721
rect 1072 5635 1078 5687
rect 1130 5675 1136 5687
rect 1555 5678 1613 5684
rect 1555 5675 1567 5678
rect 1130 5647 1567 5675
rect 1130 5635 1136 5647
rect 1555 5644 1567 5647
rect 1601 5644 1613 5678
rect 1555 5638 1613 5644
rect 2896 5635 2902 5687
rect 2954 5675 2960 5687
rect 4435 5678 4493 5684
rect 2954 5647 2999 5675
rect 2954 5635 2960 5647
rect 4435 5644 4447 5678
rect 4481 5675 4493 5678
rect 4912 5675 4918 5687
rect 4481 5647 4918 5675
rect 4481 5644 4493 5647
rect 4435 5638 4493 5644
rect 4912 5635 4918 5647
rect 4970 5635 4976 5687
rect 5200 5675 5206 5687
rect 5161 5647 5206 5675
rect 5200 5635 5206 5647
rect 5258 5635 5264 5687
rect 6832 5675 6838 5687
rect 6793 5647 6838 5675
rect 6832 5635 6838 5647
rect 6890 5635 6896 5687
rect 7216 5635 7222 5687
rect 7274 5675 7280 5687
rect 7603 5678 7661 5684
rect 7603 5675 7615 5678
rect 7274 5647 7615 5675
rect 7274 5635 7280 5647
rect 7603 5644 7615 5647
rect 7649 5644 7661 5678
rect 7603 5638 7661 5644
rect 7987 5678 8045 5684
rect 7987 5644 7999 5678
rect 8033 5675 8045 5678
rect 8371 5678 8429 5684
rect 8371 5675 8383 5678
rect 8033 5647 8383 5675
rect 8033 5644 8045 5647
rect 7987 5638 8045 5644
rect 8371 5644 8383 5647
rect 8417 5644 8429 5678
rect 8371 5638 8429 5644
rect 8752 5635 8758 5687
rect 8810 5675 8816 5687
rect 9619 5678 9677 5684
rect 9619 5675 9631 5678
rect 8810 5647 9631 5675
rect 8810 5635 8816 5647
rect 9619 5644 9631 5647
rect 9665 5644 9677 5678
rect 9619 5638 9677 5644
rect 10192 5635 10198 5687
rect 10250 5675 10256 5687
rect 10387 5678 10445 5684
rect 10387 5675 10399 5678
rect 10250 5647 10399 5675
rect 10250 5635 10256 5647
rect 10387 5644 10399 5647
rect 10433 5644 10445 5678
rect 10387 5638 10445 5644
rect 10480 5635 10486 5687
rect 10538 5675 10544 5687
rect 11155 5678 11213 5684
rect 11155 5675 11167 5678
rect 10538 5647 11167 5675
rect 10538 5635 10544 5647
rect 11155 5644 11167 5647
rect 11201 5644 11213 5678
rect 12592 5675 12598 5687
rect 12553 5647 12598 5675
rect 11155 5638 11213 5644
rect 12592 5635 12598 5647
rect 12650 5635 12656 5687
rect 13459 5678 13517 5684
rect 13459 5644 13471 5678
rect 13505 5675 13517 5678
rect 13648 5675 13654 5687
rect 13505 5647 13654 5675
rect 13505 5644 13517 5647
rect 13459 5638 13517 5644
rect 13648 5635 13654 5647
rect 13706 5635 13712 5687
rect 14992 5675 14998 5687
rect 14953 5647 14998 5675
rect 14992 5635 14998 5647
rect 15050 5635 15056 5687
rect 15856 5675 15862 5687
rect 15817 5647 15862 5675
rect 15856 5635 15862 5647
rect 15914 5635 15920 5687
rect 16144 5635 16150 5687
rect 16202 5675 16208 5687
rect 16531 5678 16589 5684
rect 16531 5675 16543 5678
rect 16202 5647 16543 5675
rect 16202 5635 16208 5647
rect 16531 5644 16543 5647
rect 16577 5644 16589 5678
rect 16531 5638 16589 5644
rect 17296 5635 17302 5687
rect 17354 5675 17360 5687
rect 18736 5675 18742 5687
rect 17354 5647 17399 5675
rect 18697 5647 18742 5675
rect 17354 5635 17360 5647
rect 18736 5635 18742 5647
rect 18794 5635 18800 5687
rect 20176 5675 20182 5687
rect 20137 5647 20182 5675
rect 20176 5635 20182 5647
rect 20234 5635 20240 5687
rect 20560 5635 20566 5687
rect 20618 5675 20624 5687
rect 20947 5678 21005 5684
rect 20947 5675 20959 5678
rect 20618 5647 20959 5675
rect 20618 5635 20624 5647
rect 20947 5644 20959 5647
rect 20993 5644 21005 5678
rect 21712 5675 21718 5687
rect 21673 5647 21718 5675
rect 20947 5638 21005 5644
rect 21712 5635 21718 5647
rect 21770 5635 21776 5687
rect 22498 5684 22526 5721
rect 26032 5709 26038 5761
rect 26090 5749 26096 5761
rect 26090 5721 27038 5749
rect 26090 5709 26096 5721
rect 22483 5678 22541 5684
rect 22483 5644 22495 5678
rect 22529 5644 22541 5678
rect 22483 5638 22541 5644
rect 23152 5635 23158 5687
rect 23210 5675 23216 5687
rect 23251 5678 23309 5684
rect 23251 5675 23263 5678
rect 23210 5647 23263 5675
rect 23210 5635 23216 5647
rect 23251 5644 23263 5647
rect 23297 5644 23309 5678
rect 23251 5638 23309 5644
rect 23440 5635 23446 5687
rect 23498 5675 23504 5687
rect 24019 5678 24077 5684
rect 24019 5675 24031 5678
rect 23498 5647 24031 5675
rect 23498 5635 23504 5647
rect 24019 5644 24031 5647
rect 24065 5644 24077 5678
rect 24019 5638 24077 5644
rect 24592 5635 24598 5687
rect 24650 5675 24656 5687
rect 25459 5678 25517 5684
rect 25459 5675 25471 5678
rect 24650 5647 25471 5675
rect 24650 5635 24656 5647
rect 25459 5644 25471 5647
rect 25505 5644 25517 5678
rect 26224 5675 26230 5687
rect 26185 5647 26230 5675
rect 25459 5638 25517 5644
rect 26224 5635 26230 5647
rect 26282 5635 26288 5687
rect 27010 5684 27038 5721
rect 37456 5709 37462 5761
rect 37514 5749 37520 5761
rect 37514 5721 38366 5749
rect 37514 5709 37520 5721
rect 26995 5678 27053 5684
rect 26995 5644 27007 5678
rect 27041 5644 27053 5678
rect 26995 5638 27053 5644
rect 27376 5635 27382 5687
rect 27434 5675 27440 5687
rect 27763 5678 27821 5684
rect 27763 5675 27775 5678
rect 27434 5647 27775 5675
rect 27434 5635 27440 5647
rect 27763 5644 27775 5647
rect 27809 5644 27821 5678
rect 27763 5638 27821 5644
rect 27856 5635 27862 5687
rect 27914 5675 27920 5687
rect 28531 5678 28589 5684
rect 28531 5675 28543 5678
rect 27914 5647 28543 5675
rect 27914 5635 27920 5647
rect 28531 5644 28543 5647
rect 28577 5644 28589 5678
rect 28531 5638 28589 5644
rect 28816 5635 28822 5687
rect 28874 5675 28880 5687
rect 29299 5678 29357 5684
rect 29299 5675 29311 5678
rect 28874 5647 29311 5675
rect 28874 5635 28880 5647
rect 29299 5644 29311 5647
rect 29345 5644 29357 5678
rect 29299 5638 29357 5644
rect 30256 5635 30262 5687
rect 30314 5675 30320 5687
rect 30739 5678 30797 5684
rect 30739 5675 30751 5678
rect 30314 5647 30751 5675
rect 30314 5635 30320 5647
rect 30739 5644 30751 5647
rect 30785 5644 30797 5678
rect 30739 5638 30797 5644
rect 30832 5635 30838 5687
rect 30890 5675 30896 5687
rect 31507 5678 31565 5684
rect 31507 5675 31519 5678
rect 30890 5647 31519 5675
rect 30890 5635 30896 5647
rect 31507 5644 31519 5647
rect 31553 5644 31565 5678
rect 31507 5638 31565 5644
rect 31696 5635 31702 5687
rect 31754 5675 31760 5687
rect 32275 5678 32333 5684
rect 32275 5675 32287 5678
rect 31754 5647 32287 5675
rect 31754 5635 31760 5647
rect 32275 5644 32287 5647
rect 32321 5644 32333 5678
rect 33136 5675 33142 5687
rect 33097 5647 33142 5675
rect 32275 5638 32333 5644
rect 33136 5635 33142 5647
rect 33194 5635 33200 5687
rect 33232 5635 33238 5687
rect 33290 5675 33296 5687
rect 33811 5678 33869 5684
rect 33811 5675 33823 5678
rect 33290 5647 33823 5675
rect 33290 5635 33296 5647
rect 33811 5644 33823 5647
rect 33857 5644 33869 5678
rect 33811 5638 33869 5644
rect 34675 5678 34733 5684
rect 34675 5644 34687 5678
rect 34721 5675 34733 5678
rect 34768 5675 34774 5687
rect 34721 5647 34774 5675
rect 34721 5644 34733 5647
rect 34675 5638 34733 5644
rect 34768 5635 34774 5647
rect 34826 5635 34832 5687
rect 36112 5675 36118 5687
rect 36073 5647 36118 5675
rect 36112 5635 36118 5647
rect 36170 5635 36176 5687
rect 36208 5635 36214 5687
rect 36266 5675 36272 5687
rect 36787 5678 36845 5684
rect 36787 5675 36799 5678
rect 36266 5647 36799 5675
rect 36266 5635 36272 5647
rect 36787 5644 36799 5647
rect 36833 5644 36845 5678
rect 37552 5675 37558 5687
rect 37513 5647 37558 5675
rect 36787 5638 36845 5644
rect 37552 5635 37558 5647
rect 37610 5635 37616 5687
rect 38338 5684 38366 5721
rect 38323 5678 38381 5684
rect 38323 5644 38335 5678
rect 38369 5644 38381 5678
rect 39088 5675 39094 5687
rect 39049 5647 39094 5675
rect 38323 5638 38381 5644
rect 39088 5635 39094 5647
rect 39146 5635 39152 5687
rect 39280 5635 39286 5687
rect 39338 5675 39344 5687
rect 39859 5678 39917 5684
rect 39859 5675 39871 5678
rect 39338 5647 39871 5675
rect 39338 5635 39344 5647
rect 39859 5644 39871 5647
rect 39905 5644 39917 5678
rect 39859 5638 39917 5644
rect 40720 5635 40726 5687
rect 40778 5675 40784 5687
rect 41299 5678 41357 5684
rect 41299 5675 41311 5678
rect 40778 5647 41311 5675
rect 40778 5635 40784 5647
rect 41299 5644 41311 5647
rect 41345 5644 41357 5678
rect 41299 5638 41357 5644
rect 41776 5635 41782 5687
rect 41834 5675 41840 5687
rect 42067 5678 42125 5684
rect 42067 5675 42079 5678
rect 41834 5647 42079 5675
rect 41834 5635 41840 5647
rect 42067 5644 42079 5647
rect 42113 5644 42125 5678
rect 42067 5638 42125 5644
rect 42256 5635 42262 5687
rect 42314 5675 42320 5687
rect 42835 5678 42893 5684
rect 42835 5675 42847 5678
rect 42314 5647 42847 5675
rect 42314 5635 42320 5647
rect 42835 5644 42847 5647
rect 42881 5644 42893 5678
rect 42835 5638 42893 5644
rect 43216 5635 43222 5687
rect 43274 5675 43280 5687
rect 43603 5678 43661 5684
rect 43603 5675 43615 5678
rect 43274 5647 43615 5675
rect 43274 5635 43280 5647
rect 43603 5644 43615 5647
rect 43649 5644 43661 5678
rect 43603 5638 43661 5644
rect 43696 5635 43702 5687
rect 43754 5675 43760 5687
rect 44371 5678 44429 5684
rect 44371 5675 44383 5678
rect 43754 5647 44383 5675
rect 43754 5635 43760 5647
rect 44371 5644 44383 5647
rect 44417 5644 44429 5678
rect 45136 5675 45142 5687
rect 45097 5647 45142 5675
rect 44371 5638 44429 5644
rect 45136 5635 45142 5647
rect 45194 5635 45200 5687
rect 46096 5635 46102 5687
rect 46154 5675 46160 5687
rect 46579 5678 46637 5684
rect 46579 5675 46591 5678
rect 46154 5647 46591 5675
rect 46154 5635 46160 5647
rect 46579 5644 46591 5647
rect 46625 5644 46637 5678
rect 46579 5638 46637 5644
rect 46672 5635 46678 5687
rect 46730 5675 46736 5687
rect 47347 5678 47405 5684
rect 47347 5675 47359 5678
rect 46730 5647 47359 5675
rect 46730 5635 46736 5647
rect 47347 5644 47359 5647
rect 47393 5644 47405 5678
rect 47347 5638 47405 5644
rect 47536 5635 47542 5687
rect 47594 5675 47600 5687
rect 48115 5678 48173 5684
rect 48115 5675 48127 5678
rect 47594 5647 48127 5675
rect 47594 5635 47600 5647
rect 48115 5644 48127 5647
rect 48161 5644 48173 5678
rect 48115 5638 48173 5644
rect 48979 5678 49037 5684
rect 48979 5644 48991 5678
rect 49025 5675 49037 5678
rect 49072 5675 49078 5687
rect 49025 5647 49078 5675
rect 49025 5644 49037 5647
rect 48979 5638 49037 5644
rect 49072 5635 49078 5647
rect 49130 5635 49136 5687
rect 49648 5675 49654 5687
rect 49609 5647 49654 5675
rect 49648 5635 49654 5647
rect 49706 5635 49712 5687
rect 50515 5678 50573 5684
rect 50515 5644 50527 5678
rect 50561 5675 50573 5678
rect 50704 5675 50710 5687
rect 50561 5647 50710 5675
rect 50561 5644 50573 5647
rect 50515 5638 50573 5644
rect 50704 5635 50710 5647
rect 50762 5635 50768 5687
rect 52144 5675 52150 5687
rect 52105 5647 52150 5675
rect 52144 5635 52150 5647
rect 52202 5635 52208 5687
rect 52528 5635 52534 5687
rect 52586 5675 52592 5687
rect 52915 5678 52973 5684
rect 52915 5675 52927 5678
rect 52586 5647 52927 5675
rect 52586 5635 52592 5647
rect 52915 5644 52927 5647
rect 52961 5644 52973 5678
rect 53680 5675 53686 5687
rect 53641 5647 53686 5675
rect 52915 5638 52973 5644
rect 53680 5635 53686 5647
rect 53738 5635 53744 5687
rect 54451 5678 54509 5684
rect 54451 5644 54463 5678
rect 54497 5644 54509 5678
rect 54451 5638 54509 5644
rect 55987 5678 56045 5684
rect 55987 5644 55999 5678
rect 56033 5644 56045 5678
rect 57424 5675 57430 5687
rect 57385 5647 57430 5675
rect 55987 5638 56045 5644
rect 5968 5601 5974 5613
rect 5929 5573 5974 5601
rect 5968 5561 5974 5573
rect 6026 5561 6032 5613
rect 6067 5604 6125 5610
rect 6067 5570 6079 5604
rect 6113 5601 6125 5604
rect 50800 5601 50806 5613
rect 6113 5573 50806 5601
rect 6113 5570 6125 5573
rect 6067 5564 6125 5570
rect 50800 5561 50806 5573
rect 50858 5561 50864 5613
rect 53584 5561 53590 5613
rect 53642 5601 53648 5613
rect 54466 5601 54494 5638
rect 53642 5573 54494 5601
rect 56002 5601 56030 5638
rect 57424 5635 57430 5647
rect 57482 5635 57488 5687
rect 59632 5601 59638 5613
rect 56002 5573 59638 5601
rect 53642 5561 53648 5573
rect 59632 5561 59638 5573
rect 59690 5561 59696 5613
rect 7600 5487 7606 5539
rect 7658 5527 7664 5539
rect 7987 5530 8045 5536
rect 7987 5527 7999 5530
rect 7658 5499 7999 5527
rect 7658 5487 7664 5499
rect 7987 5496 7999 5499
rect 8033 5496 8045 5530
rect 7987 5490 8045 5496
rect 17584 5413 17590 5465
rect 17642 5453 17648 5465
rect 17872 5453 17878 5465
rect 17642 5425 17878 5453
rect 17642 5413 17648 5425
rect 17872 5413 17878 5425
rect 17930 5413 17936 5465
rect 17971 5456 18029 5462
rect 17971 5422 17983 5456
rect 18017 5453 18029 5456
rect 18259 5456 18317 5462
rect 18259 5453 18271 5456
rect 18017 5425 18271 5453
rect 18017 5422 18029 5425
rect 17971 5416 18029 5422
rect 18259 5422 18271 5425
rect 18305 5453 18317 5456
rect 29488 5453 29494 5465
rect 18305 5425 29494 5453
rect 18305 5422 18317 5425
rect 18259 5416 18317 5422
rect 29488 5413 29494 5425
rect 29546 5413 29552 5465
rect 33520 5413 33526 5465
rect 33578 5453 33584 5465
rect 55411 5456 55469 5462
rect 55411 5453 55423 5456
rect 33578 5425 55423 5453
rect 33578 5413 33584 5425
rect 55411 5422 55423 5425
rect 55457 5422 55469 5456
rect 55411 5416 55469 5422
rect 1152 5354 58848 5376
rect 1152 5302 4294 5354
rect 4346 5302 4358 5354
rect 4410 5302 4422 5354
rect 4474 5302 4486 5354
rect 4538 5302 35014 5354
rect 35066 5302 35078 5354
rect 35130 5302 35142 5354
rect 35194 5302 35206 5354
rect 35258 5302 58848 5354
rect 1152 5280 58848 5302
rect 7120 5191 7126 5243
rect 7178 5231 7184 5243
rect 38128 5231 38134 5243
rect 7178 5203 38134 5231
rect 7178 5191 7184 5203
rect 38128 5191 38134 5203
rect 38186 5191 38192 5243
rect 4720 5117 4726 5169
rect 4778 5157 4784 5169
rect 7507 5160 7565 5166
rect 7507 5157 7519 5160
rect 4778 5129 7519 5157
rect 4778 5117 4784 5129
rect 7507 5126 7519 5129
rect 7553 5157 7565 5160
rect 7553 5129 8640 5157
rect 7553 5126 7565 5129
rect 7507 5120 7565 5126
rect 11056 5117 11062 5169
rect 11114 5157 11120 5169
rect 20464 5157 20470 5169
rect 11114 5129 20470 5157
rect 11114 5117 11120 5129
rect 20464 5117 20470 5129
rect 20522 5117 20528 5169
rect 3568 5043 3574 5095
rect 3626 5083 3632 5095
rect 3626 5055 7968 5083
rect 3626 5043 3632 5055
rect 304 4969 310 5021
rect 362 5009 368 5021
rect 1555 5012 1613 5018
rect 1555 5009 1567 5012
rect 362 4981 1567 5009
rect 362 4969 368 4981
rect 1555 4978 1567 4981
rect 1601 4978 1613 5012
rect 1555 4972 1613 4978
rect 1840 4969 1846 5021
rect 1898 5009 1904 5021
rect 2323 5012 2381 5018
rect 2323 5009 2335 5012
rect 1898 4981 2335 5009
rect 1898 4969 1904 4981
rect 2323 4978 2335 4981
rect 2369 4978 2381 5012
rect 3088 5009 3094 5021
rect 3049 4981 3094 5009
rect 2323 4972 2381 4978
rect 3088 4969 3094 4981
rect 3146 4969 3152 5021
rect 4144 5009 4150 5021
rect 4105 4981 4150 5009
rect 4144 4969 4150 4981
rect 4202 4969 4208 5021
rect 5392 5009 5398 5021
rect 5353 4981 5398 5009
rect 5392 4969 5398 4981
rect 5450 4969 5456 5021
rect 6064 4969 6070 5021
rect 6122 5009 6128 5021
rect 6931 5012 6989 5018
rect 6931 5009 6943 5012
rect 6122 4981 6943 5009
rect 6122 4969 6128 4981
rect 6931 4978 6943 4981
rect 6977 4978 6989 5012
rect 9232 5009 9238 5021
rect 9193 4981 9238 5009
rect 6931 4972 6989 4978
rect 9232 4969 9238 4981
rect 9290 4969 9296 5021
rect 10099 5012 10157 5018
rect 10099 4978 10111 5012
rect 10145 5009 10157 5012
rect 10576 5009 10582 5021
rect 10145 4981 10582 5009
rect 10145 4978 10157 4981
rect 10099 4972 10157 4978
rect 10576 4969 10582 4981
rect 10634 4969 10640 5021
rect 10867 5012 10925 5018
rect 10867 4978 10879 5012
rect 10913 5009 10925 5012
rect 11056 5009 11062 5021
rect 10913 4981 11062 5009
rect 10913 4978 10925 4981
rect 10867 4972 10925 4978
rect 11056 4969 11062 4981
rect 11114 4969 11120 5021
rect 11824 4969 11830 5021
rect 11882 5009 11888 5021
rect 12211 5012 12269 5018
rect 12211 5009 12223 5012
rect 11882 4981 12223 5009
rect 11882 4969 11888 4981
rect 12211 4978 12223 4981
rect 12257 4978 12269 5012
rect 12976 5009 12982 5021
rect 12937 4981 12982 5009
rect 12211 4972 12269 4978
rect 12976 4969 12982 4981
rect 13034 4969 13040 5021
rect 13936 5009 13942 5021
rect 13897 4981 13942 5009
rect 13936 4969 13942 4981
rect 13994 4969 14000 5021
rect 14416 4969 14422 5021
rect 14474 5009 14480 5021
rect 14707 5012 14765 5018
rect 14707 5009 14719 5012
rect 14474 4981 14719 5009
rect 14474 4969 14480 4981
rect 14707 4978 14719 4981
rect 14753 4978 14765 5012
rect 14707 4972 14765 4978
rect 14800 4969 14806 5021
rect 14858 5009 14864 5021
rect 15475 5012 15533 5018
rect 15475 5009 15487 5012
rect 14858 4981 15487 5009
rect 14858 4969 14864 4981
rect 15475 4978 15487 4981
rect 15521 4978 15533 5012
rect 15475 4972 15533 4978
rect 16339 5012 16397 5018
rect 16339 4978 16351 5012
rect 16385 5009 16397 5012
rect 16432 5009 16438 5021
rect 16385 4981 16438 5009
rect 16385 4978 16397 4981
rect 16339 4972 16397 4978
rect 16432 4969 16438 4981
rect 16490 4969 16496 5021
rect 17488 5009 17494 5021
rect 17449 4981 17494 5009
rect 17488 4969 17494 4981
rect 17546 4969 17552 5021
rect 18256 5009 18262 5021
rect 18217 4981 18262 5009
rect 18256 4969 18262 4981
rect 18314 4969 18320 5021
rect 19024 5009 19030 5021
rect 18985 4981 19030 5009
rect 19024 4969 19030 4981
rect 19082 4969 19088 5021
rect 19120 4969 19126 5021
rect 19178 5009 19184 5021
rect 19795 5012 19853 5018
rect 19795 5009 19807 5012
rect 19178 4981 19807 5009
rect 19178 4969 19184 4981
rect 19795 4978 19807 4981
rect 19841 4978 19853 5012
rect 20656 5009 20662 5021
rect 20617 4981 20662 5009
rect 19795 4972 19853 4978
rect 20656 4969 20662 4981
rect 20714 4969 20720 5021
rect 20848 4969 20854 5021
rect 20906 5009 20912 5021
rect 21331 5012 21389 5018
rect 21331 5009 21343 5012
rect 20906 4981 21343 5009
rect 20906 4969 20912 4981
rect 21331 4978 21343 4981
rect 21377 4978 21389 5012
rect 22768 5009 22774 5021
rect 22729 4981 22774 5009
rect 21331 4972 21389 4978
rect 22768 4969 22774 4981
rect 22826 4969 22832 5021
rect 23536 5009 23542 5021
rect 23497 4981 23542 5009
rect 23536 4969 23542 4981
rect 23594 4969 23600 5021
rect 24307 5012 24365 5018
rect 24307 4978 24319 5012
rect 24353 4978 24365 5012
rect 25072 5009 25078 5021
rect 25033 4981 25078 5009
rect 24307 4972 24365 4978
rect 23056 4895 23062 4947
rect 23114 4935 23120 4947
rect 24322 4935 24350 4972
rect 25072 4969 25078 4981
rect 25130 4969 25136 5021
rect 25840 5009 25846 5021
rect 25801 4981 25846 5009
rect 25840 4969 25846 4981
rect 25898 4969 25904 5021
rect 26608 5009 26614 5021
rect 26569 4981 26614 5009
rect 26608 4969 26614 4981
rect 26666 4969 26672 5021
rect 28048 5009 28054 5021
rect 28009 4981 28054 5009
rect 28048 4969 28054 4981
rect 28106 4969 28112 5021
rect 28912 5009 28918 5021
rect 28873 4981 28918 5009
rect 28912 4969 28918 4981
rect 28970 4969 28976 5021
rect 29296 4969 29302 5021
rect 29354 5009 29360 5021
rect 29587 5012 29645 5018
rect 29587 5009 29599 5012
rect 29354 4981 29599 5009
rect 29354 4969 29360 4981
rect 29587 4978 29599 4981
rect 29633 4978 29645 5012
rect 30352 5009 30358 5021
rect 30313 4981 30358 5009
rect 29587 4972 29645 4978
rect 30352 4969 30358 4981
rect 30410 4969 30416 5021
rect 30448 4969 30454 5021
rect 30506 5009 30512 5021
rect 31123 5012 31181 5018
rect 31123 5009 31135 5012
rect 30506 4981 31135 5009
rect 30506 4969 30512 4981
rect 31123 4978 31135 4981
rect 31169 4978 31181 5012
rect 31888 5009 31894 5021
rect 31849 4981 31894 5009
rect 31123 4972 31181 4978
rect 31888 4969 31894 4981
rect 31946 4969 31952 5021
rect 33328 5009 33334 5021
rect 33289 4981 33334 5009
rect 33328 4969 33334 4981
rect 33386 4969 33392 5021
rect 34096 5009 34102 5021
rect 34057 4981 34102 5009
rect 34096 4969 34102 4981
rect 34154 4969 34160 5021
rect 34864 5009 34870 5021
rect 34825 4981 34870 5009
rect 34864 4969 34870 4981
rect 34922 4969 34928 5021
rect 35635 5012 35693 5018
rect 35635 4978 35647 5012
rect 35681 4978 35693 5012
rect 36400 5009 36406 5021
rect 36361 4981 36406 5009
rect 35635 4972 35693 4978
rect 23114 4907 24350 4935
rect 23114 4895 23120 4907
rect 34576 4895 34582 4947
rect 34634 4935 34640 4947
rect 35650 4935 35678 4972
rect 36400 4969 36406 4981
rect 36458 4969 36464 5021
rect 36688 4969 36694 5021
rect 36746 5009 36752 5021
rect 37171 5012 37229 5018
rect 37171 5009 37183 5012
rect 36746 4981 37183 5009
rect 36746 4969 36752 4981
rect 37171 4978 37183 4981
rect 37217 4978 37229 5012
rect 38608 5009 38614 5021
rect 38569 4981 38614 5009
rect 37171 4972 37229 4978
rect 38608 4969 38614 4981
rect 38666 4969 38672 5021
rect 39376 5009 39382 5021
rect 39337 4981 39382 5009
rect 39376 4969 39382 4981
rect 39434 4969 39440 5021
rect 40144 5009 40150 5021
rect 40105 4981 40150 5009
rect 40144 4969 40150 4981
rect 40202 4969 40208 5021
rect 40912 5009 40918 5021
rect 40873 4981 40918 5009
rect 40912 4969 40918 4981
rect 40970 4969 40976 5021
rect 41680 5009 41686 5021
rect 41641 4981 41686 5009
rect 41680 4969 41686 4981
rect 41738 4969 41744 5021
rect 42064 4969 42070 5021
rect 42122 5009 42128 5021
rect 42451 5012 42509 5018
rect 42451 5009 42463 5012
rect 42122 4981 42463 5009
rect 42122 4969 42128 4981
rect 42451 4978 42463 4981
rect 42497 4978 42509 5012
rect 42451 4972 42509 4978
rect 43504 4969 43510 5021
rect 43562 5009 43568 5021
rect 43891 5012 43949 5018
rect 43891 5009 43903 5012
rect 43562 4981 43903 5009
rect 43562 4969 43568 4981
rect 43891 4978 43903 4981
rect 43937 4978 43949 5012
rect 44752 5009 44758 5021
rect 44713 4981 44758 5009
rect 43891 4972 43949 4978
rect 44752 4969 44758 4981
rect 44810 4969 44816 5021
rect 45424 5009 45430 5021
rect 45385 4981 45430 5009
rect 45424 4969 45430 4981
rect 45482 4969 45488 5021
rect 46192 5009 46198 5021
rect 46153 4981 46198 5009
rect 46192 4969 46198 4981
rect 46250 4969 46256 5021
rect 46288 4969 46294 5021
rect 46346 5009 46352 5021
rect 46963 5012 47021 5018
rect 46963 5009 46975 5012
rect 46346 4981 46975 5009
rect 46346 4969 46352 4981
rect 46963 4978 46975 4981
rect 47009 4978 47021 5012
rect 46963 4972 47021 4978
rect 47632 4969 47638 5021
rect 47690 5009 47696 5021
rect 47731 5012 47789 5018
rect 47731 5009 47743 5012
rect 47690 4981 47743 5009
rect 47690 4969 47696 4981
rect 47731 4978 47743 4981
rect 47777 4978 47789 5012
rect 49360 5009 49366 5021
rect 49321 4981 49366 5009
rect 47731 4972 47789 4978
rect 49360 4969 49366 4981
rect 49418 4969 49424 5021
rect 50416 5009 50422 5021
rect 50377 4981 50422 5009
rect 50416 4969 50422 4981
rect 50474 4969 50480 5021
rect 50896 4969 50902 5021
rect 50954 5009 50960 5021
rect 51091 5012 51149 5018
rect 51091 5009 51103 5012
rect 50954 4981 51103 5009
rect 50954 4969 50960 4981
rect 51091 4978 51103 4981
rect 51137 4978 51149 5012
rect 51856 5009 51862 5021
rect 51817 4981 51862 5009
rect 51091 4972 51149 4978
rect 51856 4969 51862 4981
rect 51914 4969 51920 5021
rect 51952 4969 51958 5021
rect 52010 5009 52016 5021
rect 52627 5012 52685 5018
rect 52627 5009 52639 5012
rect 52010 4981 52639 5009
rect 52010 4969 52016 4981
rect 52627 4978 52639 4981
rect 52673 4978 52685 5012
rect 52627 4972 52685 4978
rect 53296 4969 53302 5021
rect 53354 5009 53360 5021
rect 54451 5012 54509 5018
rect 54451 5009 54463 5012
rect 53354 4981 54463 5009
rect 53354 4969 53360 4981
rect 54451 4978 54463 4981
rect 54497 4978 54509 5012
rect 54451 4972 54509 4978
rect 55603 5012 55661 5018
rect 55603 4978 55615 5012
rect 55649 4978 55661 5012
rect 55603 4972 55661 4978
rect 56371 5012 56429 5018
rect 56371 4978 56383 5012
rect 56417 4978 56429 5012
rect 57040 5009 57046 5021
rect 57001 4981 57046 5009
rect 56371 4972 56429 4978
rect 34634 4907 35678 4935
rect 34634 4895 34640 4907
rect 55618 4861 55646 4972
rect 56386 4935 56414 4972
rect 57040 4969 57046 4981
rect 57098 4969 57104 5021
rect 57808 4935 57814 4947
rect 56386 4907 57814 4935
rect 57808 4895 57814 4907
rect 57866 4895 57872 4947
rect 59248 4861 59254 4873
rect 2866 4833 7646 4861
rect 2128 4747 2134 4799
rect 2186 4787 2192 4799
rect 2866 4787 2894 4833
rect 2186 4759 2894 4787
rect 7618 4787 7646 4833
rect 8242 4787 8270 4847
rect 55618 4833 59254 4861
rect 59248 4821 59254 4833
rect 59306 4821 59312 4873
rect 7618 4759 8270 4787
rect 2186 4747 2192 4759
rect 1152 4688 58848 4710
rect 1152 4636 19654 4688
rect 19706 4636 19718 4688
rect 19770 4636 19782 4688
rect 19834 4636 19846 4688
rect 19898 4636 50374 4688
rect 50426 4636 50438 4688
rect 50490 4636 50502 4688
rect 50554 4636 50566 4688
rect 50618 4636 58848 4688
rect 1152 4614 58848 4636
rect 11152 4525 11158 4577
rect 11210 4565 11216 4577
rect 15763 4568 15821 4574
rect 15763 4565 15775 4568
rect 11210 4537 15775 4565
rect 11210 4525 11216 4537
rect 15763 4534 15775 4537
rect 15809 4534 15821 4568
rect 15763 4528 15821 4534
rect 20464 4525 20470 4577
rect 20522 4565 20528 4577
rect 20563 4568 20621 4574
rect 20563 4565 20575 4568
rect 20522 4537 20575 4565
rect 20522 4525 20528 4537
rect 20563 4534 20575 4537
rect 20609 4534 20621 4568
rect 38128 4565 38134 4577
rect 38089 4537 38134 4565
rect 20563 4528 20621 4534
rect 38128 4525 38134 4537
rect 38186 4525 38192 4577
rect 54835 4568 54893 4574
rect 54835 4534 54847 4568
rect 54881 4565 54893 4568
rect 55123 4568 55181 4574
rect 55123 4565 55135 4568
rect 54881 4537 55135 4565
rect 54881 4534 54893 4537
rect 54835 4528 54893 4534
rect 55123 4534 55135 4537
rect 55169 4565 55181 4568
rect 57328 4565 57334 4577
rect 55169 4537 57334 4565
rect 55169 4534 55181 4537
rect 55123 4528 55181 4534
rect 57328 4525 57334 4537
rect 57386 4525 57392 4577
rect 10768 4451 10774 4503
rect 10826 4451 10832 4503
rect 11440 4451 11446 4503
rect 11498 4491 11504 4503
rect 16531 4494 16589 4500
rect 16531 4491 16543 4494
rect 11498 4463 16543 4491
rect 11498 4451 11504 4463
rect 16531 4460 16543 4463
rect 16577 4460 16589 4494
rect 16531 4454 16589 4460
rect 17299 4494 17357 4500
rect 17299 4460 17311 4494
rect 17345 4460 17357 4494
rect 17299 4454 17357 4460
rect 784 4377 790 4429
rect 842 4417 848 4429
rect 10786 4417 10814 4451
rect 17314 4417 17342 4454
rect 842 4389 2366 4417
rect 10786 4389 17342 4417
rect 38146 4417 38174 4525
rect 38323 4420 38381 4426
rect 38323 4417 38335 4420
rect 38146 4389 38335 4417
rect 842 4377 848 4389
rect 1168 4303 1174 4355
rect 1226 4343 1232 4355
rect 2338 4352 2366 4389
rect 38323 4386 38335 4389
rect 38369 4386 38381 4420
rect 38323 4380 38381 4386
rect 1555 4346 1613 4352
rect 1555 4343 1567 4346
rect 1226 4315 1567 4343
rect 1226 4303 1232 4315
rect 1555 4312 1567 4315
rect 1601 4312 1613 4346
rect 1555 4306 1613 4312
rect 2323 4346 2381 4352
rect 2323 4312 2335 4346
rect 2369 4312 2381 4346
rect 3091 4346 3149 4352
rect 3091 4343 3103 4346
rect 2323 4306 2381 4312
rect 2866 4315 3103 4343
rect 1360 4229 1366 4281
rect 1418 4269 1424 4281
rect 2866 4269 2894 4315
rect 3091 4312 3103 4315
rect 3137 4312 3149 4346
rect 3091 4306 3149 4312
rect 4339 4346 4397 4352
rect 4339 4312 4351 4346
rect 4385 4312 4397 4346
rect 4339 4306 4397 4312
rect 1418 4241 2894 4269
rect 1418 4229 1424 4241
rect 3760 4229 3766 4281
rect 3818 4269 3824 4281
rect 4354 4269 4382 4306
rect 4720 4303 4726 4355
rect 4778 4343 4784 4355
rect 5107 4346 5165 4352
rect 5107 4343 5119 4346
rect 4778 4315 5119 4343
rect 4778 4303 4784 4315
rect 5107 4312 5119 4315
rect 5153 4312 5165 4346
rect 5875 4346 5933 4352
rect 5875 4343 5887 4346
rect 5107 4306 5165 4312
rect 5602 4315 5887 4343
rect 3818 4241 4382 4269
rect 3818 4229 3824 4241
rect 3472 4155 3478 4207
rect 3530 4195 3536 4207
rect 4912 4195 4918 4207
rect 3530 4167 4918 4195
rect 3530 4155 3536 4167
rect 4912 4155 4918 4167
rect 4970 4155 4976 4207
rect 5104 4155 5110 4207
rect 5162 4195 5168 4207
rect 5602 4195 5630 4315
rect 5875 4312 5887 4315
rect 5921 4312 5933 4346
rect 5875 4306 5933 4312
rect 6643 4346 6701 4352
rect 6643 4312 6655 4346
rect 6689 4312 6701 4346
rect 7408 4343 7414 4355
rect 7369 4315 7414 4343
rect 6643 4306 6701 4312
rect 5680 4229 5686 4281
rect 5738 4269 5744 4281
rect 6658 4269 6686 4306
rect 7408 4303 7414 4315
rect 7466 4303 7472 4355
rect 8179 4346 8237 4352
rect 8179 4312 8191 4346
rect 8225 4312 8237 4346
rect 9616 4343 9622 4355
rect 9577 4315 9622 4343
rect 8179 4306 8237 4312
rect 5738 4241 6686 4269
rect 5738 4229 5744 4241
rect 5162 4167 5630 4195
rect 5162 4155 5168 4167
rect 6448 4155 6454 4207
rect 6506 4195 6512 4207
rect 8194 4195 8222 4306
rect 9616 4303 9622 4315
rect 9674 4303 9680 4355
rect 10384 4343 10390 4355
rect 10345 4315 10390 4343
rect 10384 4303 10390 4315
rect 10442 4303 10448 4355
rect 10768 4303 10774 4355
rect 10826 4343 10832 4355
rect 11155 4346 11213 4352
rect 11155 4343 11167 4346
rect 10826 4315 11167 4343
rect 10826 4303 10832 4315
rect 11155 4312 11167 4315
rect 11201 4312 11213 4346
rect 11923 4346 11981 4352
rect 11923 4343 11935 4346
rect 11155 4306 11213 4312
rect 11266 4315 11935 4343
rect 9808 4229 9814 4281
rect 9866 4269 9872 4281
rect 10192 4269 10198 4281
rect 9866 4241 10198 4269
rect 9866 4229 9872 4241
rect 10192 4229 10198 4241
rect 10250 4229 10256 4281
rect 6506 4167 8222 4195
rect 6506 4155 6512 4167
rect 11152 4155 11158 4207
rect 11210 4195 11216 4207
rect 11266 4195 11294 4315
rect 11923 4312 11935 4315
rect 11969 4312 11981 4346
rect 11923 4306 11981 4312
rect 12691 4346 12749 4352
rect 12691 4312 12703 4346
rect 12737 4312 12749 4346
rect 13552 4343 13558 4355
rect 13513 4315 13558 4343
rect 12691 4306 12749 4312
rect 11440 4229 11446 4281
rect 11498 4269 11504 4281
rect 12706 4269 12734 4306
rect 13552 4303 13558 4315
rect 13610 4303 13616 4355
rect 15472 4343 15478 4355
rect 15433 4315 15478 4343
rect 15472 4303 15478 4315
rect 15530 4303 15536 4355
rect 15952 4303 15958 4355
rect 16010 4343 16016 4355
rect 16243 4346 16301 4352
rect 16243 4343 16255 4346
rect 16010 4315 16255 4343
rect 16010 4303 16016 4315
rect 16243 4312 16255 4315
rect 16289 4312 16301 4346
rect 16243 4306 16301 4312
rect 17011 4346 17069 4352
rect 17011 4312 17023 4346
rect 17057 4312 17069 4346
rect 17779 4346 17837 4352
rect 17779 4343 17791 4346
rect 17011 4306 17069 4312
rect 17266 4315 17791 4343
rect 11498 4241 12734 4269
rect 11498 4229 11504 4241
rect 11210 4167 11294 4195
rect 11210 4155 11216 4167
rect 16240 4155 16246 4207
rect 16298 4195 16304 4207
rect 17026 4195 17054 4306
rect 16298 4167 17054 4195
rect 16298 4155 16304 4167
rect 976 4081 982 4133
rect 1034 4121 1040 4133
rect 2320 4121 2326 4133
rect 1034 4093 2326 4121
rect 1034 4081 1040 4093
rect 2320 4081 2326 4093
rect 2378 4081 2384 4133
rect 2416 4081 2422 4133
rect 2474 4121 2480 4133
rect 5008 4121 5014 4133
rect 2474 4093 5014 4121
rect 2474 4081 2480 4093
rect 5008 4081 5014 4093
rect 5066 4081 5072 4133
rect 9040 4081 9046 4133
rect 9098 4121 9104 4133
rect 11056 4121 11062 4133
rect 9098 4093 11062 4121
rect 9098 4081 9104 4093
rect 11056 4081 11062 4093
rect 11114 4081 11120 4133
rect 16912 4081 16918 4133
rect 16970 4121 16976 4133
rect 17266 4121 17294 4315
rect 17779 4312 17791 4315
rect 17825 4312 17837 4346
rect 17779 4306 17837 4312
rect 18547 4346 18605 4352
rect 18547 4312 18559 4346
rect 18593 4312 18605 4346
rect 20272 4343 20278 4355
rect 20233 4315 20278 4343
rect 18547 4306 18605 4312
rect 17680 4229 17686 4281
rect 17738 4269 17744 4281
rect 18562 4269 18590 4306
rect 20272 4303 20278 4315
rect 20330 4303 20336 4355
rect 21040 4343 21046 4355
rect 21001 4315 21046 4343
rect 21040 4303 21046 4315
rect 21098 4303 21104 4355
rect 21808 4343 21814 4355
rect 21769 4315 21814 4343
rect 21808 4303 21814 4315
rect 21866 4303 21872 4355
rect 23248 4343 23254 4355
rect 23209 4315 23254 4343
rect 23248 4303 23254 4315
rect 23306 4303 23312 4355
rect 24019 4346 24077 4352
rect 24019 4312 24031 4346
rect 24065 4312 24077 4346
rect 25456 4343 25462 4355
rect 25417 4315 25462 4343
rect 24019 4306 24077 4312
rect 17738 4241 18590 4269
rect 17738 4229 17744 4241
rect 22000 4229 22006 4281
rect 22058 4269 22064 4281
rect 24034 4269 24062 4306
rect 25456 4303 25462 4315
rect 25514 4303 25520 4355
rect 26128 4303 26134 4355
rect 26186 4343 26192 4355
rect 26227 4346 26285 4352
rect 26227 4343 26239 4346
rect 26186 4315 26239 4343
rect 26186 4303 26192 4315
rect 26227 4312 26239 4315
rect 26273 4312 26285 4346
rect 26227 4306 26285 4312
rect 26512 4303 26518 4355
rect 26570 4343 26576 4355
rect 26995 4346 27053 4352
rect 26995 4343 27007 4346
rect 26570 4315 27007 4343
rect 26570 4303 26576 4315
rect 26995 4312 27007 4315
rect 27041 4312 27053 4346
rect 28336 4343 28342 4355
rect 28297 4315 28342 4343
rect 26995 4306 27053 4312
rect 28336 4303 28342 4315
rect 28394 4303 28400 4355
rect 29104 4343 29110 4355
rect 29065 4315 29110 4343
rect 29104 4303 29110 4315
rect 29162 4303 29168 4355
rect 30928 4343 30934 4355
rect 30889 4315 30934 4343
rect 30928 4303 30934 4315
rect 30986 4303 30992 4355
rect 31696 4343 31702 4355
rect 31657 4315 31702 4343
rect 31696 4303 31702 4315
rect 31754 4303 31760 4355
rect 32752 4343 32758 4355
rect 32713 4315 32758 4343
rect 32752 4303 32758 4315
rect 32810 4303 32816 4355
rect 33904 4343 33910 4355
rect 33865 4315 33910 4343
rect 33904 4303 33910 4315
rect 33962 4303 33968 4355
rect 34576 4303 34582 4355
rect 34634 4343 34640 4355
rect 34675 4346 34733 4352
rect 34675 4343 34687 4346
rect 34634 4315 34687 4343
rect 34634 4303 34640 4315
rect 34675 4312 34687 4315
rect 34721 4312 34733 4346
rect 36019 4346 36077 4352
rect 36019 4343 36031 4346
rect 34675 4306 34733 4312
rect 34786 4315 36031 4343
rect 22058 4241 24062 4269
rect 22058 4229 22064 4241
rect 34192 4229 34198 4281
rect 34250 4269 34256 4281
rect 34786 4269 34814 4315
rect 36019 4312 36031 4315
rect 36065 4312 36077 4346
rect 36784 4343 36790 4355
rect 36745 4315 36790 4343
rect 36019 4306 36077 4312
rect 36784 4303 36790 4315
rect 36842 4303 36848 4355
rect 37555 4346 37613 4352
rect 37555 4343 37567 4346
rect 37426 4315 37567 4343
rect 34250 4241 34814 4269
rect 34250 4229 34256 4241
rect 37168 4229 37174 4281
rect 37226 4269 37232 4281
rect 37426 4269 37454 4315
rect 37555 4312 37567 4315
rect 37601 4312 37613 4346
rect 38992 4343 38998 4355
rect 38953 4315 38998 4343
rect 37555 4306 37613 4312
rect 38992 4303 38998 4315
rect 39050 4303 39056 4355
rect 39760 4343 39766 4355
rect 39721 4315 39766 4343
rect 39760 4303 39766 4315
rect 39818 4303 39824 4355
rect 41968 4343 41974 4355
rect 41929 4315 41974 4343
rect 41968 4303 41974 4315
rect 42026 4303 42032 4355
rect 42352 4303 42358 4355
rect 42410 4343 42416 4355
rect 42739 4346 42797 4352
rect 42739 4343 42751 4346
rect 42410 4315 42751 4343
rect 42410 4303 42416 4315
rect 42739 4312 42751 4315
rect 42785 4312 42797 4346
rect 42739 4306 42797 4312
rect 43408 4303 43414 4355
rect 43466 4343 43472 4355
rect 43507 4346 43565 4352
rect 43507 4343 43519 4346
rect 43466 4315 43519 4343
rect 43466 4303 43472 4315
rect 43507 4312 43519 4315
rect 43553 4312 43565 4346
rect 44944 4343 44950 4355
rect 44905 4315 44950 4343
rect 43507 4306 43565 4312
rect 44944 4303 44950 4315
rect 45002 4303 45008 4355
rect 46768 4343 46774 4355
rect 46729 4315 46774 4343
rect 46768 4303 46774 4315
rect 46826 4303 46832 4355
rect 47539 4346 47597 4352
rect 47539 4312 47551 4346
rect 47585 4312 47597 4346
rect 47539 4306 47597 4312
rect 37226 4241 37454 4269
rect 37226 4229 37232 4241
rect 44464 4229 44470 4281
rect 44522 4269 44528 4281
rect 45136 4269 45142 4281
rect 44522 4241 45142 4269
rect 44522 4229 44528 4241
rect 45136 4229 45142 4241
rect 45194 4229 45200 4281
rect 47440 4229 47446 4281
rect 47498 4269 47504 4281
rect 47554 4269 47582 4306
rect 47824 4303 47830 4355
rect 47882 4343 47888 4355
rect 48307 4346 48365 4352
rect 48307 4343 48319 4346
rect 47882 4315 48319 4343
rect 47882 4303 47888 4315
rect 48307 4312 48319 4315
rect 48353 4312 48365 4346
rect 48307 4306 48365 4312
rect 49075 4346 49133 4352
rect 49075 4312 49087 4346
rect 49121 4312 49133 4346
rect 49075 4306 49133 4312
rect 49843 4346 49901 4352
rect 49843 4312 49855 4346
rect 49889 4312 49901 4346
rect 49843 4306 49901 4312
rect 50611 4346 50669 4352
rect 50611 4312 50623 4346
rect 50657 4312 50669 4346
rect 50611 4306 50669 4312
rect 51859 4346 51917 4352
rect 51859 4312 51871 4346
rect 51905 4312 51917 4346
rect 52624 4343 52630 4355
rect 52585 4315 52630 4343
rect 51859 4306 51917 4312
rect 47498 4241 47582 4269
rect 47498 4229 47504 4241
rect 48592 4229 48598 4281
rect 48650 4269 48656 4281
rect 49090 4269 49118 4306
rect 48650 4241 49118 4269
rect 48650 4229 48656 4241
rect 43792 4155 43798 4207
rect 43850 4195 43856 4207
rect 47152 4195 47158 4207
rect 43850 4167 47158 4195
rect 43850 4155 43856 4167
rect 47152 4155 47158 4167
rect 47210 4155 47216 4207
rect 48976 4155 48982 4207
rect 49034 4195 49040 4207
rect 49858 4195 49886 4306
rect 49936 4229 49942 4281
rect 49994 4269 50000 4281
rect 50626 4269 50654 4306
rect 49994 4241 50654 4269
rect 49994 4229 50000 4241
rect 50992 4229 50998 4281
rect 51050 4269 51056 4281
rect 51874 4269 51902 4306
rect 52624 4303 52630 4315
rect 52682 4303 52688 4355
rect 53395 4346 53453 4352
rect 53395 4343 53407 4346
rect 53266 4315 53407 4343
rect 51050 4241 51902 4269
rect 51050 4229 51056 4241
rect 53008 4229 53014 4281
rect 53066 4269 53072 4281
rect 53266 4269 53294 4315
rect 53395 4312 53407 4315
rect 53441 4312 53453 4346
rect 53395 4306 53453 4312
rect 54064 4303 54070 4355
rect 54122 4343 54128 4355
rect 54163 4346 54221 4352
rect 54163 4343 54175 4346
rect 54122 4315 54175 4343
rect 54122 4303 54128 4315
rect 54163 4312 54175 4315
rect 54209 4312 54221 4346
rect 55600 4343 55606 4355
rect 55561 4315 55606 4343
rect 54163 4306 54221 4312
rect 55600 4303 55606 4315
rect 55658 4303 55664 4355
rect 56656 4303 56662 4355
rect 56714 4343 56720 4355
rect 57139 4346 57197 4352
rect 57139 4343 57151 4346
rect 56714 4315 57151 4343
rect 56714 4303 56720 4315
rect 57139 4312 57151 4315
rect 57185 4312 57197 4346
rect 57139 4306 57197 4312
rect 53066 4241 53294 4269
rect 53066 4229 53072 4241
rect 56848 4229 56854 4281
rect 56906 4269 56912 4281
rect 59152 4269 59158 4281
rect 56906 4241 59158 4269
rect 56906 4229 56912 4241
rect 59152 4229 59158 4241
rect 59210 4229 59216 4281
rect 49034 4167 49886 4195
rect 49034 4155 49040 4167
rect 56368 4155 56374 4207
rect 56426 4195 56432 4207
rect 58288 4195 58294 4207
rect 56426 4167 58294 4195
rect 56426 4155 56432 4167
rect 58288 4155 58294 4167
rect 58346 4155 58352 4207
rect 16970 4093 17294 4121
rect 16970 4081 16976 4093
rect 17872 4081 17878 4133
rect 17930 4121 17936 4133
rect 20944 4121 20950 4133
rect 17930 4093 20950 4121
rect 17930 4081 17936 4093
rect 20944 4081 20950 4093
rect 21002 4081 21008 4133
rect 21520 4081 21526 4133
rect 21578 4121 21584 4133
rect 22864 4121 22870 4133
rect 21578 4093 22870 4121
rect 21578 4081 21584 4093
rect 22864 4081 22870 4093
rect 22922 4081 22928 4133
rect 24976 4081 24982 4133
rect 25034 4121 25040 4133
rect 26608 4121 26614 4133
rect 25034 4093 26614 4121
rect 25034 4081 25040 4093
rect 26608 4081 26614 4093
rect 26666 4081 26672 4133
rect 40048 4081 40054 4133
rect 40106 4121 40112 4133
rect 41680 4121 41686 4133
rect 40106 4093 41686 4121
rect 40106 4081 40112 4093
rect 41680 4081 41686 4093
rect 41738 4081 41744 4133
rect 45328 4081 45334 4133
rect 45386 4121 45392 4133
rect 46288 4121 46294 4133
rect 45386 4093 46294 4121
rect 45386 4081 45392 4093
rect 46288 4081 46294 4093
rect 46346 4081 46352 4133
rect 48112 4081 48118 4133
rect 48170 4121 48176 4133
rect 49072 4121 49078 4133
rect 48170 4093 49078 4121
rect 48170 4081 48176 4093
rect 49072 4081 49078 4093
rect 49130 4081 49136 4133
rect 49168 4081 49174 4133
rect 49226 4121 49232 4133
rect 50704 4121 50710 4133
rect 49226 4093 50710 4121
rect 49226 4081 49232 4093
rect 50704 4081 50710 4093
rect 50762 4081 50768 4133
rect 56272 4081 56278 4133
rect 56330 4121 56336 4133
rect 58000 4121 58006 4133
rect 56330 4093 58006 4121
rect 56330 4081 56336 4093
rect 58000 4081 58006 4093
rect 58058 4081 58064 4133
rect 1152 4022 58848 4044
rect 1152 3970 4294 4022
rect 4346 3970 4358 4022
rect 4410 3970 4422 4022
rect 4474 3970 4486 4022
rect 4538 3970 35014 4022
rect 35066 3970 35078 4022
rect 35130 3970 35142 4022
rect 35194 3970 35206 4022
rect 35258 3970 58848 4022
rect 1152 3948 58848 3970
rect 1936 3859 1942 3911
rect 1994 3899 2000 3911
rect 2992 3899 2998 3911
rect 1994 3871 2998 3899
rect 1994 3859 2000 3871
rect 2992 3859 2998 3871
rect 3050 3859 3056 3911
rect 8272 3859 8278 3911
rect 8330 3899 8336 3911
rect 10576 3899 10582 3911
rect 8330 3871 10582 3899
rect 8330 3859 8336 3871
rect 10576 3859 10582 3871
rect 10634 3859 10640 3911
rect 13168 3859 13174 3911
rect 13226 3899 13232 3911
rect 13939 3902 13997 3908
rect 13939 3899 13951 3902
rect 13226 3871 13951 3899
rect 13226 3859 13232 3871
rect 13939 3868 13951 3871
rect 13985 3868 13997 3902
rect 13939 3862 13997 3868
rect 14032 3859 14038 3911
rect 14090 3899 14096 3911
rect 15475 3902 15533 3908
rect 15475 3899 15487 3902
rect 14090 3871 15487 3899
rect 14090 3859 14096 3871
rect 15475 3868 15487 3871
rect 15521 3868 15533 3902
rect 15475 3862 15533 3868
rect 17779 3902 17837 3908
rect 17779 3868 17791 3902
rect 17825 3899 17837 3902
rect 18160 3899 18166 3911
rect 17825 3871 18166 3899
rect 17825 3868 17837 3871
rect 17779 3862 17837 3868
rect 18160 3859 18166 3871
rect 18218 3859 18224 3911
rect 18544 3899 18550 3911
rect 18505 3871 18550 3899
rect 18544 3859 18550 3871
rect 18602 3859 18608 3911
rect 21232 3859 21238 3911
rect 21290 3899 21296 3911
rect 22768 3899 22774 3911
rect 21290 3871 22774 3899
rect 21290 3859 21296 3871
rect 22768 3859 22774 3871
rect 22826 3859 22832 3911
rect 23920 3859 23926 3911
rect 23978 3899 23984 3911
rect 25072 3899 25078 3911
rect 23978 3871 25078 3899
rect 23978 3859 23984 3871
rect 25072 3859 25078 3871
rect 25130 3859 25136 3911
rect 27472 3859 27478 3911
rect 27530 3899 27536 3911
rect 28912 3899 28918 3911
rect 27530 3871 28918 3899
rect 27530 3859 27536 3871
rect 28912 3859 28918 3871
rect 28970 3859 28976 3911
rect 29008 3859 29014 3911
rect 29066 3899 29072 3911
rect 30352 3899 30358 3911
rect 29066 3871 30358 3899
rect 29066 3859 29072 3871
rect 30352 3859 30358 3871
rect 30410 3859 30416 3911
rect 38512 3859 38518 3911
rect 38570 3899 38576 3911
rect 40144 3899 40150 3911
rect 38570 3871 40150 3899
rect 38570 3859 38576 3871
rect 40144 3859 40150 3871
rect 40202 3859 40208 3911
rect 41296 3859 41302 3911
rect 41354 3899 41360 3911
rect 41488 3899 41494 3911
rect 41354 3871 41494 3899
rect 41354 3859 41360 3871
rect 41488 3859 41494 3871
rect 41546 3859 41552 3911
rect 43792 3899 43798 3911
rect 41698 3871 43798 3899
rect 496 3785 502 3837
rect 554 3825 560 3837
rect 1648 3825 1654 3837
rect 554 3797 1654 3825
rect 554 3785 560 3797
rect 1648 3785 1654 3797
rect 1706 3785 1712 3837
rect 2320 3785 2326 3837
rect 2378 3825 2384 3837
rect 3088 3825 3094 3837
rect 2378 3797 3094 3825
rect 2378 3785 2384 3797
rect 3088 3785 3094 3797
rect 3146 3785 3152 3837
rect 7888 3785 7894 3837
rect 7946 3825 7952 3837
rect 9232 3825 9238 3837
rect 7946 3797 9238 3825
rect 7946 3785 7952 3797
rect 9232 3785 9238 3797
rect 9290 3785 9296 3837
rect 12016 3785 12022 3837
rect 12074 3825 12080 3837
rect 13648 3825 13654 3837
rect 12074 3797 13654 3825
rect 12074 3785 12080 3797
rect 13648 3785 13654 3797
rect 13706 3785 13712 3837
rect 15280 3785 15286 3837
rect 15338 3785 15344 3837
rect 16528 3785 16534 3837
rect 16586 3825 16592 3837
rect 17296 3825 17302 3837
rect 16586 3797 17302 3825
rect 16586 3785 16592 3797
rect 17296 3785 17302 3797
rect 17354 3785 17360 3837
rect 19408 3785 19414 3837
rect 19466 3825 19472 3837
rect 20656 3825 20662 3837
rect 19466 3797 20662 3825
rect 19466 3785 19472 3797
rect 20656 3785 20662 3797
rect 20714 3785 20720 3837
rect 24208 3785 24214 3837
rect 24266 3825 24272 3837
rect 25840 3825 25846 3837
rect 24266 3797 25846 3825
rect 24266 3785 24272 3797
rect 25840 3785 25846 3797
rect 25898 3785 25904 3837
rect 26416 3785 26422 3837
rect 26474 3825 26480 3837
rect 28048 3825 28054 3837
rect 26474 3797 28054 3825
rect 26474 3785 26480 3797
rect 28048 3785 28054 3797
rect 28106 3785 28112 3837
rect 29392 3785 29398 3837
rect 29450 3825 29456 3837
rect 30448 3825 30454 3837
rect 29450 3797 30454 3825
rect 29450 3785 29456 3797
rect 30448 3785 30454 3797
rect 30506 3785 30512 3837
rect 33424 3785 33430 3837
rect 33482 3825 33488 3837
rect 34864 3825 34870 3837
rect 33482 3797 34870 3825
rect 33482 3785 33488 3797
rect 34864 3785 34870 3797
rect 34922 3785 34928 3837
rect 35632 3785 35638 3837
rect 35690 3825 35696 3837
rect 36400 3825 36406 3837
rect 35690 3797 36406 3825
rect 35690 3785 35696 3797
rect 36400 3785 36406 3797
rect 36458 3785 36464 3837
rect 37840 3785 37846 3837
rect 37898 3825 37904 3837
rect 39376 3825 39382 3837
rect 37898 3797 39382 3825
rect 37898 3785 37904 3797
rect 39376 3785 39382 3797
rect 39434 3785 39440 3837
rect 2992 3711 2998 3763
rect 3050 3751 3056 3763
rect 3280 3751 3286 3763
rect 3050 3723 3286 3751
rect 3050 3711 3056 3723
rect 3280 3711 3286 3723
rect 3338 3711 3344 3763
rect 3376 3711 3382 3763
rect 3434 3751 3440 3763
rect 15298 3751 15326 3785
rect 20083 3754 20141 3760
rect 20083 3751 20095 3754
rect 3434 3723 4670 3751
rect 15298 3723 20095 3751
rect 3434 3711 3440 3723
rect 112 3637 118 3689
rect 170 3677 176 3689
rect 1555 3680 1613 3686
rect 1555 3677 1567 3680
rect 170 3649 1567 3677
rect 170 3637 176 3649
rect 1555 3646 1567 3649
rect 1601 3646 1613 3680
rect 1555 3640 1613 3646
rect 1648 3637 1654 3689
rect 1706 3677 1712 3689
rect 2323 3680 2381 3686
rect 2323 3677 2335 3680
rect 1706 3649 2335 3677
rect 1706 3637 1712 3649
rect 2323 3646 2335 3649
rect 2369 3646 2381 3680
rect 2323 3640 2381 3646
rect 2704 3637 2710 3689
rect 2762 3677 2768 3689
rect 4642 3686 4670 3723
rect 20083 3720 20095 3723
rect 20129 3720 20141 3754
rect 20083 3714 20141 3720
rect 28720 3711 28726 3763
rect 28778 3751 28784 3763
rect 28778 3723 29630 3751
rect 28778 3711 28784 3723
rect 3091 3680 3149 3686
rect 3091 3677 3103 3680
rect 2762 3649 3103 3677
rect 2762 3637 2768 3649
rect 3091 3646 3103 3649
rect 3137 3646 3149 3680
rect 3091 3640 3149 3646
rect 3859 3680 3917 3686
rect 3859 3646 3871 3680
rect 3905 3646 3917 3680
rect 3859 3640 3917 3646
rect 4627 3680 4685 3686
rect 4627 3646 4639 3680
rect 4673 3646 4685 3680
rect 5584 3677 5590 3689
rect 5545 3649 5590 3677
rect 4627 3640 4685 3646
rect 3088 3489 3094 3541
rect 3146 3529 3152 3541
rect 3874 3529 3902 3640
rect 5584 3637 5590 3649
rect 5642 3637 5648 3689
rect 6352 3637 6358 3689
rect 6410 3677 6416 3689
rect 6931 3680 6989 3686
rect 6931 3677 6943 3680
rect 6410 3649 6943 3677
rect 6410 3637 6416 3649
rect 6931 3646 6943 3649
rect 6977 3646 6989 3680
rect 6931 3640 6989 3646
rect 7024 3637 7030 3689
rect 7082 3677 7088 3689
rect 7699 3680 7757 3686
rect 7699 3677 7711 3680
rect 7082 3649 7711 3677
rect 7082 3637 7088 3649
rect 7699 3646 7711 3649
rect 7745 3646 7757 3680
rect 7699 3640 7757 3646
rect 7792 3637 7798 3689
rect 7850 3677 7856 3689
rect 8467 3680 8525 3686
rect 8467 3677 8479 3680
rect 7850 3649 8479 3677
rect 7850 3637 7856 3649
rect 8467 3646 8479 3649
rect 8513 3646 8525 3680
rect 8467 3640 8525 3646
rect 8560 3637 8566 3689
rect 8618 3677 8624 3689
rect 9235 3680 9293 3686
rect 9235 3677 9247 3680
rect 8618 3649 9247 3677
rect 8618 3637 8624 3649
rect 9235 3646 9247 3649
rect 9281 3646 9293 3680
rect 9235 3640 9293 3646
rect 9328 3637 9334 3689
rect 9386 3677 9392 3689
rect 10003 3680 10061 3686
rect 10003 3677 10015 3680
rect 9386 3649 10015 3677
rect 9386 3637 9392 3649
rect 10003 3646 10015 3649
rect 10049 3646 10061 3680
rect 10003 3640 10061 3646
rect 10771 3680 10829 3686
rect 10771 3646 10783 3680
rect 10817 3646 10829 3680
rect 10771 3640 10829 3646
rect 12979 3680 13037 3686
rect 12979 3646 12991 3680
rect 13025 3677 13037 3680
rect 13168 3677 13174 3689
rect 13025 3649 13174 3677
rect 13025 3646 13037 3649
rect 12979 3640 13037 3646
rect 8080 3563 8086 3615
rect 8138 3603 8144 3615
rect 9712 3603 9718 3615
rect 8138 3575 9718 3603
rect 8138 3563 8144 3575
rect 9712 3563 9718 3575
rect 9770 3563 9776 3615
rect 3146 3501 3902 3529
rect 3146 3489 3152 3501
rect 5104 3489 5110 3541
rect 5162 3529 5168 3541
rect 5968 3529 5974 3541
rect 5162 3501 5974 3529
rect 5162 3489 5168 3501
rect 5968 3489 5974 3501
rect 6026 3489 6032 3541
rect 10000 3489 10006 3541
rect 10058 3529 10064 3541
rect 10786 3529 10814 3640
rect 13168 3637 13174 3649
rect 13226 3637 13232 3689
rect 13648 3677 13654 3689
rect 13609 3649 13654 3677
rect 13648 3637 13654 3649
rect 13706 3637 13712 3689
rect 14032 3637 14038 3689
rect 14090 3677 14096 3689
rect 14419 3680 14477 3686
rect 14419 3677 14431 3680
rect 14090 3649 14431 3677
rect 14090 3637 14096 3649
rect 14419 3646 14431 3649
rect 14465 3646 14477 3680
rect 14419 3640 14477 3646
rect 14800 3637 14806 3689
rect 14858 3677 14864 3689
rect 15187 3680 15245 3686
rect 15187 3677 15199 3680
rect 14858 3649 15199 3677
rect 14858 3637 14864 3649
rect 15187 3646 15199 3649
rect 15233 3646 15245 3680
rect 15187 3640 15245 3646
rect 15280 3637 15286 3689
rect 15338 3677 15344 3689
rect 15955 3680 16013 3686
rect 15955 3677 15967 3680
rect 15338 3649 15967 3677
rect 15338 3637 15344 3649
rect 15955 3646 15967 3649
rect 16001 3646 16013 3680
rect 15955 3640 16013 3646
rect 17392 3637 17398 3689
rect 17450 3677 17456 3689
rect 17491 3680 17549 3686
rect 17491 3677 17503 3680
rect 17450 3649 17503 3677
rect 17450 3637 17456 3649
rect 17491 3646 17503 3649
rect 17537 3646 17549 3680
rect 17491 3640 17549 3646
rect 18064 3637 18070 3689
rect 18122 3677 18128 3689
rect 18259 3680 18317 3686
rect 18259 3677 18271 3680
rect 18122 3649 18271 3677
rect 18122 3637 18128 3649
rect 18259 3646 18271 3649
rect 18305 3646 18317 3680
rect 18259 3640 18317 3646
rect 18448 3637 18454 3689
rect 18506 3677 18512 3689
rect 19027 3680 19085 3686
rect 19027 3677 19039 3680
rect 18506 3649 19039 3677
rect 18506 3637 18512 3649
rect 19027 3646 19039 3649
rect 19073 3646 19085 3680
rect 19027 3640 19085 3646
rect 19216 3637 19222 3689
rect 19274 3677 19280 3689
rect 19795 3680 19853 3686
rect 19795 3677 19807 3680
rect 19274 3649 19807 3677
rect 19274 3637 19280 3649
rect 19795 3646 19807 3649
rect 19841 3646 19853 3680
rect 19795 3640 19853 3646
rect 20656 3637 20662 3689
rect 20714 3677 20720 3689
rect 21331 3680 21389 3686
rect 21331 3677 21343 3680
rect 20714 3649 21343 3677
rect 20714 3637 20720 3649
rect 21331 3646 21343 3649
rect 21377 3646 21389 3680
rect 21331 3640 21389 3646
rect 22096 3637 22102 3689
rect 22154 3677 22160 3689
rect 22771 3680 22829 3686
rect 22771 3677 22783 3680
rect 22154 3649 22783 3677
rect 22154 3637 22160 3649
rect 22771 3646 22783 3649
rect 22817 3646 22829 3680
rect 22771 3640 22829 3646
rect 22864 3637 22870 3689
rect 22922 3677 22928 3689
rect 23539 3680 23597 3686
rect 23539 3677 23551 3680
rect 22922 3649 23551 3677
rect 22922 3637 22928 3649
rect 23539 3646 23551 3649
rect 23585 3646 23597 3680
rect 23539 3640 23597 3646
rect 23632 3637 23638 3689
rect 23690 3677 23696 3689
rect 24307 3680 24365 3686
rect 24307 3677 24319 3680
rect 23690 3649 24319 3677
rect 23690 3637 23696 3649
rect 24307 3646 24319 3649
rect 24353 3646 24365 3680
rect 24307 3640 24365 3646
rect 24400 3637 24406 3689
rect 24458 3677 24464 3689
rect 25075 3680 25133 3686
rect 25075 3677 25087 3680
rect 24458 3649 25087 3677
rect 24458 3637 24464 3649
rect 25075 3646 25087 3649
rect 25121 3646 25133 3680
rect 25075 3640 25133 3646
rect 25843 3680 25901 3686
rect 25843 3646 25855 3680
rect 25889 3646 25901 3680
rect 25843 3640 25901 3646
rect 26611 3680 26669 3686
rect 26611 3646 26623 3680
rect 26657 3646 26669 3680
rect 26611 3640 26669 3646
rect 19984 3563 19990 3615
rect 20042 3603 20048 3615
rect 20755 3606 20813 3612
rect 20755 3603 20767 3606
rect 20042 3575 20767 3603
rect 20042 3563 20048 3575
rect 20755 3572 20767 3575
rect 20801 3572 20813 3606
rect 20755 3566 20813 3572
rect 24688 3563 24694 3615
rect 24746 3603 24752 3615
rect 25858 3603 25886 3640
rect 24746 3575 25886 3603
rect 24746 3563 24752 3575
rect 10058 3501 10814 3529
rect 10058 3489 10064 3501
rect 15088 3489 15094 3541
rect 15146 3529 15152 3541
rect 15146 3501 20702 3529
rect 15146 3489 15152 3501
rect 592 3415 598 3467
rect 650 3455 656 3467
rect 1456 3455 1462 3467
rect 650 3427 1462 3455
rect 650 3415 656 3427
rect 1456 3415 1462 3427
rect 1514 3415 1520 3467
rect 3280 3415 3286 3467
rect 3338 3455 3344 3467
rect 3952 3455 3958 3467
rect 3338 3427 3958 3455
rect 3338 3415 3344 3427
rect 3952 3415 3958 3427
rect 4010 3415 4016 3467
rect 17296 3415 17302 3467
rect 17354 3455 17360 3467
rect 17488 3455 17494 3467
rect 17354 3427 17494 3455
rect 17354 3415 17360 3427
rect 17488 3415 17494 3427
rect 17546 3415 17552 3467
rect 20674 3464 20702 3501
rect 25840 3489 25846 3541
rect 25898 3529 25904 3541
rect 26626 3529 26654 3640
rect 27280 3637 27286 3689
rect 27338 3677 27344 3689
rect 29602 3686 29630 3723
rect 37744 3711 37750 3763
rect 37802 3751 37808 3763
rect 41698 3751 41726 3871
rect 43792 3859 43798 3871
rect 43850 3859 43856 3911
rect 43984 3859 43990 3911
rect 44042 3899 44048 3911
rect 44752 3899 44758 3911
rect 44042 3871 44758 3899
rect 44042 3859 44048 3871
rect 44752 3859 44758 3871
rect 44810 3859 44816 3911
rect 46288 3859 46294 3911
rect 46346 3899 46352 3911
rect 47632 3899 47638 3911
rect 46346 3871 47638 3899
rect 46346 3859 46352 3871
rect 47632 3859 47638 3871
rect 47690 3859 47696 3911
rect 48496 3859 48502 3911
rect 48554 3899 48560 3911
rect 49648 3899 49654 3911
rect 48554 3871 49654 3899
rect 48554 3859 48560 3871
rect 49648 3859 49654 3871
rect 49706 3859 49712 3911
rect 51376 3859 51382 3911
rect 51434 3899 51440 3911
rect 51856 3899 51862 3911
rect 51434 3871 51862 3899
rect 51434 3859 51440 3871
rect 51856 3859 51862 3871
rect 51914 3859 51920 3911
rect 55984 3859 55990 3911
rect 56042 3899 56048 3911
rect 57904 3899 57910 3911
rect 56042 3871 57910 3899
rect 56042 3859 56048 3871
rect 57904 3859 57910 3871
rect 57962 3859 57968 3911
rect 44080 3785 44086 3837
rect 44138 3825 44144 3837
rect 45424 3825 45430 3837
rect 44138 3797 45430 3825
rect 44138 3785 44144 3797
rect 45424 3785 45430 3797
rect 45482 3785 45488 3837
rect 46096 3785 46102 3837
rect 46154 3825 46160 3837
rect 47056 3825 47062 3837
rect 46154 3797 47062 3825
rect 46154 3785 46160 3797
rect 47056 3785 47062 3797
rect 47114 3785 47120 3837
rect 49072 3785 49078 3837
rect 49130 3825 49136 3837
rect 50032 3825 50038 3837
rect 49130 3797 50038 3825
rect 49130 3785 49136 3797
rect 50032 3785 50038 3797
rect 50090 3785 50096 3837
rect 37802 3723 41726 3751
rect 37802 3711 37808 3723
rect 45232 3711 45238 3763
rect 45290 3751 45296 3763
rect 45290 3723 46238 3751
rect 45290 3711 45296 3723
rect 28051 3680 28109 3686
rect 28051 3677 28063 3680
rect 27338 3649 28063 3677
rect 27338 3637 27344 3649
rect 28051 3646 28063 3649
rect 28097 3646 28109 3680
rect 28051 3640 28109 3646
rect 28819 3680 28877 3686
rect 28819 3646 28831 3680
rect 28865 3646 28877 3680
rect 28819 3640 28877 3646
rect 29587 3680 29645 3686
rect 29587 3646 29599 3680
rect 29633 3646 29645 3680
rect 29587 3640 29645 3646
rect 30355 3680 30413 3686
rect 30355 3646 30367 3680
rect 30401 3646 30413 3680
rect 30355 3640 30413 3646
rect 25898 3501 26654 3529
rect 25898 3489 25904 3501
rect 28048 3489 28054 3541
rect 28106 3529 28112 3541
rect 28834 3529 28862 3640
rect 29488 3563 29494 3615
rect 29546 3603 29552 3615
rect 30370 3603 30398 3640
rect 30448 3637 30454 3689
rect 30506 3677 30512 3689
rect 31123 3680 31181 3686
rect 31123 3677 31135 3680
rect 30506 3649 31135 3677
rect 30506 3637 30512 3649
rect 31123 3646 31135 3649
rect 31169 3646 31181 3680
rect 31123 3640 31181 3646
rect 31312 3637 31318 3689
rect 31370 3677 31376 3689
rect 31891 3680 31949 3686
rect 31891 3677 31903 3680
rect 31370 3649 31903 3677
rect 31370 3637 31376 3649
rect 31891 3646 31903 3649
rect 31937 3646 31949 3680
rect 31891 3640 31949 3646
rect 32464 3637 32470 3689
rect 32522 3677 32528 3689
rect 33331 3680 33389 3686
rect 33331 3677 33343 3680
rect 32522 3649 33343 3677
rect 32522 3637 32528 3649
rect 33331 3646 33343 3649
rect 33377 3646 33389 3680
rect 33331 3640 33389 3646
rect 33520 3637 33526 3689
rect 33578 3677 33584 3689
rect 34099 3680 34157 3686
rect 34099 3677 34111 3680
rect 33578 3649 34111 3677
rect 33578 3637 33584 3649
rect 34099 3646 34111 3649
rect 34145 3646 34157 3680
rect 34099 3640 34157 3646
rect 34288 3637 34294 3689
rect 34346 3677 34352 3689
rect 34867 3680 34925 3686
rect 34867 3677 34879 3680
rect 34346 3649 34879 3677
rect 34346 3637 34352 3649
rect 34867 3646 34879 3649
rect 34913 3646 34925 3680
rect 34867 3640 34925 3646
rect 34960 3637 34966 3689
rect 35018 3677 35024 3689
rect 35635 3680 35693 3686
rect 35635 3677 35647 3680
rect 35018 3649 35647 3677
rect 35018 3637 35024 3649
rect 35635 3646 35647 3649
rect 35681 3646 35693 3680
rect 35635 3640 35693 3646
rect 35728 3637 35734 3689
rect 35786 3677 35792 3689
rect 36403 3680 36461 3686
rect 36403 3677 36415 3680
rect 35786 3649 36415 3677
rect 35786 3637 35792 3649
rect 36403 3646 36415 3649
rect 36449 3646 36461 3680
rect 36403 3640 36461 3646
rect 36496 3637 36502 3689
rect 36554 3677 36560 3689
rect 37171 3680 37229 3686
rect 37171 3677 37183 3680
rect 36554 3649 37183 3677
rect 36554 3637 36560 3649
rect 37171 3646 37183 3649
rect 37217 3646 37229 3680
rect 37171 3640 37229 3646
rect 37936 3637 37942 3689
rect 37994 3677 38000 3689
rect 38611 3680 38669 3686
rect 38611 3677 38623 3680
rect 37994 3649 38623 3677
rect 37994 3637 38000 3649
rect 38611 3646 38623 3649
rect 38657 3646 38669 3680
rect 38611 3640 38669 3646
rect 38704 3637 38710 3689
rect 38762 3677 38768 3689
rect 39379 3680 39437 3686
rect 39379 3677 39391 3680
rect 38762 3649 39391 3677
rect 38762 3637 38768 3649
rect 39379 3646 39391 3649
rect 39425 3646 39437 3680
rect 39379 3640 39437 3646
rect 40147 3680 40205 3686
rect 40147 3646 40159 3680
rect 40193 3646 40205 3680
rect 40147 3640 40205 3646
rect 40915 3680 40973 3686
rect 40915 3646 40927 3680
rect 40961 3646 40973 3680
rect 40915 3640 40973 3646
rect 29546 3575 30398 3603
rect 29546 3563 29552 3575
rect 32848 3563 32854 3615
rect 32906 3603 32912 3615
rect 33712 3603 33718 3615
rect 32906 3575 33718 3603
rect 32906 3563 32912 3575
rect 33712 3563 33718 3575
rect 33770 3563 33776 3615
rect 28106 3501 28862 3529
rect 28106 3489 28112 3501
rect 28912 3489 28918 3541
rect 28970 3529 28976 3541
rect 29776 3529 29782 3541
rect 28970 3501 29782 3529
rect 28970 3489 28976 3501
rect 29776 3489 29782 3501
rect 29834 3489 29840 3541
rect 30448 3489 30454 3541
rect 30506 3529 30512 3541
rect 31888 3529 31894 3541
rect 30506 3501 31894 3529
rect 30506 3489 30512 3501
rect 31888 3489 31894 3501
rect 31946 3489 31952 3541
rect 35920 3489 35926 3541
rect 35978 3529 35984 3541
rect 36688 3529 36694 3541
rect 35978 3501 36694 3529
rect 35978 3489 35984 3501
rect 36688 3489 36694 3501
rect 36746 3489 36752 3541
rect 39376 3489 39382 3541
rect 39434 3529 39440 3541
rect 40162 3529 40190 3640
rect 39434 3501 40190 3529
rect 39434 3489 39440 3501
rect 20659 3458 20717 3464
rect 20659 3424 20671 3458
rect 20705 3424 20717 3458
rect 20659 3418 20717 3424
rect 36016 3415 36022 3467
rect 36074 3455 36080 3467
rect 36208 3455 36214 3467
rect 36074 3427 36214 3455
rect 36074 3415 36080 3427
rect 36208 3415 36214 3427
rect 36266 3415 36272 3467
rect 37072 3415 37078 3467
rect 37130 3455 37136 3467
rect 38608 3455 38614 3467
rect 37130 3427 38614 3455
rect 37130 3415 37136 3427
rect 38608 3415 38614 3427
rect 38666 3415 38672 3467
rect 40144 3415 40150 3467
rect 40202 3455 40208 3467
rect 40930 3455 40958 3640
rect 41008 3637 41014 3689
rect 41066 3677 41072 3689
rect 41683 3680 41741 3686
rect 41683 3677 41695 3680
rect 41066 3649 41695 3677
rect 41066 3637 41072 3649
rect 41683 3646 41695 3649
rect 41729 3646 41741 3680
rect 41683 3640 41741 3646
rect 42451 3680 42509 3686
rect 42451 3646 42463 3680
rect 42497 3646 42509 3680
rect 42451 3640 42509 3646
rect 41584 3563 41590 3615
rect 41642 3603 41648 3615
rect 42466 3603 42494 3640
rect 42736 3637 42742 3689
rect 42794 3677 42800 3689
rect 46210 3686 46238 3723
rect 43891 3680 43949 3686
rect 43891 3677 43903 3680
rect 42794 3649 43903 3677
rect 42794 3637 42800 3649
rect 43891 3646 43903 3649
rect 43937 3646 43949 3680
rect 44659 3680 44717 3686
rect 44659 3677 44671 3680
rect 43891 3640 43949 3646
rect 44002 3649 44671 3677
rect 41642 3575 42494 3603
rect 41642 3563 41648 3575
rect 43792 3563 43798 3615
rect 43850 3603 43856 3615
rect 44002 3603 44030 3649
rect 44659 3646 44671 3649
rect 44705 3646 44717 3680
rect 44659 3640 44717 3646
rect 45427 3680 45485 3686
rect 45427 3646 45439 3680
rect 45473 3646 45485 3680
rect 45427 3640 45485 3646
rect 46195 3680 46253 3686
rect 46195 3646 46207 3680
rect 46241 3646 46253 3680
rect 46195 3640 46253 3646
rect 46963 3680 47021 3686
rect 46963 3646 46975 3680
rect 47009 3646 47021 3680
rect 46963 3640 47021 3646
rect 43850 3575 44030 3603
rect 43850 3563 43856 3575
rect 44560 3563 44566 3615
rect 44618 3603 44624 3615
rect 45442 3603 45470 3640
rect 44618 3575 45470 3603
rect 44618 3563 44624 3575
rect 46000 3563 46006 3615
rect 46058 3603 46064 3615
rect 46978 3603 47006 3640
rect 47152 3637 47158 3689
rect 47210 3677 47216 3689
rect 47731 3680 47789 3686
rect 47731 3677 47743 3680
rect 47210 3649 47743 3677
rect 47210 3637 47216 3649
rect 47731 3646 47743 3649
rect 47777 3646 47789 3680
rect 47731 3640 47789 3646
rect 48208 3637 48214 3689
rect 48266 3677 48272 3689
rect 49171 3680 49229 3686
rect 49171 3677 49183 3680
rect 48266 3649 49183 3677
rect 48266 3637 48272 3649
rect 49171 3646 49183 3649
rect 49217 3646 49229 3680
rect 49171 3640 49229 3646
rect 50515 3680 50573 3686
rect 50515 3646 50527 3680
rect 50561 3677 50573 3680
rect 50704 3677 50710 3689
rect 50561 3649 50710 3677
rect 50561 3646 50573 3649
rect 50515 3640 50573 3646
rect 50704 3637 50710 3649
rect 50762 3637 50768 3689
rect 50800 3637 50806 3689
rect 50858 3677 50864 3689
rect 51187 3680 51245 3686
rect 51187 3677 51199 3680
rect 50858 3649 51199 3677
rect 50858 3637 50864 3649
rect 51187 3646 51199 3649
rect 51233 3646 51245 3680
rect 51187 3640 51245 3646
rect 51280 3637 51286 3689
rect 51338 3677 51344 3689
rect 51955 3680 52013 3686
rect 51955 3677 51967 3680
rect 51338 3649 51967 3677
rect 51338 3637 51344 3649
rect 51955 3646 51967 3649
rect 52001 3646 52013 3680
rect 51955 3640 52013 3646
rect 52048 3637 52054 3689
rect 52106 3677 52112 3689
rect 52723 3680 52781 3686
rect 52723 3677 52735 3680
rect 52106 3649 52735 3677
rect 52106 3637 52112 3649
rect 52723 3646 52735 3649
rect 52769 3646 52781 3680
rect 52723 3640 52781 3646
rect 53392 3637 53398 3689
rect 53450 3677 53456 3689
rect 54451 3680 54509 3686
rect 54451 3677 54463 3680
rect 53450 3649 54463 3677
rect 53450 3637 53456 3649
rect 54451 3646 54463 3649
rect 54497 3646 54509 3680
rect 54451 3640 54509 3646
rect 55219 3680 55277 3686
rect 55219 3646 55231 3680
rect 55265 3646 55277 3680
rect 55219 3640 55277 3646
rect 46058 3575 47006 3603
rect 46058 3563 46064 3575
rect 47632 3563 47638 3615
rect 47690 3603 47696 3615
rect 48400 3603 48406 3615
rect 47690 3575 48406 3603
rect 47690 3563 47696 3575
rect 48400 3563 48406 3575
rect 48458 3563 48464 3615
rect 54352 3563 54358 3615
rect 54410 3603 54416 3615
rect 55234 3603 55262 3640
rect 55312 3637 55318 3689
rect 55370 3677 55376 3689
rect 55987 3680 56045 3686
rect 55987 3677 55999 3680
rect 55370 3649 55999 3677
rect 55370 3637 55376 3649
rect 55987 3646 55999 3649
rect 56033 3646 56045 3680
rect 55987 3640 56045 3646
rect 56755 3680 56813 3686
rect 56755 3646 56767 3680
rect 56801 3646 56813 3680
rect 56755 3640 56813 3646
rect 57523 3680 57581 3686
rect 57523 3646 57535 3680
rect 57569 3646 57581 3680
rect 57523 3640 57581 3646
rect 54410 3575 55262 3603
rect 54410 3563 54416 3575
rect 55888 3563 55894 3615
rect 55946 3603 55952 3615
rect 56770 3603 56798 3640
rect 55946 3575 56798 3603
rect 55946 3563 55952 3575
rect 44752 3489 44758 3541
rect 44810 3529 44816 3541
rect 46192 3529 46198 3541
rect 44810 3501 46198 3529
rect 44810 3489 44816 3501
rect 46192 3489 46198 3501
rect 46250 3489 46256 3541
rect 51280 3489 51286 3541
rect 51338 3529 51344 3541
rect 51568 3529 51574 3541
rect 51338 3501 51574 3529
rect 51338 3489 51344 3501
rect 51568 3489 51574 3501
rect 51626 3489 51632 3541
rect 52048 3489 52054 3541
rect 52106 3529 52112 3541
rect 52240 3529 52246 3541
rect 52106 3501 52246 3529
rect 52106 3489 52112 3501
rect 52240 3489 52246 3501
rect 52298 3489 52304 3541
rect 56272 3489 56278 3541
rect 56330 3529 56336 3541
rect 57538 3529 57566 3640
rect 56330 3501 57566 3529
rect 56330 3489 56336 3501
rect 40202 3427 40958 3455
rect 40202 3415 40208 3427
rect 42544 3415 42550 3467
rect 42602 3455 42608 3467
rect 43504 3455 43510 3467
rect 42602 3427 43510 3455
rect 42602 3415 42608 3427
rect 43504 3415 43510 3427
rect 43562 3415 43568 3467
rect 1152 3356 58848 3378
rect 1152 3304 19654 3356
rect 19706 3304 19718 3356
rect 19770 3304 19782 3356
rect 19834 3304 19846 3356
rect 19898 3304 50374 3356
rect 50426 3304 50438 3356
rect 50490 3304 50502 3356
rect 50554 3304 50566 3356
rect 50618 3304 58848 3356
rect 1152 3282 58848 3304
rect 1456 3193 1462 3245
rect 1514 3233 1520 3245
rect 2224 3233 2230 3245
rect 1514 3205 2230 3233
rect 1514 3193 1520 3205
rect 2224 3193 2230 3205
rect 2282 3193 2288 3245
rect 3952 3193 3958 3245
rect 4010 3233 4016 3245
rect 5200 3233 5206 3245
rect 4010 3205 5206 3233
rect 4010 3193 4016 3205
rect 5200 3193 5206 3205
rect 5258 3193 5264 3245
rect 12304 3193 12310 3245
rect 12362 3233 12368 3245
rect 13072 3233 13078 3245
rect 12362 3205 13078 3233
rect 12362 3193 12368 3205
rect 13072 3193 13078 3205
rect 13130 3193 13136 3245
rect 13264 3233 13270 3245
rect 13225 3205 13270 3233
rect 13264 3193 13270 3205
rect 13322 3193 13328 3245
rect 13360 3193 13366 3245
rect 13418 3233 13424 3245
rect 14035 3236 14093 3242
rect 14035 3233 14047 3236
rect 13418 3205 14047 3233
rect 13418 3193 13424 3205
rect 14035 3202 14047 3205
rect 14081 3202 14093 3236
rect 14035 3196 14093 3202
rect 14128 3193 14134 3245
rect 14186 3233 14192 3245
rect 15379 3236 15437 3242
rect 15379 3233 15391 3236
rect 14186 3205 15391 3233
rect 14186 3193 14192 3205
rect 15379 3202 15391 3205
rect 15425 3202 15437 3236
rect 15379 3196 15437 3202
rect 17584 3193 17590 3245
rect 17642 3233 17648 3245
rect 18067 3236 18125 3242
rect 18067 3233 18079 3236
rect 17642 3205 18079 3233
rect 17642 3193 17648 3205
rect 18067 3202 18079 3205
rect 18113 3202 18125 3236
rect 18067 3196 18125 3202
rect 20755 3236 20813 3242
rect 20755 3202 20767 3236
rect 20801 3233 20813 3236
rect 20944 3233 20950 3245
rect 20801 3205 20950 3233
rect 20801 3202 20813 3205
rect 20755 3196 20813 3202
rect 20944 3193 20950 3205
rect 21002 3193 21008 3245
rect 22768 3193 22774 3245
rect 22826 3233 22832 3245
rect 23152 3233 23158 3245
rect 22826 3205 23158 3233
rect 22826 3193 22832 3205
rect 23152 3193 23158 3205
rect 23210 3193 23216 3245
rect 28240 3193 28246 3245
rect 28298 3233 28304 3245
rect 29296 3233 29302 3245
rect 28298 3205 29302 3233
rect 28298 3193 28304 3205
rect 29296 3193 29302 3205
rect 29354 3193 29360 3245
rect 31888 3193 31894 3245
rect 31946 3233 31952 3245
rect 33328 3233 33334 3245
rect 31946 3205 33334 3233
rect 31946 3193 31952 3205
rect 33328 3193 33334 3205
rect 33386 3193 33392 3245
rect 33808 3193 33814 3245
rect 33866 3233 33872 3245
rect 35056 3233 35062 3245
rect 33866 3205 35062 3233
rect 33866 3193 33872 3205
rect 35056 3193 35062 3205
rect 35114 3193 35120 3245
rect 36688 3193 36694 3245
rect 36746 3233 36752 3245
rect 37552 3233 37558 3245
rect 36746 3205 37558 3233
rect 36746 3193 36752 3205
rect 37552 3193 37558 3205
rect 37610 3193 37616 3245
rect 41488 3193 41494 3245
rect 41546 3233 41552 3245
rect 41776 3233 41782 3245
rect 41546 3205 41782 3233
rect 41546 3193 41552 3205
rect 41776 3193 41782 3205
rect 41834 3193 41840 3245
rect 43312 3233 43318 3245
rect 43273 3205 43318 3233
rect 43312 3193 43318 3205
rect 43370 3193 43376 3245
rect 44176 3233 44182 3245
rect 43426 3205 44182 3233
rect 208 3119 214 3171
rect 266 3159 272 3171
rect 1744 3159 1750 3171
rect 266 3131 1750 3159
rect 266 3119 272 3131
rect 1744 3119 1750 3131
rect 1802 3119 1808 3171
rect 12208 3119 12214 3171
rect 12266 3159 12272 3171
rect 12976 3159 12982 3171
rect 12266 3131 12982 3159
rect 12266 3119 12272 3131
rect 12976 3119 12982 3131
rect 13034 3119 13040 3171
rect 13744 3159 13750 3171
rect 13090 3131 13750 3159
rect 13090 3097 13118 3131
rect 13744 3119 13750 3131
rect 13802 3119 13808 3171
rect 17776 3119 17782 3171
rect 17834 3159 17840 3171
rect 18835 3162 18893 3168
rect 18835 3159 18847 3162
rect 17834 3131 18847 3159
rect 17834 3119 17840 3131
rect 18835 3128 18847 3131
rect 18881 3128 18893 3162
rect 18835 3122 18893 3128
rect 19792 3119 19798 3171
rect 19850 3159 19856 3171
rect 20176 3159 20182 3171
rect 19850 3131 20182 3159
rect 19850 3119 19856 3131
rect 20176 3119 20182 3131
rect 20234 3119 20240 3171
rect 22384 3119 22390 3171
rect 22442 3159 22448 3171
rect 23536 3159 23542 3171
rect 22442 3131 23542 3159
rect 22442 3119 22448 3131
rect 23536 3119 23542 3131
rect 23594 3119 23600 3171
rect 25360 3119 25366 3171
rect 25418 3159 25424 3171
rect 26224 3159 26230 3171
rect 25418 3131 26230 3159
rect 25418 3119 25424 3131
rect 26224 3119 26230 3131
rect 26282 3119 26288 3171
rect 32656 3119 32662 3171
rect 32714 3159 32720 3171
rect 34096 3159 34102 3171
rect 32714 3131 34102 3159
rect 32714 3119 32720 3131
rect 34096 3119 34102 3131
rect 34154 3119 34160 3171
rect 34672 3119 34678 3171
rect 34730 3159 34736 3171
rect 35344 3159 35350 3171
rect 34730 3131 35350 3159
rect 34730 3119 34736 3131
rect 35344 3119 35350 3131
rect 35402 3119 35408 3171
rect 36208 3119 36214 3171
rect 36266 3159 36272 3171
rect 36266 3131 37406 3159
rect 36266 3119 36272 3131
rect 13072 3045 13078 3097
rect 13130 3045 13136 3097
rect 17488 3045 17494 3097
rect 17546 3085 17552 3097
rect 18352 3085 18358 3097
rect 17546 3057 18358 3085
rect 17546 3045 17552 3057
rect 18352 3045 18358 3057
rect 18410 3045 18416 3097
rect 19600 3045 19606 3097
rect 19658 3085 19664 3097
rect 19658 3057 20606 3085
rect 19658 3045 19664 3057
rect 16 2971 22 3023
rect 74 3011 80 3023
rect 1555 3014 1613 3020
rect 1555 3011 1567 3014
rect 74 2983 1567 3011
rect 74 2971 80 2983
rect 1555 2980 1567 2983
rect 1601 2980 1613 3014
rect 2323 3014 2381 3020
rect 2323 3011 2335 3014
rect 1555 2974 1613 2980
rect 1666 2983 2335 3011
rect 688 2897 694 2949
rect 746 2937 752 2949
rect 1666 2937 1694 2983
rect 2323 2980 2335 2983
rect 2369 2980 2381 3014
rect 3091 3014 3149 3020
rect 3091 3011 3103 3014
rect 2323 2974 2381 2980
rect 2866 2983 3103 3011
rect 746 2909 1694 2937
rect 746 2897 752 2909
rect 2128 2897 2134 2949
rect 2186 2937 2192 2949
rect 2866 2937 2894 2983
rect 3091 2980 3103 2983
rect 3137 2980 3149 3014
rect 4912 3011 4918 3023
rect 4873 2983 4918 3011
rect 3091 2974 3149 2980
rect 4912 2971 4918 2983
rect 4970 2971 4976 3023
rect 5200 2971 5206 3023
rect 5258 3011 5264 3023
rect 5683 3014 5741 3020
rect 5683 3011 5695 3014
rect 5258 2983 5695 3011
rect 5258 2971 5264 2983
rect 5683 2980 5695 2983
rect 5729 2980 5741 3014
rect 5683 2974 5741 2980
rect 5968 2971 5974 3023
rect 6026 3011 6032 3023
rect 7027 3014 7085 3020
rect 7027 3011 7039 3014
rect 6026 2983 7039 3011
rect 6026 2971 6032 2983
rect 7027 2980 7039 2983
rect 7073 2980 7085 3014
rect 7027 2974 7085 2980
rect 7795 3014 7853 3020
rect 7795 2980 7807 3014
rect 7841 2980 7853 3014
rect 7795 2974 7853 2980
rect 2186 2909 2894 2937
rect 2186 2897 2192 2909
rect 6736 2897 6742 2949
rect 6794 2937 6800 2949
rect 7810 2937 7838 2974
rect 8176 2971 8182 3023
rect 8234 3011 8240 3023
rect 9715 3014 9773 3020
rect 9715 3011 9727 3014
rect 8234 2983 9727 3011
rect 8234 2971 8240 2983
rect 9715 2980 9727 2983
rect 9761 2980 9773 3014
rect 9715 2974 9773 2980
rect 10483 3014 10541 3020
rect 10483 2980 10495 3014
rect 10529 2980 10541 3014
rect 10483 2974 10541 2980
rect 6794 2909 7838 2937
rect 6794 2897 6800 2909
rect 8944 2897 8950 2949
rect 9002 2937 9008 2949
rect 10498 2937 10526 2974
rect 11728 2971 11734 3023
rect 11786 3011 11792 3023
rect 12400 3011 12406 3023
rect 11786 2983 12406 3011
rect 11786 2971 11792 2983
rect 12400 2971 12406 2983
rect 12458 2971 12464 3023
rect 12976 3011 12982 3023
rect 12937 2983 12982 3011
rect 12976 2971 12982 2983
rect 13034 2971 13040 3023
rect 13360 2971 13366 3023
rect 13418 3011 13424 3023
rect 13747 3014 13805 3020
rect 13747 3011 13759 3014
rect 13418 2983 13759 3011
rect 13418 2971 13424 2983
rect 13747 2980 13759 2983
rect 13793 2980 13805 3014
rect 13747 2974 13805 2980
rect 14512 2971 14518 3023
rect 14570 3011 14576 3023
rect 15091 3014 15149 3020
rect 15091 3011 15103 3014
rect 14570 2983 15103 3011
rect 14570 2971 14576 2983
rect 15091 2980 15103 2983
rect 15137 2980 15149 3014
rect 16624 3011 16630 3023
rect 16585 2983 16630 3011
rect 15091 2974 15149 2980
rect 16624 2971 16630 2983
rect 16682 2971 16688 3023
rect 17008 2971 17014 3023
rect 17066 3011 17072 3023
rect 17779 3014 17837 3020
rect 17779 3011 17791 3014
rect 17066 2983 17791 3011
rect 17066 2971 17072 2983
rect 17779 2980 17791 2983
rect 17825 2980 17837 3014
rect 18547 3014 18605 3020
rect 18547 3011 18559 3014
rect 17779 2974 17837 2980
rect 17890 2983 18559 3011
rect 9002 2909 10526 2937
rect 9002 2897 9008 2909
rect 15376 2897 15382 2949
rect 15434 2937 15440 2949
rect 16432 2937 16438 2949
rect 15434 2909 16438 2937
rect 15434 2897 15440 2909
rect 16432 2897 16438 2909
rect 16490 2897 16496 2949
rect 17680 2897 17686 2949
rect 17738 2937 17744 2949
rect 17890 2937 17918 2983
rect 18547 2980 18559 2983
rect 18593 2980 18605 3014
rect 18547 2974 18605 2980
rect 18832 2971 18838 3023
rect 18890 3011 18896 3023
rect 20467 3014 20525 3020
rect 20467 3011 20479 3014
rect 18890 2983 20479 3011
rect 18890 2971 18896 2983
rect 20467 2980 20479 2983
rect 20513 2980 20525 3014
rect 20578 3011 20606 3057
rect 20944 3045 20950 3097
rect 21002 3085 21008 3097
rect 21712 3085 21718 3097
rect 21002 3057 21718 3085
rect 21002 3045 21008 3057
rect 21712 3045 21718 3057
rect 21770 3045 21776 3097
rect 22480 3045 22486 3097
rect 22538 3085 22544 3097
rect 22538 3057 23966 3085
rect 22538 3045 22544 3057
rect 21235 3014 21293 3020
rect 21235 3011 21247 3014
rect 20578 2983 21247 3011
rect 20467 2974 20525 2980
rect 21235 2980 21247 2983
rect 21281 2980 21293 3014
rect 21235 2974 21293 2980
rect 21424 2971 21430 3023
rect 21482 3011 21488 3023
rect 23938 3020 23966 3057
rect 25072 3045 25078 3097
rect 25130 3085 25136 3097
rect 25130 3057 26654 3085
rect 25130 3045 25136 3057
rect 23155 3014 23213 3020
rect 23155 3011 23167 3014
rect 21482 2983 23167 3011
rect 21482 2971 21488 2983
rect 23155 2980 23167 2983
rect 23201 2980 23213 3014
rect 23155 2974 23213 2980
rect 23923 3014 23981 3020
rect 23923 2980 23935 3014
rect 23969 2980 23981 3014
rect 23923 2974 23981 2980
rect 24016 2971 24022 3023
rect 24074 3011 24080 3023
rect 26626 3020 26654 3057
rect 27664 3045 27670 3097
rect 27722 3085 27728 3097
rect 27722 3057 29342 3085
rect 27722 3045 27728 3057
rect 25843 3014 25901 3020
rect 25843 3011 25855 3014
rect 24074 2983 25855 3011
rect 24074 2971 24080 2983
rect 25843 2980 25855 2983
rect 25889 2980 25901 3014
rect 25843 2974 25901 2980
rect 26611 3014 26669 3020
rect 26611 2980 26623 3014
rect 26657 2980 26669 3014
rect 26611 2974 26669 2980
rect 26896 2971 26902 3023
rect 26954 3011 26960 3023
rect 29314 3020 29342 3057
rect 30544 3045 30550 3097
rect 30602 3085 30608 3097
rect 30602 3057 32030 3085
rect 30602 3045 30608 3057
rect 28531 3014 28589 3020
rect 28531 3011 28543 3014
rect 26954 2983 28543 3011
rect 26954 2971 26960 2983
rect 28531 2980 28543 2983
rect 28577 2980 28589 3014
rect 28531 2974 28589 2980
rect 29299 3014 29357 3020
rect 29299 2980 29311 3014
rect 29345 2980 29357 3014
rect 29299 2974 29357 2980
rect 29872 2971 29878 3023
rect 29930 3011 29936 3023
rect 32002 3020 32030 3057
rect 32080 3045 32086 3097
rect 32138 3085 32144 3097
rect 32138 3057 33278 3085
rect 32138 3045 32144 3057
rect 31219 3014 31277 3020
rect 31219 3011 31231 3014
rect 29930 2983 31231 3011
rect 29930 2971 29936 2983
rect 31219 2980 31231 2983
rect 31265 2980 31277 3014
rect 31219 2974 31277 2980
rect 31987 3014 32045 3020
rect 31987 2980 31999 3014
rect 32033 2980 32045 3014
rect 31987 2974 32045 2980
rect 32272 2971 32278 3023
rect 32330 3011 32336 3023
rect 33136 3011 33142 3023
rect 32330 2983 33142 3011
rect 32330 2971 32336 2983
rect 33136 2971 33142 2983
rect 33194 2971 33200 3023
rect 33250 3011 33278 3057
rect 33328 3045 33334 3097
rect 33386 3085 33392 3097
rect 33386 3057 34718 3085
rect 33386 3045 33392 3057
rect 34690 3020 34718 3057
rect 35440 3045 35446 3097
rect 35498 3085 35504 3097
rect 35498 3057 36638 3085
rect 35498 3045 35504 3057
rect 33907 3014 33965 3020
rect 33907 3011 33919 3014
rect 33250 2983 33919 3011
rect 33907 2980 33919 2983
rect 33953 2980 33965 3014
rect 33907 2974 33965 2980
rect 34675 3014 34733 3020
rect 34675 2980 34687 3014
rect 34721 2980 34733 3014
rect 34675 2974 34733 2980
rect 35344 2971 35350 3023
rect 35402 3011 35408 3023
rect 36112 3011 36118 3023
rect 35402 2983 36118 3011
rect 35402 2971 35408 2983
rect 36112 2971 36118 2983
rect 36170 2971 36176 3023
rect 36610 3020 36638 3057
rect 37378 3020 37406 3131
rect 39664 3119 39670 3171
rect 39722 3159 39728 3171
rect 40912 3159 40918 3171
rect 39722 3131 40918 3159
rect 39722 3119 39728 3131
rect 40912 3119 40918 3131
rect 40970 3119 40976 3171
rect 41104 3119 41110 3171
rect 41162 3159 41168 3171
rect 42064 3159 42070 3171
rect 41162 3131 42070 3159
rect 41162 3119 41168 3131
rect 42064 3119 42070 3131
rect 42122 3119 42128 3171
rect 38320 3045 38326 3097
rect 38378 3085 38384 3097
rect 38378 3057 40094 3085
rect 38378 3045 38384 3057
rect 36595 3014 36653 3020
rect 36595 2980 36607 3014
rect 36641 2980 36653 3014
rect 36595 2974 36653 2980
rect 37363 3014 37421 3020
rect 37363 2980 37375 3014
rect 37409 2980 37421 3014
rect 37363 2974 37421 2980
rect 37552 2971 37558 3023
rect 37610 3011 37616 3023
rect 40066 3020 40094 3057
rect 41200 3045 41206 3097
rect 41258 3085 41264 3097
rect 43330 3085 43358 3193
rect 41258 3057 42782 3085
rect 41258 3045 41264 3057
rect 39283 3014 39341 3020
rect 39283 3011 39295 3014
rect 37610 2983 39295 3011
rect 37610 2971 37616 2983
rect 39283 2980 39295 2983
rect 39329 2980 39341 3014
rect 39283 2974 39341 2980
rect 40051 3014 40109 3020
rect 40051 2980 40063 3014
rect 40097 2980 40109 3014
rect 40051 2974 40109 2980
rect 40528 2971 40534 3023
rect 40586 3011 40592 3023
rect 42754 3020 42782 3057
rect 43234 3057 43358 3085
rect 41971 3014 42029 3020
rect 41971 3011 41983 3014
rect 40586 2983 41983 3011
rect 40586 2971 40592 2983
rect 41971 2980 41983 2983
rect 42017 2980 42029 3014
rect 41971 2974 42029 2980
rect 42739 3014 42797 3020
rect 42739 2980 42751 3014
rect 42785 2980 42797 3014
rect 42739 2974 42797 2980
rect 17738 2909 17918 2937
rect 17738 2897 17744 2909
rect 17968 2897 17974 2949
rect 18026 2937 18032 2949
rect 18256 2937 18262 2949
rect 18026 2909 18262 2937
rect 18026 2897 18032 2909
rect 18256 2897 18262 2909
rect 18314 2897 18320 2949
rect 18352 2897 18358 2949
rect 18410 2937 18416 2949
rect 19024 2937 19030 2949
rect 18410 2909 19030 2937
rect 18410 2897 18416 2909
rect 19024 2897 19030 2909
rect 19082 2897 19088 2949
rect 19219 2940 19277 2946
rect 19219 2906 19231 2940
rect 19265 2937 19277 2940
rect 19507 2940 19565 2946
rect 19507 2937 19519 2940
rect 19265 2909 19519 2937
rect 19265 2906 19277 2909
rect 19219 2900 19277 2906
rect 19507 2906 19519 2909
rect 19553 2937 19565 2940
rect 37744 2937 37750 2949
rect 19553 2909 37750 2937
rect 19553 2906 19565 2909
rect 19507 2900 19565 2906
rect 37744 2897 37750 2909
rect 37802 2897 37808 2949
rect 38128 2897 38134 2949
rect 38186 2937 38192 2949
rect 39088 2937 39094 2949
rect 38186 2909 39094 2937
rect 38186 2897 38192 2909
rect 39088 2897 39094 2909
rect 39146 2897 39152 2949
rect 40723 2940 40781 2946
rect 40723 2906 40735 2940
rect 40769 2937 40781 2940
rect 41011 2940 41069 2946
rect 41011 2937 41023 2940
rect 40769 2909 41023 2937
rect 40769 2906 40781 2909
rect 40723 2900 40781 2906
rect 41011 2906 41023 2909
rect 41057 2937 41069 2940
rect 41776 2937 41782 2949
rect 41057 2909 41782 2937
rect 41057 2906 41069 2909
rect 41011 2900 41069 2906
rect 41776 2897 41782 2909
rect 41834 2897 41840 2949
rect 43234 2937 43262 3057
rect 43312 2971 43318 3023
rect 43370 3011 43376 3023
rect 43426 3011 43454 3205
rect 44176 3193 44182 3205
rect 44234 3193 44240 3245
rect 55312 3193 55318 3245
rect 55370 3233 55376 3245
rect 55504 3233 55510 3245
rect 55370 3205 55510 3233
rect 55370 3193 55376 3205
rect 55504 3193 55510 3205
rect 55562 3193 55568 3245
rect 58192 3233 58198 3245
rect 55618 3205 58198 3233
rect 44368 3119 44374 3171
rect 44426 3159 44432 3171
rect 55618 3159 55646 3205
rect 58192 3193 58198 3205
rect 58250 3193 58256 3245
rect 44426 3131 55646 3159
rect 44426 3119 44432 3131
rect 57712 3119 57718 3171
rect 57770 3159 57776 3171
rect 59440 3159 59446 3171
rect 57770 3131 59446 3159
rect 57770 3119 57776 3131
rect 59440 3119 59446 3131
rect 59498 3119 59504 3171
rect 44176 3045 44182 3097
rect 44234 3085 44240 3097
rect 51763 3088 51821 3094
rect 44234 3057 45470 3085
rect 44234 3045 44240 3057
rect 45442 3020 45470 3057
rect 51763 3054 51775 3088
rect 51809 3085 51821 3088
rect 52432 3085 52438 3097
rect 51809 3057 52438 3085
rect 51809 3054 51821 3057
rect 51763 3048 51821 3054
rect 52432 3045 52438 3057
rect 52490 3045 52496 3097
rect 43370 2983 43454 3011
rect 44659 3014 44717 3020
rect 43370 2971 43376 2983
rect 44659 2980 44671 3014
rect 44705 2980 44717 3014
rect 44659 2974 44717 2980
rect 45427 3014 45485 3020
rect 45427 2980 45439 3014
rect 45473 2980 45485 3014
rect 45427 2974 45485 2980
rect 43507 2940 43565 2946
rect 43507 2937 43519 2940
rect 43234 2909 43519 2937
rect 43507 2906 43519 2909
rect 43553 2906 43565 2940
rect 43507 2900 43565 2906
rect 44368 2897 44374 2949
rect 44426 2937 44432 2949
rect 44674 2937 44702 2974
rect 45616 2971 45622 3023
rect 45674 3011 45680 3023
rect 47347 3014 47405 3020
rect 47347 3011 47359 3014
rect 45674 2983 47359 3011
rect 45674 2971 45680 2983
rect 47347 2980 47359 2983
rect 47393 2980 47405 3014
rect 47347 2974 47405 2980
rect 48115 3014 48173 3020
rect 48115 2980 48127 3014
rect 48161 2980 48173 3014
rect 48115 2974 48173 2980
rect 44426 2909 44702 2937
rect 44426 2897 44432 2909
rect 46384 2897 46390 2949
rect 46442 2937 46448 2949
rect 48130 2937 48158 2974
rect 49648 2971 49654 3023
rect 49706 3011 49712 3023
rect 50035 3014 50093 3020
rect 50035 3011 50047 3014
rect 49706 2983 50047 3011
rect 49706 2971 49712 2983
rect 50035 2980 50047 2983
rect 50081 2980 50093 3014
rect 50035 2974 50093 2980
rect 50803 3014 50861 3020
rect 50803 2980 50815 3014
rect 50849 2980 50861 3014
rect 50803 2974 50861 2980
rect 50818 2937 50846 2974
rect 51472 2971 51478 3023
rect 51530 3011 51536 3023
rect 52723 3014 52781 3020
rect 52723 3011 52735 3014
rect 51530 2983 52735 3011
rect 51530 2971 51536 2983
rect 52723 2980 52735 2983
rect 52769 2980 52781 3014
rect 53491 3014 53549 3020
rect 53491 3011 53503 3014
rect 52723 2974 52781 2980
rect 52834 2983 53503 3011
rect 46442 2909 48158 2937
rect 50050 2909 50846 2937
rect 46442 2897 46448 2909
rect 50050 2875 50078 2909
rect 52240 2897 52246 2949
rect 52298 2937 52304 2949
rect 52834 2937 52862 2983
rect 53491 2980 53503 2983
rect 53537 2980 53549 3014
rect 53491 2974 53549 2980
rect 53776 2971 53782 3023
rect 53834 3011 53840 3023
rect 55411 3014 55469 3020
rect 55411 3011 55423 3014
rect 53834 2983 55423 3011
rect 53834 2971 53840 2983
rect 55411 2980 55423 2983
rect 55457 2980 55469 3014
rect 55411 2974 55469 2980
rect 56179 3014 56237 3020
rect 56179 2980 56191 3014
rect 56225 2980 56237 3014
rect 56179 2974 56237 2980
rect 52298 2909 52862 2937
rect 52298 2897 52304 2909
rect 52912 2897 52918 2949
rect 52970 2937 52976 2949
rect 53680 2937 53686 2949
rect 52970 2909 53686 2937
rect 52970 2897 52976 2909
rect 53680 2897 53686 2909
rect 53738 2897 53744 2949
rect 54832 2897 54838 2949
rect 54890 2937 54896 2949
rect 56194 2937 56222 2974
rect 54890 2909 56222 2937
rect 54890 2897 54896 2909
rect 8755 2866 8813 2872
rect 8755 2832 8767 2866
rect 8801 2863 8813 2866
rect 8801 2835 40334 2863
rect 8801 2832 8813 2835
rect 8755 2826 8813 2832
rect 16051 2792 16109 2798
rect 16051 2758 16063 2792
rect 16097 2789 16109 2792
rect 16816 2789 16822 2801
rect 16097 2761 16822 2789
rect 16097 2758 16109 2761
rect 16051 2752 16109 2758
rect 16816 2749 16822 2761
rect 16874 2749 16880 2801
rect 27760 2749 27766 2801
rect 27818 2789 27824 2801
rect 27952 2789 27958 2801
rect 27818 2761 27958 2789
rect 27818 2749 27824 2761
rect 27952 2749 27958 2761
rect 28010 2749 28016 2801
rect 32944 2789 32950 2801
rect 32905 2761 32950 2789
rect 32944 2749 32950 2761
rect 33002 2749 33008 2801
rect 40306 2789 40334 2835
rect 50032 2823 50038 2875
rect 50090 2823 50096 2875
rect 52816 2789 52822 2801
rect 40306 2761 52822 2789
rect 52816 2749 52822 2761
rect 52874 2749 52880 2801
rect 54448 2789 54454 2801
rect 54409 2761 54454 2789
rect 54448 2749 54454 2761
rect 54506 2749 54512 2801
rect 1152 2690 58848 2712
rect 1152 2638 4294 2690
rect 4346 2638 4358 2690
rect 4410 2638 4422 2690
rect 4474 2638 4486 2690
rect 4538 2638 35014 2690
rect 35066 2638 35078 2690
rect 35130 2638 35142 2690
rect 35194 2638 35206 2690
rect 35258 2638 58848 2690
rect 1152 2616 58848 2638
rect 3952 2527 3958 2579
rect 4010 2567 4016 2579
rect 4240 2567 4246 2579
rect 4010 2539 4246 2567
rect 4010 2527 4016 2539
rect 4240 2527 4246 2539
rect 4298 2527 4304 2579
rect 4336 2527 4342 2579
rect 4394 2567 4400 2579
rect 4816 2567 4822 2579
rect 4394 2539 4822 2567
rect 4394 2527 4400 2539
rect 4816 2527 4822 2539
rect 4874 2527 4880 2579
rect 7984 2527 7990 2579
rect 8042 2567 8048 2579
rect 32944 2567 32950 2579
rect 8042 2539 32950 2567
rect 8042 2527 8048 2539
rect 32944 2527 32950 2539
rect 33002 2527 33008 2579
rect 35152 2527 35158 2579
rect 35210 2567 35216 2579
rect 35536 2567 35542 2579
rect 35210 2539 35542 2567
rect 35210 2527 35216 2539
rect 35536 2527 35542 2539
rect 35594 2527 35600 2579
rect 5776 2453 5782 2505
rect 5834 2493 5840 2505
rect 54448 2493 54454 2505
rect 5834 2465 54454 2493
rect 5834 2453 5840 2465
rect 54448 2453 54454 2465
rect 54506 2453 54512 2505
rect 20176 2379 20182 2431
rect 20234 2419 20240 2431
rect 20848 2419 20854 2431
rect 20234 2391 20854 2419
rect 20234 2379 20240 2391
rect 20848 2379 20854 2391
rect 20906 2379 20912 2431
rect 4720 2009 4726 2061
rect 4778 2049 4784 2061
rect 5296 2049 5302 2061
rect 4778 2021 5302 2049
rect 4778 2009 4784 2021
rect 5296 2009 5302 2021
rect 5354 2009 5360 2061
rect 4528 1861 4534 1913
rect 4586 1901 4592 1913
rect 4816 1901 4822 1913
rect 4586 1873 4822 1901
rect 4586 1861 4592 1873
rect 4816 1861 4822 1873
rect 4874 1861 4880 1913
rect 30352 1713 30358 1765
rect 30410 1753 30416 1765
rect 31504 1753 31510 1765
rect 30410 1725 31510 1753
rect 30410 1713 30416 1725
rect 31504 1713 31510 1725
rect 31562 1713 31568 1765
rect 34864 1713 34870 1765
rect 34922 1753 34928 1765
rect 35632 1753 35638 1765
rect 34922 1725 35638 1753
rect 34922 1713 34928 1725
rect 35632 1713 35638 1725
rect 35690 1713 35696 1765
rect 41008 1713 41014 1765
rect 41066 1753 41072 1765
rect 41296 1753 41302 1765
rect 41066 1725 41302 1753
rect 41066 1713 41072 1725
rect 41296 1713 41302 1725
rect 41354 1713 41360 1765
rect 54352 1713 54358 1765
rect 54410 1753 54416 1765
rect 54640 1753 54646 1765
rect 54410 1725 54646 1753
rect 54410 1713 54416 1725
rect 54640 1713 54646 1725
rect 54698 1713 54704 1765
rect 35632 1565 35638 1617
rect 35690 1605 35696 1617
rect 35920 1605 35926 1617
rect 35690 1577 35926 1605
rect 35690 1565 35696 1577
rect 35920 1565 35926 1577
rect 35978 1565 35984 1617
rect 36304 1491 36310 1543
rect 36362 1491 36368 1543
rect 50512 1491 50518 1543
rect 50570 1531 50576 1543
rect 51088 1531 51094 1543
rect 50570 1503 51094 1531
rect 50570 1491 50576 1503
rect 51088 1491 51094 1503
rect 51146 1491 51152 1543
rect 33232 1417 33238 1469
rect 33290 1457 33296 1469
rect 33712 1457 33718 1469
rect 33290 1429 33718 1457
rect 33290 1417 33296 1429
rect 33712 1417 33718 1429
rect 33770 1417 33776 1469
rect 34672 1417 34678 1469
rect 34730 1457 34736 1469
rect 35440 1457 35446 1469
rect 34730 1429 35446 1457
rect 34730 1417 34736 1429
rect 35440 1417 35446 1429
rect 35498 1417 35504 1469
rect 36322 1173 36350 1491
rect 45424 1417 45430 1469
rect 45482 1457 45488 1469
rect 45712 1457 45718 1469
rect 45482 1429 45718 1457
rect 45482 1417 45488 1429
rect 45712 1417 45718 1429
rect 45770 1417 45776 1469
rect 50704 1417 50710 1469
rect 50762 1457 50768 1469
rect 50896 1457 50902 1469
rect 50762 1429 50902 1457
rect 50762 1417 50768 1429
rect 50896 1417 50902 1429
rect 50954 1417 50960 1469
rect 43312 1269 43318 1321
rect 43370 1309 43376 1321
rect 43984 1309 43990 1321
rect 43370 1281 43990 1309
rect 43370 1269 43376 1281
rect 43984 1269 43990 1281
rect 44042 1269 44048 1321
rect 50896 1269 50902 1321
rect 50954 1309 50960 1321
rect 51568 1309 51574 1321
rect 50954 1281 51574 1309
rect 50954 1269 50960 1281
rect 51568 1269 51574 1281
rect 51626 1269 51632 1321
rect 36304 1121 36310 1173
rect 36362 1121 36368 1173
rect 45136 1047 45142 1099
rect 45194 1087 45200 1099
rect 45328 1087 45334 1099
rect 45194 1059 45334 1087
rect 45194 1047 45200 1059
rect 45328 1047 45334 1059
rect 45386 1047 45392 1099
rect 43024 899 43030 951
rect 43082 939 43088 951
rect 44368 939 44374 951
rect 43082 911 44374 939
rect 43082 899 43088 911
rect 44368 899 44374 911
rect 44426 899 44432 951
<< via1 >>
rect 4294 57250 4346 57302
rect 4358 57250 4410 57302
rect 4422 57250 4474 57302
rect 4486 57250 4538 57302
rect 35014 57250 35066 57302
rect 35078 57250 35130 57302
rect 35142 57250 35194 57302
rect 35206 57250 35258 57302
rect 1750 56991 1802 57043
rect 214 56917 266 56969
rect 3286 56991 3338 57043
rect 4918 56917 4970 56969
rect 9622 56991 9674 57043
rect 11254 56991 11306 57043
rect 6454 56917 6506 56969
rect 8086 56960 8138 56969
rect 8086 56926 8095 56960
rect 8095 56926 8129 56960
rect 8129 56926 8138 56960
rect 8086 56917 8138 56926
rect 16438 56991 16490 57043
rect 29110 56991 29162 57043
rect 12790 56917 12842 56969
rect 14422 56917 14474 56969
rect 15958 56917 16010 56969
rect 17494 56917 17546 56969
rect 19126 56917 19178 56969
rect 20662 56917 20714 56969
rect 22294 56917 22346 56969
rect 23830 56917 23882 56969
rect 25462 56917 25514 56969
rect 26998 56917 27050 56969
rect 28630 56917 28682 56969
rect 30166 56917 30218 56969
rect 31702 56960 31754 56969
rect 31702 56926 31711 56960
rect 31711 56926 31745 56960
rect 31745 56926 31754 56960
rect 31702 56917 31754 56926
rect 33334 56917 33386 56969
rect 34870 56960 34922 56969
rect 34870 56926 34879 56960
rect 34879 56926 34913 56960
rect 34913 56926 34922 56960
rect 34870 56917 34922 56926
rect 38038 56960 38090 56969
rect 38038 56926 38047 56960
rect 38047 56926 38081 56960
rect 38081 56926 38090 56960
rect 38038 56917 38090 56926
rect 41206 56917 41258 56969
rect 44374 56917 44426 56969
rect 47542 56960 47594 56969
rect 47542 56926 47551 56960
rect 47551 56926 47585 56960
rect 47585 56926 47594 56960
rect 47542 56917 47594 56926
rect 49942 56917 49994 56969
rect 52150 56917 52202 56969
rect 53878 56960 53930 56969
rect 53878 56926 53887 56960
rect 53887 56926 53921 56960
rect 53921 56926 53930 56960
rect 53878 56917 53930 56926
rect 2038 56843 2090 56895
rect 3574 56843 3626 56895
rect 5110 56886 5162 56895
rect 5110 56852 5119 56886
rect 5119 56852 5153 56886
rect 5153 56852 5162 56886
rect 5110 56843 5162 56852
rect 7222 56886 7274 56895
rect 7222 56852 7231 56886
rect 7231 56852 7265 56886
rect 7265 56852 7274 56886
rect 11254 56886 11306 56895
rect 7222 56843 7274 56852
rect 11254 56852 11263 56886
rect 11263 56852 11297 56886
rect 11297 56852 11306 56886
rect 11254 56843 11306 56852
rect 12982 56886 13034 56895
rect 12982 56852 12991 56886
rect 12991 56852 13025 56886
rect 13025 56852 13034 56886
rect 12982 56843 13034 56852
rect 16150 56886 16202 56895
rect 16150 56852 16159 56886
rect 16159 56852 16193 56886
rect 16193 56852 16202 56886
rect 16150 56843 16202 56852
rect 17974 56886 18026 56895
rect 17974 56852 17983 56886
rect 17983 56852 18017 56886
rect 18017 56852 18026 56886
rect 17974 56843 18026 56852
rect 19318 56886 19370 56895
rect 19318 56852 19327 56886
rect 19327 56852 19361 56886
rect 19361 56852 19370 56886
rect 19318 56843 19370 56852
rect 20854 56886 20906 56895
rect 20854 56852 20863 56886
rect 20863 56852 20897 56886
rect 20897 56852 20906 56886
rect 20854 56843 20906 56852
rect 24022 56886 24074 56895
rect 24022 56852 24031 56886
rect 24031 56852 24065 56886
rect 24065 56852 24074 56886
rect 24022 56843 24074 56852
rect 27190 56886 27242 56895
rect 27190 56852 27199 56886
rect 27199 56852 27233 56886
rect 27233 56852 27242 56886
rect 27190 56843 27242 56852
rect 28822 56886 28874 56895
rect 28822 56852 28831 56886
rect 28831 56852 28865 56886
rect 28865 56852 28874 56886
rect 28822 56843 28874 56852
rect 32566 56886 32618 56895
rect 32566 56852 32575 56886
rect 32575 56852 32609 56886
rect 32609 56852 32618 56886
rect 32566 56843 32618 56852
rect 34102 56886 34154 56895
rect 34102 56852 34111 56886
rect 34111 56852 34145 56886
rect 34145 56852 34154 56886
rect 34102 56843 34154 56852
rect 36502 56843 36554 56895
rect 39670 56843 39722 56895
rect 26710 56769 26762 56821
rect 42838 56843 42890 56895
rect 45910 56843 45962 56895
rect 49078 56843 49130 56895
rect 50710 56843 50762 56895
rect 52246 56843 52298 56895
rect 55414 56843 55466 56895
rect 57046 56886 57098 56895
rect 57046 56852 57055 56886
rect 57055 56852 57089 56886
rect 57089 56852 57098 56886
rect 57046 56843 57098 56852
rect 47926 56769 47978 56821
rect 54838 56769 54890 56821
rect 9814 56738 9866 56747
rect 9814 56704 9823 56738
rect 9823 56704 9857 56738
rect 9857 56704 9866 56738
rect 9814 56695 9866 56704
rect 36694 56738 36746 56747
rect 36694 56704 36703 56738
rect 36703 56704 36737 56738
rect 36737 56704 36746 56738
rect 36694 56695 36746 56704
rect 39766 56738 39818 56747
rect 39766 56704 39775 56738
rect 39775 56704 39809 56738
rect 39809 56704 39818 56738
rect 39766 56695 39818 56704
rect 40438 56738 40490 56747
rect 40438 56704 40447 56738
rect 40447 56704 40481 56738
rect 40481 56704 40490 56738
rect 40438 56695 40490 56704
rect 40822 56738 40874 56747
rect 40822 56704 40831 56738
rect 40831 56704 40865 56738
rect 40865 56704 40874 56738
rect 40822 56695 40874 56704
rect 42934 56738 42986 56747
rect 42934 56704 42943 56738
rect 42943 56704 42977 56738
rect 42977 56704 42986 56738
rect 42934 56695 42986 56704
rect 46102 56695 46154 56747
rect 48694 56738 48746 56747
rect 48694 56704 48703 56738
rect 48703 56704 48737 56738
rect 48737 56704 48746 56738
rect 48694 56695 48746 56704
rect 50806 56738 50858 56747
rect 50806 56704 50815 56738
rect 50815 56704 50849 56738
rect 50849 56704 50858 56738
rect 50806 56695 50858 56704
rect 52822 56738 52874 56747
rect 52822 56704 52831 56738
rect 52831 56704 52865 56738
rect 52865 56704 52874 56738
rect 52822 56695 52874 56704
rect 55414 56695 55466 56747
rect 56758 56738 56810 56747
rect 56758 56704 56767 56738
rect 56767 56704 56801 56738
rect 56801 56704 56810 56738
rect 56758 56695 56810 56704
rect 19654 56584 19706 56636
rect 19718 56584 19770 56636
rect 19782 56584 19834 56636
rect 19846 56584 19898 56636
rect 50374 56584 50426 56636
rect 50438 56584 50490 56636
rect 50502 56584 50554 56636
rect 50566 56584 50618 56636
rect 694 56473 746 56525
rect 2230 56473 2282 56525
rect 2806 56473 2858 56525
rect 3862 56473 3914 56525
rect 5398 56473 5450 56525
rect 5974 56473 6026 56525
rect 7030 56473 7082 56525
rect 8566 56473 8618 56525
rect 10198 56473 10250 56525
rect 10678 56473 10730 56525
rect 11734 56473 11786 56525
rect 12310 56473 12362 56525
rect 13366 56473 13418 56525
rect 14902 56473 14954 56525
rect 17014 56473 17066 56525
rect 18070 56473 18122 56525
rect 18742 56473 18794 56525
rect 21238 56473 21290 56525
rect 21718 56473 21770 56525
rect 22774 56473 22826 56525
rect 24406 56516 24458 56525
rect 24406 56482 24415 56516
rect 24415 56482 24449 56516
rect 24449 56482 24458 56516
rect 24406 56473 24458 56482
rect 25942 56473 25994 56525
rect 26518 56473 26570 56525
rect 27574 56473 27626 56525
rect 28054 56473 28106 56525
rect 29686 56516 29738 56525
rect 29686 56482 29695 56516
rect 29695 56482 29729 56516
rect 29729 56482 29738 56516
rect 29686 56473 29738 56482
rect 30646 56473 30698 56525
rect 32278 56473 32330 56525
rect 33814 56473 33866 56525
rect 34390 56473 34442 56525
rect 36022 56473 36074 56525
rect 37558 56473 37610 56525
rect 38614 56473 38666 56525
rect 40150 56516 40202 56525
rect 40150 56482 40159 56516
rect 40159 56482 40193 56516
rect 40193 56482 40202 56516
rect 40150 56473 40202 56482
rect 41782 56473 41834 56525
rect 42262 56473 42314 56525
rect 43318 56473 43370 56525
rect 43894 56473 43946 56525
rect 44950 56473 45002 56525
rect 46486 56473 46538 56525
rect 48022 56473 48074 56525
rect 49654 56473 49706 56525
rect 50134 56473 50186 56525
rect 52918 56516 52970 56525
rect 52918 56482 52927 56516
rect 52927 56482 52961 56516
rect 52961 56482 52970 56516
rect 52918 56473 52970 56482
rect 53302 56473 53354 56525
rect 54358 56473 54410 56525
rect 54934 56473 54986 56525
rect 55990 56516 56042 56525
rect 55990 56482 55999 56516
rect 55999 56482 56033 56516
rect 56033 56482 56042 56516
rect 55990 56473 56042 56482
rect 16534 56399 16586 56451
rect 56758 56399 56810 56451
rect 13750 56325 13802 56377
rect 43318 56325 43370 56377
rect 3766 56251 3818 56303
rect 15190 56251 15242 56303
rect 26422 56251 26474 56303
rect 36022 56251 36074 56303
rect 1750 56220 1802 56229
rect 1750 56186 1759 56220
rect 1759 56186 1793 56220
rect 1793 56186 1802 56220
rect 1750 56177 1802 56186
rect 2518 56220 2570 56229
rect 2518 56186 2527 56220
rect 2527 56186 2561 56220
rect 2561 56186 2570 56220
rect 2518 56177 2570 56186
rect 3382 56177 3434 56229
rect 5206 56177 5258 56229
rect 5590 56220 5642 56229
rect 5590 56186 5599 56220
rect 5599 56186 5633 56220
rect 5633 56186 5642 56220
rect 5590 56177 5642 56186
rect 6358 56220 6410 56229
rect 6358 56186 6367 56220
rect 6367 56186 6401 56220
rect 6401 56186 6410 56220
rect 6358 56177 6410 56186
rect 6454 56177 6506 56229
rect 10774 56220 10826 56229
rect 10774 56186 10783 56220
rect 10783 56186 10817 56220
rect 10817 56186 10826 56220
rect 10774 56177 10826 56186
rect 11926 56220 11978 56229
rect 11926 56186 11935 56220
rect 11935 56186 11969 56220
rect 11969 56186 11978 56220
rect 11926 56177 11978 56186
rect 12694 56220 12746 56229
rect 12694 56186 12703 56220
rect 12703 56186 12737 56220
rect 12737 56186 12746 56220
rect 12694 56177 12746 56186
rect 15094 56220 15146 56229
rect 15094 56186 15103 56220
rect 15103 56186 15137 56220
rect 15137 56186 15146 56220
rect 15094 56177 15146 56186
rect 15766 56220 15818 56229
rect 15766 56186 15775 56220
rect 15775 56186 15809 56220
rect 15809 56186 15818 56220
rect 15766 56177 15818 56186
rect 15382 56103 15434 56155
rect 16630 56177 16682 56229
rect 18262 56220 18314 56229
rect 18262 56186 18271 56220
rect 18271 56186 18305 56220
rect 18305 56186 18314 56220
rect 18262 56177 18314 56186
rect 18742 56220 18794 56229
rect 18742 56186 18751 56220
rect 18751 56186 18785 56220
rect 18785 56186 18794 56220
rect 18742 56177 18794 56186
rect 19990 56220 20042 56229
rect 19990 56186 19999 56220
rect 19999 56186 20033 56220
rect 20033 56186 20042 56220
rect 19990 56177 20042 56186
rect 21046 56220 21098 56229
rect 19510 56103 19562 56155
rect 21046 56186 21055 56220
rect 21055 56186 21089 56220
rect 21089 56186 21098 56220
rect 21046 56177 21098 56186
rect 21814 56220 21866 56229
rect 21814 56186 21823 56220
rect 21823 56186 21857 56220
rect 21857 56186 21866 56220
rect 21814 56177 21866 56186
rect 22966 56220 23018 56229
rect 22966 56186 22975 56220
rect 22975 56186 23009 56220
rect 23009 56186 23018 56220
rect 22966 56177 23018 56186
rect 24310 56220 24362 56229
rect 24310 56186 24319 56220
rect 24319 56186 24353 56220
rect 24353 56186 24362 56220
rect 24310 56177 24362 56186
rect 26518 56220 26570 56229
rect 26518 56186 26527 56220
rect 26527 56186 26561 56220
rect 26561 56186 26570 56220
rect 26518 56177 26570 56186
rect 27670 56220 27722 56229
rect 27670 56186 27679 56220
rect 27679 56186 27713 56220
rect 27713 56186 27722 56220
rect 27670 56177 27722 56186
rect 28150 56220 28202 56229
rect 28150 56186 28159 56220
rect 28159 56186 28193 56220
rect 28193 56186 28202 56220
rect 28150 56177 28202 56186
rect 29590 56220 29642 56229
rect 29590 56186 29599 56220
rect 29599 56186 29633 56220
rect 29633 56186 29642 56220
rect 29590 56177 29642 56186
rect 30934 56220 30986 56229
rect 30934 56186 30943 56220
rect 30943 56186 30977 56220
rect 30977 56186 30986 56220
rect 30934 56177 30986 56186
rect 31318 56220 31370 56229
rect 31318 56186 31327 56220
rect 31327 56186 31361 56220
rect 31361 56186 31370 56220
rect 31318 56177 31370 56186
rect 32470 56220 32522 56229
rect 31222 56103 31274 56155
rect 32470 56186 32479 56220
rect 32479 56186 32513 56220
rect 32513 56186 32522 56220
rect 32470 56177 32522 56186
rect 32854 56220 32906 56229
rect 32854 56186 32863 56220
rect 32863 56186 32897 56220
rect 32897 56186 32906 56220
rect 32854 56177 32906 56186
rect 34006 56220 34058 56229
rect 32758 56103 32810 56155
rect 34006 56186 34015 56220
rect 34015 56186 34049 56220
rect 34049 56186 34058 56220
rect 34006 56177 34058 56186
rect 34774 56220 34826 56229
rect 34774 56186 34783 56220
rect 34783 56186 34817 56220
rect 34817 56186 34826 56220
rect 34774 56177 34826 56186
rect 35830 56220 35882 56229
rect 35830 56186 35839 56220
rect 35839 56186 35873 56220
rect 35873 56186 35882 56220
rect 35830 56177 35882 56186
rect 36598 56220 36650 56229
rect 35446 56103 35498 56155
rect 36598 56186 36607 56220
rect 36607 56186 36641 56220
rect 36641 56186 36650 56220
rect 36598 56177 36650 56186
rect 40246 56220 40298 56229
rect 40246 56186 40255 56220
rect 40255 56186 40289 56220
rect 40289 56186 40298 56220
rect 40246 56177 40298 56186
rect 42070 56177 42122 56229
rect 42358 56220 42410 56229
rect 42358 56186 42367 56220
rect 42367 56186 42401 56220
rect 42401 56186 42410 56220
rect 42358 56177 42410 56186
rect 43414 56220 43466 56229
rect 43414 56186 43423 56220
rect 43423 56186 43457 56220
rect 43457 56186 43466 56220
rect 43414 56177 43466 56186
rect 46678 56220 46730 56229
rect 46678 56186 46687 56220
rect 46687 56186 46721 56220
rect 46721 56186 46730 56220
rect 46678 56177 46730 56186
rect 46870 56251 46922 56303
rect 49174 56325 49226 56377
rect 52150 56325 52202 56377
rect 47926 56177 47978 56229
rect 48214 56220 48266 56229
rect 48214 56186 48223 56220
rect 48223 56186 48257 56220
rect 48257 56186 48266 56220
rect 48214 56177 48266 56186
rect 48886 56220 48938 56229
rect 48886 56186 48895 56220
rect 48895 56186 48929 56220
rect 48929 56186 48938 56220
rect 48886 56177 48938 56186
rect 49654 56251 49706 56303
rect 37078 56103 37130 56155
rect 40822 56103 40874 56155
rect 48598 56103 48650 56155
rect 49846 56220 49898 56229
rect 49846 56186 49855 56220
rect 49855 56186 49889 56220
rect 49889 56186 49898 56220
rect 54358 56251 54410 56303
rect 58582 56251 58634 56303
rect 49846 56177 49898 56186
rect 53014 56220 53066 56229
rect 51190 56103 51242 56155
rect 53014 56186 53023 56220
rect 53023 56186 53057 56220
rect 53057 56186 53066 56220
rect 53014 56177 53066 56186
rect 53398 56220 53450 56229
rect 53398 56186 53407 56220
rect 53407 56186 53441 56220
rect 53441 56186 53450 56220
rect 53398 56177 53450 56186
rect 54454 56220 54506 56229
rect 54454 56186 54463 56220
rect 54463 56186 54497 56220
rect 54497 56186 54506 56220
rect 54454 56177 54506 56186
rect 55510 56220 55562 56229
rect 55510 56186 55519 56220
rect 55519 56186 55553 56220
rect 55553 56186 55562 56220
rect 55510 56177 55562 56186
rect 4294 55918 4346 55970
rect 4358 55918 4410 55970
rect 4422 55918 4474 55970
rect 4486 55918 4538 55970
rect 35014 55918 35066 55970
rect 35078 55918 35130 55970
rect 35142 55918 35194 55970
rect 35206 55918 35258 55970
rect 26326 55733 26378 55785
rect 1174 55659 1226 55711
rect 4630 55659 4682 55711
rect 7510 55659 7562 55711
rect 9142 55659 9194 55711
rect 13846 55659 13898 55711
rect 20182 55659 20234 55711
rect 23350 55659 23402 55711
rect 24886 55659 24938 55711
rect 39094 55659 39146 55711
rect 40726 55659 40778 55711
rect 45430 55659 45482 55711
rect 46966 55659 47018 55711
rect 51766 55659 51818 55711
rect 56470 55659 56522 55711
rect 57526 55659 57578 55711
rect 36022 55585 36074 55637
rect 4630 55511 4682 55563
rect 7702 55554 7754 55563
rect 7702 55520 7711 55554
rect 7711 55520 7745 55554
rect 7745 55520 7754 55554
rect 7702 55511 7754 55520
rect 8470 55554 8522 55563
rect 8470 55520 8479 55554
rect 8479 55520 8513 55554
rect 8513 55520 8522 55554
rect 8470 55511 8522 55520
rect 9238 55554 9290 55563
rect 9238 55520 9247 55554
rect 9247 55520 9281 55554
rect 9281 55520 9290 55554
rect 9238 55511 9290 55520
rect 14038 55554 14090 55563
rect 14038 55520 14047 55554
rect 14047 55520 14081 55554
rect 14081 55520 14090 55554
rect 14038 55511 14090 55520
rect 20470 55511 20522 55563
rect 23446 55554 23498 55563
rect 23446 55520 23455 55554
rect 23455 55520 23489 55554
rect 23489 55520 23498 55554
rect 23446 55511 23498 55520
rect 1846 55363 1898 55415
rect 24694 55406 24746 55415
rect 24694 55372 24703 55406
rect 24703 55372 24737 55406
rect 24737 55372 24746 55406
rect 24694 55363 24746 55372
rect 28630 55363 28682 55415
rect 38902 55511 38954 55563
rect 40918 55554 40970 55563
rect 40918 55520 40927 55554
rect 40927 55520 40961 55554
rect 40961 55520 40970 55554
rect 40918 55511 40970 55520
rect 45238 55511 45290 55563
rect 46486 55511 46538 55563
rect 32374 55437 32426 55489
rect 29782 55406 29834 55415
rect 29782 55372 29791 55406
rect 29791 55372 29825 55406
rect 29825 55372 29834 55406
rect 29782 55363 29834 55372
rect 38902 55406 38954 55415
rect 38902 55372 38911 55406
rect 38911 55372 38945 55406
rect 38945 55372 38954 55406
rect 38902 55363 38954 55372
rect 45238 55406 45290 55415
rect 45238 55372 45247 55406
rect 45247 55372 45281 55406
rect 45281 55372 45290 55406
rect 45238 55363 45290 55372
rect 46486 55363 46538 55415
rect 56662 55554 56714 55563
rect 56662 55520 56671 55554
rect 56671 55520 56705 55554
rect 56705 55520 56714 55554
rect 56662 55511 56714 55520
rect 57526 55511 57578 55563
rect 50710 55363 50762 55415
rect 51574 55406 51626 55415
rect 51574 55372 51583 55406
rect 51583 55372 51617 55406
rect 51617 55372 51626 55406
rect 51574 55363 51626 55372
rect 55606 55406 55658 55415
rect 55606 55372 55615 55406
rect 55615 55372 55649 55406
rect 55649 55372 55658 55406
rect 55606 55363 55658 55372
rect 19654 55252 19706 55304
rect 19718 55252 19770 55304
rect 19782 55252 19834 55304
rect 19846 55252 19898 55304
rect 50374 55252 50426 55304
rect 50438 55252 50490 55304
rect 50502 55252 50554 55304
rect 50566 55252 50618 55304
rect 12022 55141 12074 55193
rect 24694 55141 24746 55193
rect 26710 55184 26762 55193
rect 26710 55150 26719 55184
rect 26719 55150 26753 55184
rect 26753 55150 26762 55184
rect 26710 55141 26762 55150
rect 59158 55141 59210 55193
rect 30166 55067 30218 55119
rect 55606 55067 55658 55119
rect 20566 54993 20618 55045
rect 32374 54993 32426 55045
rect 54358 54993 54410 55045
rect 5302 54919 5354 54971
rect 28630 54919 28682 54971
rect 36790 54962 36842 54971
rect 36790 54928 36799 54962
rect 36799 54928 36833 54962
rect 36833 54928 36842 54962
rect 36790 54919 36842 54928
rect 57910 54888 57962 54897
rect 8470 54771 8522 54823
rect 57910 54854 57919 54888
rect 57919 54854 57953 54888
rect 57953 54854 57962 54888
rect 57910 54845 57962 54854
rect 51094 54771 51146 54823
rect 40918 54697 40970 54749
rect 46582 54740 46634 54749
rect 46582 54706 46591 54740
rect 46591 54706 46625 54740
rect 46625 54706 46634 54740
rect 46582 54697 46634 54706
rect 4294 54586 4346 54638
rect 4358 54586 4410 54638
rect 4422 54586 4474 54638
rect 4486 54586 4538 54638
rect 35014 54586 35066 54638
rect 35078 54586 35130 54638
rect 35142 54586 35194 54638
rect 35206 54586 35258 54638
rect 58102 54327 58154 54379
rect 33622 54179 33674 54231
rect 2134 54105 2186 54157
rect 49750 54179 49802 54231
rect 34006 54031 34058 54083
rect 57622 54074 57674 54083
rect 57622 54040 57631 54074
rect 57631 54040 57665 54074
rect 57665 54040 57674 54074
rect 57622 54031 57674 54040
rect 19654 53920 19706 53972
rect 19718 53920 19770 53972
rect 19782 53920 19834 53972
rect 19846 53920 19898 53972
rect 50374 53920 50426 53972
rect 50438 53920 50490 53972
rect 50502 53920 50554 53972
rect 50566 53920 50618 53972
rect 59638 53809 59690 53861
rect 26134 53439 26186 53491
rect 57334 53365 57386 53417
rect 57718 53365 57770 53417
rect 4294 53254 4346 53306
rect 4358 53254 4410 53306
rect 4422 53254 4474 53306
rect 4486 53254 4538 53306
rect 35014 53254 35066 53306
rect 35078 53254 35130 53306
rect 35142 53254 35194 53306
rect 35206 53254 35258 53306
rect 3286 52847 3338 52899
rect 25078 52847 25130 52899
rect 23542 52699 23594 52751
rect 19654 52588 19706 52640
rect 19718 52588 19770 52640
rect 19782 52588 19834 52640
rect 19846 52588 19898 52640
rect 50374 52588 50426 52640
rect 50438 52588 50490 52640
rect 50502 52588 50554 52640
rect 50566 52588 50618 52640
rect 11926 52181 11978 52233
rect 4294 51922 4346 51974
rect 4358 51922 4410 51974
rect 4422 51922 4474 51974
rect 4486 51922 4538 51974
rect 35014 51922 35066 51974
rect 35078 51922 35130 51974
rect 35142 51922 35194 51974
rect 35206 51922 35258 51974
rect 23062 51515 23114 51567
rect 19654 51256 19706 51308
rect 19718 51256 19770 51308
rect 19782 51256 19834 51308
rect 19846 51256 19898 51308
rect 50374 51256 50426 51308
rect 50438 51256 50490 51308
rect 50502 51256 50554 51308
rect 50566 51256 50618 51308
rect 57910 50997 57962 51049
rect 1750 50849 1802 50901
rect 9430 50744 9482 50753
rect 9430 50710 9439 50744
rect 9439 50710 9473 50744
rect 9473 50710 9482 50744
rect 9430 50701 9482 50710
rect 50230 50701 50282 50753
rect 4294 50590 4346 50642
rect 4358 50590 4410 50642
rect 4422 50590 4474 50642
rect 4486 50590 4538 50642
rect 35014 50590 35066 50642
rect 35078 50590 35130 50642
rect 35142 50590 35194 50642
rect 35206 50590 35258 50642
rect 54838 50479 54890 50531
rect 10294 50448 10346 50457
rect 10294 50414 10303 50448
rect 10303 50414 10337 50448
rect 10337 50414 10346 50448
rect 10294 50405 10346 50414
rect 19654 49924 19706 49976
rect 19718 49924 19770 49976
rect 19782 49924 19834 49976
rect 19846 49924 19898 49976
rect 50374 49924 50426 49976
rect 50438 49924 50490 49976
rect 50502 49924 50554 49976
rect 50566 49924 50618 49976
rect 10294 49665 10346 49717
rect 29110 49665 29162 49717
rect 47542 49443 47594 49495
rect 33238 49412 33290 49421
rect 33238 49378 33247 49412
rect 33247 49378 33281 49412
rect 33281 49378 33290 49412
rect 33238 49369 33290 49378
rect 44182 49412 44234 49421
rect 44182 49378 44191 49412
rect 44191 49378 44225 49412
rect 44225 49378 44234 49412
rect 44182 49369 44234 49378
rect 4294 49258 4346 49310
rect 4358 49258 4410 49310
rect 4422 49258 4474 49310
rect 4486 49258 4538 49310
rect 35014 49258 35066 49310
rect 35078 49258 35130 49310
rect 35142 49258 35194 49310
rect 35206 49258 35258 49310
rect 9046 49147 9098 49199
rect 44182 49147 44234 49199
rect 27286 49073 27338 49125
rect 33238 49073 33290 49125
rect 39478 48851 39530 48903
rect 19654 48592 19706 48644
rect 19718 48592 19770 48644
rect 19782 48592 19834 48644
rect 19846 48592 19898 48644
rect 50374 48592 50426 48644
rect 50438 48592 50490 48644
rect 50502 48592 50554 48644
rect 50566 48592 50618 48644
rect 2710 48080 2762 48089
rect 2710 48046 2719 48080
rect 2719 48046 2753 48080
rect 2753 48046 2762 48080
rect 2710 48037 2762 48046
rect 37750 48037 37802 48089
rect 4294 47926 4346 47978
rect 4358 47926 4410 47978
rect 4422 47926 4474 47978
rect 4486 47926 4538 47978
rect 35014 47926 35066 47978
rect 35078 47926 35130 47978
rect 35142 47926 35194 47978
rect 35206 47926 35258 47978
rect 2710 47815 2762 47867
rect 56950 47815 57002 47867
rect 28342 47519 28394 47571
rect 49174 47488 49226 47497
rect 49174 47454 49183 47488
rect 49183 47454 49217 47488
rect 49217 47454 49226 47488
rect 49174 47445 49226 47454
rect 19654 47260 19706 47312
rect 19718 47260 19770 47312
rect 19782 47260 19834 47312
rect 19846 47260 19898 47312
rect 50374 47260 50426 47312
rect 50438 47260 50490 47312
rect 50502 47260 50554 47312
rect 50566 47260 50618 47312
rect 48214 47001 48266 47053
rect 36406 46748 36458 46757
rect 36406 46714 36415 46748
rect 36415 46714 36449 46748
rect 36449 46714 36458 46748
rect 36406 46705 36458 46714
rect 4294 46594 4346 46646
rect 4358 46594 4410 46646
rect 4422 46594 4474 46646
rect 4486 46594 4538 46646
rect 35014 46594 35066 46646
rect 35078 46594 35130 46646
rect 35142 46594 35194 46646
rect 35206 46594 35258 46646
rect 54646 46113 54698 46165
rect 19654 45928 19706 45980
rect 19718 45928 19770 45980
rect 19782 45928 19834 45980
rect 19846 45928 19898 45980
rect 50374 45928 50426 45980
rect 50438 45928 50490 45980
rect 50502 45928 50554 45980
rect 50566 45928 50618 45980
rect 7702 45447 7754 45499
rect 12598 45416 12650 45425
rect 12598 45382 12607 45416
rect 12607 45382 12641 45416
rect 12641 45382 12650 45416
rect 12598 45373 12650 45382
rect 48790 45416 48842 45425
rect 48790 45382 48799 45416
rect 48799 45382 48833 45416
rect 48833 45382 48842 45416
rect 48790 45373 48842 45382
rect 55606 45373 55658 45425
rect 4294 45262 4346 45314
rect 4358 45262 4410 45314
rect 4422 45262 4474 45314
rect 4486 45262 4538 45314
rect 35014 45262 35066 45314
rect 35078 45262 35130 45314
rect 35142 45262 35194 45314
rect 35206 45262 35258 45314
rect 31798 45151 31850 45203
rect 48790 45151 48842 45203
rect 29014 44707 29066 44759
rect 19654 44596 19706 44648
rect 19718 44596 19770 44648
rect 19782 44596 19834 44648
rect 19846 44596 19898 44648
rect 50374 44596 50426 44648
rect 50438 44596 50490 44648
rect 50502 44596 50554 44648
rect 50566 44596 50618 44648
rect 41110 44041 41162 44093
rect 42262 44041 42314 44093
rect 52150 44084 52202 44093
rect 52150 44050 52159 44084
rect 52159 44050 52193 44084
rect 52193 44050 52202 44084
rect 52150 44041 52202 44050
rect 4294 43930 4346 43982
rect 4358 43930 4410 43982
rect 4422 43930 4474 43982
rect 4486 43930 4538 43982
rect 35014 43930 35066 43982
rect 35078 43930 35130 43982
rect 35142 43930 35194 43982
rect 35206 43930 35258 43982
rect 49558 43745 49610 43797
rect 34582 43671 34634 43723
rect 56086 43597 56138 43649
rect 23926 43449 23978 43501
rect 19654 43264 19706 43316
rect 19718 43264 19770 43316
rect 19782 43264 19834 43316
rect 19846 43264 19898 43316
rect 50374 43264 50426 43316
rect 50438 43264 50490 43316
rect 50502 43264 50554 43316
rect 50566 43264 50618 43316
rect 16438 42752 16490 42761
rect 16438 42718 16447 42752
rect 16447 42718 16481 42752
rect 16481 42718 16490 42752
rect 16438 42709 16490 42718
rect 20086 42752 20138 42761
rect 20086 42718 20095 42752
rect 20095 42718 20129 42752
rect 20129 42718 20138 42752
rect 20086 42709 20138 42718
rect 21142 42709 21194 42761
rect 52534 42752 52586 42761
rect 52534 42718 52543 42752
rect 52543 42718 52577 42752
rect 52577 42718 52586 42752
rect 52534 42709 52586 42718
rect 4294 42598 4346 42650
rect 4358 42598 4410 42650
rect 4422 42598 4474 42650
rect 4486 42598 4538 42650
rect 35014 42598 35066 42650
rect 35078 42598 35130 42650
rect 35142 42598 35194 42650
rect 35206 42598 35258 42650
rect 16438 42487 16490 42539
rect 27766 42487 27818 42539
rect 16726 42191 16778 42243
rect 3670 42043 3722 42095
rect 45334 42043 45386 42095
rect 19654 41932 19706 41984
rect 19718 41932 19770 41984
rect 19782 41932 19834 41984
rect 19846 41932 19898 41984
rect 50374 41932 50426 41984
rect 50438 41932 50490 41984
rect 50502 41932 50554 41984
rect 50566 41932 50618 41984
rect 4294 41266 4346 41318
rect 4358 41266 4410 41318
rect 4422 41266 4474 41318
rect 4486 41266 4538 41318
rect 35014 41266 35066 41318
rect 35078 41266 35130 41318
rect 35142 41266 35194 41318
rect 35206 41266 35258 41318
rect 33334 40859 33386 40911
rect 18838 40785 18890 40837
rect 33334 40711 33386 40763
rect 40246 40711 40298 40763
rect 19654 40600 19706 40652
rect 19718 40600 19770 40652
rect 19782 40600 19834 40652
rect 19846 40600 19898 40652
rect 50374 40600 50426 40652
rect 50438 40600 50490 40652
rect 50502 40600 50554 40652
rect 50566 40600 50618 40652
rect 15190 40489 15242 40541
rect 15958 40045 16010 40097
rect 23350 40088 23402 40097
rect 23350 40054 23359 40088
rect 23359 40054 23393 40088
rect 23393 40054 23402 40088
rect 23350 40045 23402 40054
rect 47254 40088 47306 40097
rect 47254 40054 47263 40088
rect 47263 40054 47297 40088
rect 47297 40054 47306 40088
rect 47254 40045 47306 40054
rect 4294 39934 4346 39986
rect 4358 39934 4410 39986
rect 4422 39934 4474 39986
rect 4486 39934 4538 39986
rect 35014 39934 35066 39986
rect 35078 39934 35130 39986
rect 35142 39934 35194 39986
rect 35206 39934 35258 39986
rect 15862 39823 15914 39875
rect 47254 39823 47306 39875
rect 49462 39527 49514 39579
rect 52918 39527 52970 39579
rect 19654 39268 19706 39320
rect 19718 39268 19770 39320
rect 19782 39268 19834 39320
rect 19846 39268 19898 39320
rect 50374 39268 50426 39320
rect 50438 39268 50490 39320
rect 50502 39268 50554 39320
rect 50566 39268 50618 39320
rect 22966 38713 23018 38765
rect 38710 38713 38762 38765
rect 4294 38602 4346 38654
rect 4358 38602 4410 38654
rect 4422 38602 4474 38654
rect 4486 38602 4538 38654
rect 35014 38602 35066 38654
rect 35078 38602 35130 38654
rect 35142 38602 35194 38654
rect 35206 38602 35258 38654
rect 6358 38195 6410 38247
rect 20470 38195 20522 38247
rect 19654 37936 19706 37988
rect 19718 37936 19770 37988
rect 19782 37936 19834 37988
rect 19846 37936 19898 37988
rect 50374 37936 50426 37988
rect 50438 37936 50490 37988
rect 50502 37936 50554 37988
rect 50566 37936 50618 37988
rect 51190 37455 51242 37507
rect 2422 37381 2474 37433
rect 6454 37381 6506 37433
rect 47350 37381 47402 37433
rect 4294 37270 4346 37322
rect 4358 37270 4410 37322
rect 4422 37270 4474 37322
rect 4486 37270 4538 37322
rect 35014 37270 35066 37322
rect 35078 37270 35130 37322
rect 35142 37270 35194 37322
rect 35206 37270 35258 37322
rect 2518 37011 2570 37063
rect 23734 37011 23786 37063
rect 28246 36906 28298 36915
rect 28246 36872 28255 36906
rect 28255 36872 28289 36906
rect 28289 36872 28298 36906
rect 28246 36863 28298 36872
rect 51574 36937 51626 36989
rect 49846 36715 49898 36767
rect 19654 36604 19706 36656
rect 19718 36604 19770 36656
rect 19782 36604 19834 36656
rect 19846 36604 19898 36656
rect 50374 36604 50426 36656
rect 50438 36604 50490 36656
rect 50502 36604 50554 36656
rect 50566 36604 50618 36656
rect 28246 36493 28298 36545
rect 45430 36493 45482 36545
rect 13942 36271 13994 36323
rect 5590 36197 5642 36249
rect 31030 36197 31082 36249
rect 37174 36271 37226 36323
rect 51286 36197 51338 36249
rect 43894 36123 43946 36175
rect 24118 36049 24170 36101
rect 37174 36049 37226 36101
rect 4294 35938 4346 35990
rect 4358 35938 4410 35990
rect 4422 35938 4474 35990
rect 4486 35938 4538 35990
rect 35014 35938 35066 35990
rect 35078 35938 35130 35990
rect 35142 35938 35194 35990
rect 35206 35938 35258 35990
rect 49942 35679 49994 35731
rect 48598 35531 48650 35583
rect 19654 35272 19706 35324
rect 19718 35272 19770 35324
rect 19782 35272 19834 35324
rect 19846 35272 19898 35324
rect 50374 35272 50426 35324
rect 50438 35272 50490 35324
rect 50502 35272 50554 35324
rect 50566 35272 50618 35324
rect 33718 34791 33770 34843
rect 11350 34717 11402 34769
rect 4294 34606 4346 34658
rect 4358 34606 4410 34658
rect 4422 34606 4474 34658
rect 4486 34606 4538 34658
rect 35014 34606 35066 34658
rect 35078 34606 35130 34658
rect 35142 34606 35194 34658
rect 35206 34606 35258 34658
rect 26998 34347 27050 34399
rect 9910 34242 9962 34251
rect 9910 34208 9919 34242
rect 9919 34208 9953 34242
rect 9953 34208 9962 34242
rect 9910 34199 9962 34208
rect 49942 34199 49994 34251
rect 48790 34051 48842 34103
rect 19654 33940 19706 33992
rect 19718 33940 19770 33992
rect 19782 33940 19834 33992
rect 19846 33940 19898 33992
rect 50374 33940 50426 33992
rect 50438 33940 50490 33992
rect 50502 33940 50554 33992
rect 50566 33940 50618 33992
rect 42070 33681 42122 33733
rect 31702 33607 31754 33659
rect 34774 33533 34826 33585
rect 44950 33533 45002 33585
rect 35350 33459 35402 33511
rect 27862 33385 27914 33437
rect 34678 33428 34730 33437
rect 34678 33394 34687 33428
rect 34687 33394 34721 33428
rect 34721 33394 34730 33428
rect 34678 33385 34730 33394
rect 38230 33428 38282 33437
rect 38230 33394 38239 33428
rect 38239 33394 38273 33428
rect 38273 33394 38282 33428
rect 38230 33385 38282 33394
rect 4294 33274 4346 33326
rect 4358 33274 4410 33326
rect 4422 33274 4474 33326
rect 4486 33274 4538 33326
rect 35014 33274 35066 33326
rect 35078 33274 35130 33326
rect 35142 33274 35194 33326
rect 35206 33274 35258 33326
rect 49654 33163 49706 33215
rect 44950 33132 45002 33141
rect 44950 33098 44959 33132
rect 44959 33098 44993 33132
rect 44993 33098 45002 33132
rect 44950 33089 45002 33098
rect 22582 32719 22634 32771
rect 19654 32608 19706 32660
rect 19718 32608 19770 32660
rect 19782 32608 19834 32660
rect 19846 32608 19898 32660
rect 50374 32608 50426 32660
rect 50438 32608 50490 32660
rect 50502 32608 50554 32660
rect 50566 32608 50618 32660
rect 2326 32096 2378 32105
rect 2326 32062 2335 32096
rect 2335 32062 2369 32096
rect 2369 32062 2378 32096
rect 2326 32053 2378 32062
rect 6742 32053 6794 32105
rect 4294 31942 4346 31994
rect 4358 31942 4410 31994
rect 4422 31942 4474 31994
rect 4486 31942 4538 31994
rect 35014 31942 35066 31994
rect 35078 31942 35130 31994
rect 35142 31942 35194 31994
rect 35206 31942 35258 31994
rect 19654 31276 19706 31328
rect 19718 31276 19770 31328
rect 19782 31276 19834 31328
rect 19846 31276 19898 31328
rect 50374 31276 50426 31328
rect 50438 31276 50490 31328
rect 50502 31276 50554 31328
rect 50566 31276 50618 31328
rect 7318 30943 7370 30995
rect 43414 30943 43466 30995
rect 53014 30869 53066 30921
rect 6646 30764 6698 30773
rect 6646 30730 6655 30764
rect 6655 30730 6689 30764
rect 6689 30730 6698 30764
rect 6646 30721 6698 30730
rect 34774 30721 34826 30773
rect 49846 30721 49898 30773
rect 4294 30610 4346 30662
rect 4358 30610 4410 30662
rect 4422 30610 4474 30662
rect 4486 30610 4538 30662
rect 35014 30610 35066 30662
rect 35078 30610 35130 30662
rect 35142 30610 35194 30662
rect 35206 30610 35258 30662
rect 32182 30320 32234 30329
rect 32182 30286 32191 30320
rect 32191 30286 32225 30320
rect 32225 30286 32234 30320
rect 32182 30277 32234 30286
rect 45142 30277 45194 30329
rect 7318 30246 7370 30255
rect 7318 30212 7327 30246
rect 7327 30212 7361 30246
rect 7361 30212 7370 30246
rect 7318 30203 7370 30212
rect 19654 29944 19706 29996
rect 19718 29944 19770 29996
rect 19782 29944 19834 29996
rect 19846 29944 19898 29996
rect 50374 29944 50426 29996
rect 50438 29944 50490 29996
rect 50502 29944 50554 29996
rect 50566 29944 50618 29996
rect 9142 29389 9194 29441
rect 11158 29389 11210 29441
rect 28150 29463 28202 29515
rect 45046 29389 45098 29441
rect 4294 29278 4346 29330
rect 4358 29278 4410 29330
rect 4422 29278 4474 29330
rect 4486 29278 4538 29330
rect 35014 29278 35066 29330
rect 35078 29278 35130 29330
rect 35142 29278 35194 29330
rect 35206 29278 35258 29330
rect 24310 29167 24362 29219
rect 9142 29093 9194 29145
rect 11158 29093 11210 29145
rect 20950 29093 21002 29145
rect 15286 29019 15338 29071
rect 41302 28871 41354 28923
rect 32662 28797 32714 28849
rect 9142 28723 9194 28775
rect 19654 28612 19706 28664
rect 19718 28612 19770 28664
rect 19782 28612 19834 28664
rect 19846 28612 19898 28664
rect 50374 28612 50426 28664
rect 50438 28612 50490 28664
rect 50502 28612 50554 28664
rect 50566 28612 50618 28664
rect 9142 28501 9194 28553
rect 10870 28501 10922 28553
rect 1846 28057 1898 28109
rect 4294 27946 4346 27998
rect 4358 27946 4410 27998
rect 4422 27946 4474 27998
rect 4486 27946 4538 27998
rect 35014 27946 35066 27998
rect 35078 27946 35130 27998
rect 35142 27946 35194 27998
rect 35206 27946 35258 27998
rect 17590 27835 17642 27887
rect 15382 27613 15434 27665
rect 22966 27582 23018 27591
rect 22966 27548 22975 27582
rect 22975 27548 23009 27582
rect 23009 27548 23018 27582
rect 22966 27539 23018 27548
rect 49654 27539 49706 27591
rect 20374 27391 20426 27443
rect 19654 27280 19706 27332
rect 19718 27280 19770 27332
rect 19782 27280 19834 27332
rect 19846 27280 19898 27332
rect 50374 27280 50426 27332
rect 50438 27280 50490 27332
rect 50502 27280 50554 27332
rect 50566 27280 50618 27332
rect 8566 26725 8618 26777
rect 18166 26725 18218 26777
rect 4294 26614 4346 26666
rect 4358 26614 4410 26666
rect 4422 26614 4474 26666
rect 4486 26614 4538 26666
rect 35014 26614 35066 26666
rect 35078 26614 35130 26666
rect 35142 26614 35194 26666
rect 35206 26614 35258 26666
rect 8230 26503 8282 26555
rect 18550 26503 18602 26555
rect 18934 26429 18986 26481
rect 8230 26318 8282 26370
rect 8518 26318 8570 26370
rect 33526 26250 33578 26259
rect 33526 26216 33535 26250
rect 33535 26216 33569 26250
rect 33569 26216 33578 26250
rect 33526 26207 33578 26216
rect 17398 26133 17450 26185
rect 17878 26059 17930 26111
rect 40438 26059 40490 26111
rect 19654 25948 19706 26000
rect 19718 25948 19770 26000
rect 19782 25948 19834 26000
rect 19846 25948 19898 26000
rect 50374 25948 50426 26000
rect 50438 25948 50490 26000
rect 50502 25948 50554 26000
rect 50566 25948 50618 26000
rect 4294 25282 4346 25334
rect 4358 25282 4410 25334
rect 4422 25282 4474 25334
rect 4486 25282 4538 25334
rect 35014 25282 35066 25334
rect 35078 25282 35130 25334
rect 35142 25282 35194 25334
rect 35206 25282 35258 25334
rect 16822 25097 16874 25149
rect 8086 24801 8138 24853
rect 11446 24801 11498 24853
rect 10774 24727 10826 24779
rect 19654 24616 19706 24668
rect 19718 24616 19770 24668
rect 19782 24616 19834 24668
rect 19846 24616 19898 24668
rect 50374 24616 50426 24668
rect 50438 24616 50490 24668
rect 50502 24616 50554 24668
rect 50566 24616 50618 24668
rect 8086 24505 8138 24557
rect 11158 24505 11210 24557
rect 18742 24209 18794 24261
rect 10966 24135 11018 24187
rect 13366 24104 13418 24113
rect 13366 24070 13375 24104
rect 13375 24070 13409 24104
rect 13409 24070 13418 24104
rect 13366 24061 13418 24070
rect 4294 23950 4346 24002
rect 4358 23950 4410 24002
rect 4422 23950 4474 24002
rect 4486 23950 4538 24002
rect 35014 23950 35066 24002
rect 35078 23950 35130 24002
rect 35142 23950 35194 24002
rect 35206 23950 35258 24002
rect 12982 23839 13034 23891
rect 13366 23839 13418 23891
rect 22678 23839 22730 23891
rect 44086 23586 44138 23595
rect 44086 23552 44095 23586
rect 44095 23552 44129 23586
rect 44129 23552 44138 23586
rect 44086 23543 44138 23552
rect 8086 23469 8138 23521
rect 16054 23395 16106 23447
rect 19654 23284 19706 23336
rect 19718 23284 19770 23336
rect 19782 23284 19834 23336
rect 19846 23284 19898 23336
rect 50374 23284 50426 23336
rect 50438 23284 50490 23336
rect 50502 23284 50554 23336
rect 50566 23284 50618 23336
rect 8086 23173 8138 23225
rect 14134 23173 14186 23225
rect 7894 22729 7946 22781
rect 44950 22729 45002 22781
rect 4294 22618 4346 22670
rect 4358 22618 4410 22670
rect 4422 22618 4474 22670
rect 4486 22618 4538 22670
rect 35014 22618 35066 22670
rect 35078 22618 35130 22670
rect 35142 22618 35194 22670
rect 35206 22618 35258 22670
rect 15478 22433 15530 22485
rect 2614 22254 2666 22263
rect 2614 22220 2623 22254
rect 2623 22220 2657 22254
rect 2657 22220 2666 22254
rect 2614 22211 2666 22220
rect 8086 22137 8138 22189
rect 13174 22137 13226 22189
rect 13462 22063 13514 22115
rect 19654 21952 19706 22004
rect 19718 21952 19770 22004
rect 19782 21952 19834 22004
rect 19846 21952 19898 22004
rect 50374 21952 50426 22004
rect 50438 21952 50490 22004
rect 50502 21952 50554 22004
rect 50566 21952 50618 22004
rect 8086 21841 8138 21893
rect 13270 21841 13322 21893
rect 32566 21841 32618 21893
rect 2614 21693 2666 21745
rect 36502 21693 36554 21745
rect 8086 21471 8138 21523
rect 55414 21471 55466 21523
rect 32278 21440 32330 21449
rect 32278 21406 32287 21440
rect 32287 21406 32321 21440
rect 32321 21406 32330 21440
rect 32278 21397 32330 21406
rect 43030 21397 43082 21449
rect 4294 21286 4346 21338
rect 4358 21286 4410 21338
rect 4422 21286 4474 21338
rect 4486 21286 4538 21338
rect 35014 21286 35066 21338
rect 35078 21286 35130 21338
rect 35142 21286 35194 21338
rect 35206 21286 35258 21338
rect 32278 21175 32330 21227
rect 44758 21175 44810 21227
rect 26422 21027 26474 21079
rect 30934 20953 30986 21005
rect 7126 20922 7178 20931
rect 7126 20888 7135 20922
rect 7135 20888 7169 20922
rect 7169 20888 7178 20922
rect 7126 20879 7178 20888
rect 29206 20879 29258 20931
rect 44854 20879 44906 20931
rect 53398 20879 53450 20931
rect 8086 20805 8138 20857
rect 16534 20805 16586 20857
rect 57718 20731 57770 20783
rect 19654 20620 19706 20672
rect 19718 20620 19770 20672
rect 19782 20620 19834 20672
rect 19846 20620 19898 20672
rect 50374 20620 50426 20672
rect 50438 20620 50490 20672
rect 50502 20620 50554 20672
rect 50566 20620 50618 20672
rect 3382 20509 3434 20561
rect 9622 20509 9674 20561
rect 12694 20509 12746 20561
rect 7126 20361 7178 20413
rect 16246 20361 16298 20413
rect 44854 20404 44906 20413
rect 44854 20370 44863 20404
rect 44863 20370 44897 20404
rect 44897 20370 44906 20404
rect 44854 20361 44906 20370
rect 9622 20330 9674 20339
rect 9622 20296 9631 20330
rect 9631 20296 9665 20330
rect 9665 20296 9674 20330
rect 9622 20287 9674 20296
rect 10582 20108 10634 20117
rect 10582 20074 10591 20108
rect 10591 20074 10625 20108
rect 10625 20074 10634 20108
rect 10582 20065 10634 20074
rect 13654 20065 13706 20117
rect 42742 20108 42794 20117
rect 42742 20074 42751 20108
rect 42751 20074 42785 20108
rect 42785 20074 42794 20108
rect 42742 20065 42794 20074
rect 43798 20065 43850 20117
rect 4294 19954 4346 20006
rect 4358 19954 4410 20006
rect 4422 19954 4474 20006
rect 4486 19954 4538 20006
rect 35014 19954 35066 20006
rect 35078 19954 35130 20006
rect 35142 19954 35194 20006
rect 35206 19954 35258 20006
rect 52822 19843 52874 19895
rect 10582 19769 10634 19821
rect 30646 19769 30698 19821
rect 55510 19621 55562 19673
rect 45910 19590 45962 19599
rect 45910 19556 45919 19590
rect 45919 19556 45953 19590
rect 45953 19556 45962 19590
rect 45910 19547 45962 19556
rect 52054 19547 52106 19599
rect 54742 19590 54794 19599
rect 54742 19556 54751 19590
rect 54751 19556 54785 19590
rect 54785 19556 54794 19590
rect 54742 19547 54794 19556
rect 50806 19473 50858 19525
rect 8758 19399 8810 19451
rect 9334 19399 9386 19451
rect 48694 19399 48746 19451
rect 19654 19288 19706 19340
rect 19718 19288 19770 19340
rect 19782 19288 19834 19340
rect 19846 19288 19898 19340
rect 50374 19288 50426 19340
rect 50438 19288 50490 19340
rect 50502 19288 50554 19340
rect 50566 19288 50618 19340
rect 8758 19177 8810 19229
rect 9334 19177 9386 19229
rect 42838 19177 42890 19229
rect 54742 19177 54794 19229
rect 36214 19103 36266 19155
rect 45910 19103 45962 19155
rect 21046 18881 21098 18933
rect 21910 18807 21962 18859
rect 25462 18733 25514 18785
rect 36118 18733 36170 18785
rect 39958 18776 40010 18785
rect 39958 18742 39967 18776
rect 39967 18742 40001 18776
rect 40001 18742 40010 18776
rect 39958 18733 40010 18742
rect 4294 18622 4346 18674
rect 4358 18622 4410 18674
rect 4422 18622 4474 18674
rect 4486 18622 4538 18674
rect 35014 18622 35066 18674
rect 35078 18622 35130 18674
rect 35142 18622 35194 18674
rect 35206 18622 35258 18674
rect 48886 18511 48938 18563
rect 46102 18363 46154 18415
rect 40342 18215 40394 18267
rect 19990 18141 20042 18193
rect 34294 18141 34346 18193
rect 14038 18067 14090 18119
rect 19654 17956 19706 18008
rect 19718 17956 19770 18008
rect 19782 17956 19834 18008
rect 19846 17956 19898 18008
rect 50374 17956 50426 18008
rect 50438 17956 50490 18008
rect 50502 17956 50554 18008
rect 50566 17956 50618 18008
rect 32470 17549 32522 17601
rect 6070 17401 6122 17453
rect 18454 17401 18506 17453
rect 4294 17290 4346 17342
rect 4358 17290 4410 17342
rect 4422 17290 4474 17342
rect 4486 17290 4538 17342
rect 35014 17290 35066 17342
rect 35078 17290 35130 17342
rect 35142 17290 35194 17342
rect 35206 17290 35258 17342
rect 42934 17179 42986 17231
rect 45238 16735 45290 16787
rect 19654 16624 19706 16676
rect 19718 16624 19770 16676
rect 19782 16624 19834 16676
rect 19846 16624 19898 16676
rect 50374 16624 50426 16676
rect 50438 16624 50490 16676
rect 50502 16624 50554 16676
rect 50566 16624 50618 16676
rect 3766 16513 3818 16565
rect 1750 16217 1802 16269
rect 3862 16143 3914 16195
rect 14710 16143 14762 16195
rect 26806 16143 26858 16195
rect 49366 16143 49418 16195
rect 16150 16069 16202 16121
rect 50038 16069 50090 16121
rect 4294 15958 4346 16010
rect 4358 15958 4410 16010
rect 4422 15958 4474 16010
rect 4486 15958 4538 16010
rect 35014 15958 35066 16010
rect 35078 15958 35130 16010
rect 35142 15958 35194 16010
rect 35206 15958 35258 16010
rect 3862 15890 3914 15899
rect 3862 15856 3871 15890
rect 3871 15856 3905 15890
rect 3905 15856 3914 15890
rect 3862 15847 3914 15856
rect 12982 15847 13034 15899
rect 16150 15890 16202 15899
rect 16150 15856 16159 15890
rect 16159 15856 16193 15890
rect 16193 15856 16202 15890
rect 16150 15847 16202 15856
rect 26806 15890 26858 15899
rect 26806 15856 26815 15890
rect 26815 15856 26849 15890
rect 26849 15856 26858 15890
rect 26806 15847 26858 15856
rect 48982 15847 49034 15899
rect 39766 15477 39818 15529
rect 42358 15403 42410 15455
rect 19654 15292 19706 15344
rect 19718 15292 19770 15344
rect 19782 15292 19834 15344
rect 19846 15292 19898 15344
rect 50374 15292 50426 15344
rect 50438 15292 50490 15344
rect 50502 15292 50554 15344
rect 50566 15292 50618 15344
rect 9622 14885 9674 14937
rect 34870 14885 34922 14937
rect 27670 14811 27722 14863
rect 27958 14737 28010 14789
rect 4294 14626 4346 14678
rect 4358 14626 4410 14678
rect 4422 14626 4474 14678
rect 4486 14626 4538 14678
rect 35014 14626 35066 14678
rect 35078 14626 35130 14678
rect 35142 14626 35194 14678
rect 35206 14626 35258 14678
rect 9622 14558 9674 14567
rect 9622 14524 9631 14558
rect 9631 14524 9665 14558
rect 9665 14524 9674 14558
rect 9622 14515 9674 14524
rect 41494 14515 41546 14567
rect 15094 14441 15146 14493
rect 53398 14441 53450 14493
rect 18262 14219 18314 14271
rect 36694 14293 36746 14345
rect 38902 14071 38954 14123
rect 19654 13960 19706 14012
rect 19718 13960 19770 14012
rect 19782 13960 19834 14012
rect 19846 13960 19898 14012
rect 50374 13960 50426 14012
rect 50438 13960 50490 14012
rect 50502 13960 50554 14012
rect 50566 13960 50618 14012
rect 21814 13849 21866 13901
rect 53590 13479 53642 13531
rect 33238 13405 33290 13457
rect 4294 13294 4346 13346
rect 4358 13294 4410 13346
rect 4422 13294 4474 13346
rect 4486 13294 4538 13346
rect 35014 13294 35066 13346
rect 35078 13294 35130 13346
rect 35142 13294 35194 13346
rect 35206 13294 35258 13346
rect 56662 13226 56714 13235
rect 56662 13192 56671 13226
rect 56671 13192 56705 13226
rect 56705 13192 56714 13226
rect 56662 13183 56714 13192
rect 36598 13109 36650 13161
rect 34102 12813 34154 12865
rect 19654 12628 19706 12680
rect 19718 12628 19770 12680
rect 19782 12628 19834 12680
rect 19846 12628 19898 12680
rect 50374 12628 50426 12680
rect 50438 12628 50490 12680
rect 50502 12628 50554 12680
rect 50566 12628 50618 12680
rect 57334 12560 57386 12569
rect 57334 12526 57343 12560
rect 57343 12526 57377 12560
rect 57377 12526 57386 12560
rect 57334 12517 57386 12526
rect 16054 12443 16106 12495
rect 15958 12221 16010 12273
rect 57526 12221 57578 12273
rect 7798 12147 7850 12199
rect 10870 12147 10922 12199
rect 9526 12073 9578 12125
rect 28822 12073 28874 12125
rect 38518 12073 38570 12125
rect 4294 11962 4346 12014
rect 4358 11962 4410 12014
rect 4422 11962 4474 12014
rect 4486 11962 4538 12014
rect 35014 11962 35066 12014
rect 35078 11962 35130 12014
rect 35142 11962 35194 12014
rect 35206 11962 35258 12014
rect 2326 11777 2378 11829
rect 7798 11777 7850 11829
rect 10486 11777 10538 11829
rect 10870 11820 10922 11829
rect 10870 11786 10879 11820
rect 10879 11786 10913 11820
rect 10913 11786 10922 11820
rect 10870 11777 10922 11786
rect 9526 11703 9578 11755
rect 32854 11777 32906 11829
rect 35830 11777 35882 11829
rect 10630 11629 10682 11681
rect 31318 11703 31370 11755
rect 59734 11777 59786 11829
rect 57142 11703 57194 11755
rect 44086 11629 44138 11681
rect 44182 11629 44234 11681
rect 44278 11598 44330 11607
rect 44278 11564 44287 11598
rect 44287 11564 44321 11598
rect 44321 11564 44330 11598
rect 44278 11555 44330 11564
rect 9526 11407 9578 11459
rect 19654 11296 19706 11348
rect 19718 11296 19770 11348
rect 19782 11296 19834 11348
rect 19846 11296 19898 11348
rect 50374 11296 50426 11348
rect 50438 11296 50490 11348
rect 50502 11296 50554 11348
rect 50566 11296 50618 11348
rect 5206 11228 5258 11237
rect 5206 11194 5215 11228
rect 5215 11194 5249 11228
rect 5249 11194 5258 11228
rect 5206 11185 5258 11194
rect 9526 11185 9578 11237
rect 27190 11185 27242 11237
rect 56950 11228 57002 11237
rect 56950 11194 56959 11228
rect 56959 11194 56993 11228
rect 56993 11194 57002 11228
rect 56950 11185 57002 11194
rect 8086 10963 8138 11015
rect 24022 10963 24074 11015
rect 8278 10815 8330 10867
rect 15766 10815 15818 10867
rect 56374 10889 56426 10941
rect 56758 10889 56810 10941
rect 6742 10741 6794 10793
rect 10678 10741 10730 10793
rect 15094 10741 15146 10793
rect 54454 10815 54506 10867
rect 4294 10630 4346 10682
rect 4358 10630 4410 10682
rect 4422 10630 4474 10682
rect 4486 10630 4538 10682
rect 35014 10630 35066 10682
rect 35078 10630 35130 10682
rect 35142 10630 35194 10682
rect 35206 10630 35258 10682
rect 10198 10519 10250 10571
rect 10678 10519 10730 10571
rect 56086 10562 56138 10571
rect 25654 10371 25706 10423
rect 8086 10297 8138 10349
rect 24694 10297 24746 10349
rect 38806 10266 38858 10275
rect 38806 10232 38815 10266
rect 38815 10232 38849 10266
rect 38849 10232 38858 10266
rect 38806 10223 38858 10232
rect 56086 10528 56095 10562
rect 56095 10528 56129 10562
rect 56129 10528 56138 10562
rect 56086 10519 56138 10528
rect 56470 10371 56522 10423
rect 29782 10149 29834 10201
rect 26518 10075 26570 10127
rect 58582 10149 58634 10201
rect 55702 10075 55754 10127
rect 56086 10075 56138 10127
rect 19654 9964 19706 10016
rect 19718 9964 19770 10016
rect 19782 9964 19834 10016
rect 19846 9964 19898 10016
rect 50374 9964 50426 10016
rect 50438 9964 50490 10016
rect 50502 9964 50554 10016
rect 50566 9964 50618 10016
rect 8182 9853 8234 9905
rect 23446 9853 23498 9905
rect 54646 9896 54698 9905
rect 8374 9705 8426 9757
rect 20854 9705 20906 9757
rect 54646 9862 54655 9896
rect 54655 9862 54689 9896
rect 54689 9862 54698 9896
rect 54646 9853 54698 9862
rect 55606 9896 55658 9905
rect 55606 9862 55615 9896
rect 55615 9862 55649 9896
rect 55649 9862 55658 9896
rect 55606 9853 55658 9862
rect 8086 9631 8138 9683
rect 19318 9631 19370 9683
rect 57622 9674 57674 9683
rect 57622 9640 57631 9674
rect 57631 9640 57665 9674
rect 57665 9640 57674 9674
rect 57622 9631 57674 9640
rect 8662 9557 8714 9609
rect 13366 9557 13418 9609
rect 17302 9557 17354 9609
rect 36790 9557 36842 9609
rect 54262 9557 54314 9609
rect 11542 9483 11594 9535
rect 24310 9483 24362 9535
rect 50710 9483 50762 9535
rect 10678 9409 10730 9461
rect 17974 9409 18026 9461
rect 25366 9409 25418 9461
rect 37270 9409 37322 9461
rect 48214 9409 48266 9461
rect 54934 9483 54986 9535
rect 55510 9557 55562 9609
rect 4294 9298 4346 9350
rect 4358 9298 4410 9350
rect 4422 9298 4474 9350
rect 4486 9298 4538 9350
rect 35014 9298 35066 9350
rect 35078 9298 35130 9350
rect 35142 9298 35194 9350
rect 35206 9298 35258 9350
rect 8182 9113 8234 9165
rect 8086 9039 8138 9091
rect 8374 9039 8426 9091
rect 10678 9187 10730 9239
rect 12022 9230 12074 9239
rect 12022 9196 12031 9230
rect 12031 9196 12065 9230
rect 12065 9196 12074 9230
rect 12022 9187 12074 9196
rect 48214 9113 48266 9165
rect 16342 9039 16394 9091
rect 22966 9039 23018 9091
rect 53398 9082 53450 9091
rect 53398 9048 53407 9082
rect 53407 9048 53441 9082
rect 53441 9048 53450 9082
rect 53398 9039 53450 9048
rect 12982 8965 13034 9017
rect 56854 8965 56906 9017
rect 57238 9008 57290 9017
rect 57238 8974 57247 9008
rect 57247 8974 57281 9008
rect 57281 8974 57290 9008
rect 57238 8965 57290 8974
rect 13750 8891 13802 8943
rect 46294 8934 46346 8943
rect 16726 8817 16778 8869
rect 18070 8817 18122 8869
rect 8086 8743 8138 8795
rect 16822 8743 16874 8795
rect 17686 8743 17738 8795
rect 46294 8900 46303 8934
rect 46303 8900 46337 8934
rect 46337 8900 46346 8934
rect 46294 8891 46346 8900
rect 49750 8817 49802 8869
rect 50230 8817 50282 8869
rect 55990 8891 56042 8943
rect 54550 8817 54602 8869
rect 53878 8743 53930 8795
rect 19654 8632 19706 8684
rect 19718 8632 19770 8684
rect 19782 8632 19834 8684
rect 19846 8632 19898 8684
rect 50374 8632 50426 8684
rect 50438 8632 50490 8684
rect 50502 8632 50554 8684
rect 50566 8632 50618 8684
rect 9910 8521 9962 8573
rect 1750 8416 1802 8425
rect 1750 8382 1759 8416
rect 1759 8382 1793 8416
rect 1793 8382 1802 8416
rect 1750 8373 1802 8382
rect 2422 8416 2474 8425
rect 2422 8382 2431 8416
rect 2431 8382 2465 8416
rect 2465 8382 2474 8416
rect 2422 8373 2474 8382
rect 3286 8416 3338 8425
rect 3286 8382 3295 8416
rect 3295 8382 3329 8416
rect 3329 8382 3338 8416
rect 3286 8373 3338 8382
rect 11734 8447 11786 8499
rect 7798 8373 7850 8425
rect 10294 8373 10346 8425
rect 11350 8416 11402 8425
rect 11350 8382 11359 8416
rect 11359 8382 11393 8416
rect 11393 8382 11402 8416
rect 11350 8373 11402 8382
rect 12214 8521 12266 8573
rect 16054 8521 16106 8573
rect 11926 8447 11978 8499
rect 34678 8521 34730 8573
rect 48598 8564 48650 8573
rect 48598 8530 48607 8564
rect 48607 8530 48641 8564
rect 48641 8530 48650 8564
rect 48598 8521 48650 8530
rect 50134 8521 50186 8573
rect 52918 8564 52970 8573
rect 13654 8416 13706 8425
rect 13654 8382 13663 8416
rect 13663 8382 13697 8416
rect 13697 8382 13706 8416
rect 13654 8373 13706 8382
rect 16054 8373 16106 8425
rect 7606 8299 7658 8351
rect 8278 8299 8330 8351
rect 20086 8373 20138 8425
rect 25654 8416 25706 8425
rect 25654 8382 25663 8416
rect 25663 8382 25697 8416
rect 25697 8382 25706 8416
rect 25654 8373 25706 8382
rect 16822 8299 16874 8351
rect 1654 8268 1706 8277
rect 1654 8234 1663 8268
rect 1663 8234 1697 8268
rect 1697 8234 1706 8268
rect 1654 8225 1706 8234
rect 2230 8151 2282 8203
rect 3286 8225 3338 8277
rect 7702 8225 7754 8277
rect 9526 8225 9578 8277
rect 10582 8268 10634 8277
rect 10582 8234 10591 8268
rect 10591 8234 10625 8268
rect 10625 8234 10634 8268
rect 10582 8225 10634 8234
rect 10678 8225 10730 8277
rect 11350 8225 11402 8277
rect 12310 8225 12362 8277
rect 12886 8225 12938 8277
rect 16054 8225 16106 8277
rect 16342 8225 16394 8277
rect 23542 8299 23594 8351
rect 52918 8530 52927 8564
rect 52927 8530 52961 8564
rect 52961 8530 52970 8564
rect 52918 8521 52970 8530
rect 49846 8299 49898 8351
rect 4822 8151 4874 8203
rect 13750 8151 13802 8203
rect 8086 8077 8138 8129
rect 9814 8077 9866 8129
rect 10582 8077 10634 8129
rect 48022 8225 48074 8277
rect 48886 8225 48938 8277
rect 17110 8151 17162 8203
rect 28054 8077 28106 8129
rect 33526 8077 33578 8129
rect 44374 8077 44426 8129
rect 48694 8151 48746 8203
rect 49462 8225 49514 8277
rect 52150 8151 52202 8203
rect 53110 8225 53162 8277
rect 53494 8225 53546 8277
rect 56950 8299 57002 8351
rect 58390 8225 58442 8277
rect 50806 8077 50858 8129
rect 59830 8151 59882 8203
rect 58966 8077 59018 8129
rect 4294 7966 4346 8018
rect 4358 7966 4410 8018
rect 4422 7966 4474 8018
rect 4486 7966 4538 8018
rect 35014 7966 35066 8018
rect 35078 7966 35130 8018
rect 35142 7966 35194 8018
rect 35206 7966 35258 8018
rect 2134 7898 2186 7907
rect 2134 7864 2143 7898
rect 2143 7864 2177 7898
rect 2177 7864 2186 7898
rect 2134 7855 2186 7864
rect 3670 7898 3722 7907
rect 3670 7864 3679 7898
rect 3679 7864 3713 7898
rect 3713 7864 3722 7898
rect 7606 7898 7658 7907
rect 3670 7855 3722 7864
rect 7606 7864 7615 7898
rect 7615 7864 7649 7898
rect 7649 7864 7658 7898
rect 7606 7855 7658 7864
rect 9046 7898 9098 7907
rect 5686 7707 5738 7759
rect 1462 7633 1514 7685
rect 9046 7864 9055 7898
rect 9055 7864 9089 7898
rect 9089 7864 9098 7898
rect 9046 7855 9098 7864
rect 28054 7855 28106 7907
rect 29014 7898 29066 7907
rect 29014 7864 29023 7898
rect 29023 7864 29057 7898
rect 29057 7864 29066 7898
rect 36502 7898 36554 7907
rect 29014 7855 29066 7864
rect 9622 7781 9674 7833
rect 8086 7707 8138 7759
rect 8374 7707 8426 7759
rect 9046 7707 9098 7759
rect 9142 7633 9194 7685
rect 10198 7676 10250 7685
rect 10198 7642 10207 7676
rect 10207 7642 10241 7676
rect 10241 7642 10250 7676
rect 10198 7633 10250 7642
rect 13750 7781 13802 7833
rect 25078 7824 25130 7833
rect 12598 7707 12650 7759
rect 12694 7707 12746 7759
rect 25078 7790 25087 7824
rect 25087 7790 25121 7824
rect 25121 7790 25130 7824
rect 25078 7781 25130 7790
rect 15862 7750 15914 7759
rect 15862 7716 15871 7750
rect 15871 7716 15905 7750
rect 15905 7716 15914 7750
rect 15862 7707 15914 7716
rect 20950 7750 21002 7759
rect 20950 7716 20959 7750
rect 20959 7716 20993 7750
rect 20993 7716 21002 7750
rect 20950 7707 21002 7716
rect 23926 7750 23978 7759
rect 23926 7716 23935 7750
rect 23935 7716 23969 7750
rect 23969 7716 23978 7750
rect 23926 7707 23978 7716
rect 24694 7750 24746 7759
rect 24694 7716 24703 7750
rect 24703 7716 24737 7750
rect 24737 7716 24746 7750
rect 24694 7707 24746 7716
rect 27766 7781 27818 7833
rect 26134 7750 26186 7759
rect 26134 7716 26143 7750
rect 26143 7716 26177 7750
rect 26177 7716 26186 7750
rect 26134 7707 26186 7716
rect 26998 7750 27050 7759
rect 26998 7716 27007 7750
rect 27007 7716 27041 7750
rect 27041 7716 27050 7750
rect 26998 7707 27050 7716
rect 36502 7864 36511 7898
rect 36511 7864 36545 7898
rect 36545 7864 36554 7898
rect 41494 7898 41546 7907
rect 36502 7855 36554 7864
rect 30166 7750 30218 7759
rect 30166 7716 30175 7750
rect 30175 7716 30209 7750
rect 30209 7716 30218 7750
rect 30166 7707 30218 7716
rect 12310 7633 12362 7685
rect 5590 7602 5642 7611
rect 5590 7568 5599 7602
rect 5599 7568 5633 7602
rect 5633 7568 5642 7602
rect 5590 7559 5642 7568
rect 11254 7559 11306 7611
rect 12502 7559 12554 7611
rect 17110 7559 17162 7611
rect 33334 7707 33386 7759
rect 33814 7707 33866 7759
rect 34582 7750 34634 7759
rect 34582 7716 34591 7750
rect 34591 7716 34625 7750
rect 34625 7716 34634 7750
rect 34582 7707 34634 7716
rect 35350 7750 35402 7759
rect 35350 7716 35359 7750
rect 35359 7716 35393 7750
rect 35393 7716 35402 7750
rect 35350 7707 35402 7716
rect 36118 7750 36170 7759
rect 36118 7716 36127 7750
rect 36127 7716 36161 7750
rect 36161 7716 36170 7750
rect 36118 7707 36170 7716
rect 41494 7864 41503 7898
rect 41503 7864 41537 7898
rect 41537 7864 41546 7898
rect 41494 7855 41546 7864
rect 42262 7898 42314 7907
rect 42262 7864 42271 7898
rect 42271 7864 42305 7898
rect 42305 7864 42314 7898
rect 42262 7855 42314 7864
rect 38806 7781 38858 7833
rect 38710 7750 38762 7759
rect 38710 7716 38719 7750
rect 38719 7716 38753 7750
rect 38753 7716 38762 7750
rect 38710 7707 38762 7716
rect 39478 7750 39530 7759
rect 39478 7716 39487 7750
rect 39487 7716 39521 7750
rect 39521 7716 39530 7750
rect 39478 7707 39530 7716
rect 38806 7633 38858 7685
rect 34486 7559 34538 7611
rect 40342 7750 40394 7759
rect 40342 7716 40351 7750
rect 40351 7716 40385 7750
rect 40385 7716 40394 7750
rect 40342 7707 40394 7716
rect 40246 7633 40298 7685
rect 41398 7707 41450 7759
rect 45046 7855 45098 7907
rect 47542 7898 47594 7907
rect 44758 7707 44810 7759
rect 47542 7864 47551 7898
rect 47551 7864 47585 7898
rect 47585 7864 47594 7898
rect 47542 7855 47594 7864
rect 46294 7707 46346 7759
rect 49558 7855 49610 7907
rect 49366 7750 49418 7759
rect 49366 7716 49375 7750
rect 49375 7716 49409 7750
rect 49409 7716 49418 7750
rect 49366 7707 49418 7716
rect 50038 7707 50090 7759
rect 59350 7781 59402 7833
rect 53590 7707 53642 7759
rect 44278 7633 44330 7685
rect 45430 7633 45482 7685
rect 49750 7633 49802 7685
rect 55798 7676 55850 7685
rect 39958 7559 40010 7611
rect 41494 7559 41546 7611
rect 45334 7559 45386 7611
rect 52822 7559 52874 7611
rect 55798 7642 55807 7676
rect 55807 7642 55841 7676
rect 55841 7642 55850 7676
rect 55798 7633 55850 7642
rect 56182 7633 56234 7685
rect 56662 7633 56714 7685
rect 58774 7559 58826 7611
rect 39478 7485 39530 7537
rect 2326 7411 2378 7463
rect 2998 7411 3050 7463
rect 3958 7454 4010 7463
rect 3958 7420 3967 7454
rect 3967 7420 4001 7454
rect 4001 7420 4010 7454
rect 3958 7411 4010 7420
rect 4054 7411 4106 7463
rect 5302 7411 5354 7463
rect 8374 7411 8426 7463
rect 8758 7411 8810 7463
rect 9910 7411 9962 7463
rect 10966 7411 11018 7463
rect 12406 7411 12458 7463
rect 15670 7411 15722 7463
rect 20758 7411 20810 7463
rect 23830 7454 23882 7463
rect 23830 7420 23839 7454
rect 23839 7420 23873 7454
rect 23873 7420 23882 7454
rect 23830 7411 23882 7420
rect 24214 7411 24266 7463
rect 24790 7411 24842 7463
rect 25558 7411 25610 7463
rect 26710 7411 26762 7463
rect 28150 7411 28202 7463
rect 29206 7411 29258 7463
rect 29590 7411 29642 7463
rect 31126 7454 31178 7463
rect 31126 7420 31135 7454
rect 31135 7420 31169 7454
rect 31169 7420 31178 7454
rect 31126 7411 31178 7420
rect 33622 7411 33674 7463
rect 34390 7411 34442 7463
rect 34678 7411 34730 7463
rect 36022 7454 36074 7463
rect 36022 7420 36031 7454
rect 36031 7420 36065 7454
rect 36065 7420 36074 7454
rect 36022 7411 36074 7420
rect 36598 7411 36650 7463
rect 38038 7411 38090 7463
rect 42454 7411 42506 7463
rect 43894 7411 43946 7463
rect 44662 7411 44714 7463
rect 45046 7411 45098 7463
rect 45814 7411 45866 7463
rect 46582 7411 46634 7463
rect 47254 7411 47306 7463
rect 48310 7411 48362 7463
rect 50038 7454 50090 7463
rect 50038 7420 50047 7454
rect 50047 7420 50081 7454
rect 50081 7420 50090 7454
rect 50038 7411 50090 7420
rect 51670 7411 51722 7463
rect 52342 7411 52394 7463
rect 52726 7411 52778 7463
rect 19654 7300 19706 7352
rect 19718 7300 19770 7352
rect 19782 7300 19834 7352
rect 19846 7300 19898 7352
rect 50374 7300 50426 7352
rect 50438 7300 50490 7352
rect 50502 7300 50554 7352
rect 50566 7300 50618 7352
rect 5590 7189 5642 7241
rect 12502 7189 12554 7241
rect 12790 7189 12842 7241
rect 12982 7189 13034 7241
rect 8854 7115 8906 7167
rect 11542 7115 11594 7167
rect 6070 7084 6122 7093
rect 6070 7050 6079 7084
rect 6079 7050 6113 7084
rect 6113 7050 6122 7084
rect 6070 7041 6122 7050
rect 17110 7189 17162 7241
rect 17974 7232 18026 7241
rect 17974 7198 17983 7232
rect 17983 7198 18017 7232
rect 18017 7198 18026 7232
rect 17974 7189 18026 7198
rect 18646 7189 18698 7241
rect 17302 7115 17354 7167
rect 1654 7010 1706 7019
rect 1654 6976 1663 7010
rect 1663 6976 1697 7010
rect 1697 6976 1706 7010
rect 1654 6967 1706 6976
rect 2518 7010 2570 7019
rect 2518 6976 2527 7010
rect 2527 6976 2561 7010
rect 2561 6976 2570 7010
rect 2518 6967 2570 6976
rect 11254 7010 11306 7019
rect 5110 6893 5162 6945
rect 5014 6819 5066 6871
rect 3670 6745 3722 6797
rect 5878 6893 5930 6945
rect 6550 6893 6602 6945
rect 6934 6893 6986 6945
rect 7798 6893 7850 6945
rect 9718 6936 9770 6945
rect 7318 6819 7370 6871
rect 9718 6902 9727 6936
rect 9727 6902 9761 6936
rect 9761 6902 9770 6936
rect 9718 6893 9770 6902
rect 9814 6936 9866 6945
rect 9814 6902 9823 6936
rect 9823 6902 9857 6936
rect 9857 6902 9866 6936
rect 9814 6893 9866 6902
rect 11254 6976 11263 7010
rect 11263 6976 11297 7010
rect 11297 6976 11306 7010
rect 11254 6967 11306 6976
rect 12694 7010 12746 7019
rect 12694 6976 12703 7010
rect 12703 6976 12737 7010
rect 12737 6976 12746 7010
rect 12694 6967 12746 6976
rect 15094 7084 15146 7093
rect 15094 7050 15103 7084
rect 15103 7050 15137 7084
rect 15137 7050 15146 7084
rect 15094 7041 15146 7050
rect 15958 7041 16010 7093
rect 18070 7084 18122 7093
rect 18070 7050 18079 7084
rect 18079 7050 18113 7084
rect 18113 7050 18122 7084
rect 18070 7041 18122 7050
rect 18934 7041 18986 7093
rect 20374 7084 20426 7093
rect 20374 7050 20383 7084
rect 20383 7050 20417 7084
rect 20417 7050 20426 7084
rect 20374 7041 20426 7050
rect 21142 7084 21194 7093
rect 21142 7050 21151 7084
rect 21151 7050 21185 7084
rect 21185 7050 21194 7084
rect 21142 7041 21194 7050
rect 21910 7084 21962 7093
rect 21910 7050 21919 7084
rect 21919 7050 21953 7084
rect 21953 7050 21962 7084
rect 21910 7041 21962 7050
rect 22678 7084 22730 7093
rect 22678 7050 22687 7084
rect 22687 7050 22721 7084
rect 22721 7050 22730 7084
rect 22678 7041 22730 7050
rect 23062 7158 23114 7167
rect 23062 7124 23071 7158
rect 23071 7124 23105 7158
rect 23105 7124 23114 7158
rect 28342 7158 28394 7167
rect 23062 7115 23114 7124
rect 23350 7041 23402 7093
rect 24310 7041 24362 7093
rect 16630 7010 16682 7019
rect 16630 6976 16639 7010
rect 16639 6976 16673 7010
rect 16673 6976 16682 7010
rect 16630 6967 16682 6976
rect 28342 7124 28351 7158
rect 28351 7124 28385 7158
rect 28385 7124 28394 7158
rect 28342 7115 28394 7124
rect 25462 7041 25514 7093
rect 26326 7084 26378 7093
rect 26326 7050 26335 7084
rect 26335 7050 26369 7084
rect 26369 7050 26378 7084
rect 26326 7041 26378 7050
rect 27286 7041 27338 7093
rect 27958 7084 28010 7093
rect 27958 7050 27967 7084
rect 27967 7050 28001 7084
rect 28001 7050 28010 7084
rect 27958 7041 28010 7050
rect 29014 7115 29066 7167
rect 32182 7115 32234 7167
rect 33718 7158 33770 7167
rect 33718 7124 33727 7158
rect 33727 7124 33761 7158
rect 33761 7124 33770 7158
rect 33718 7115 33770 7124
rect 37654 7115 37706 7167
rect 41110 7158 41162 7167
rect 41110 7124 41119 7158
rect 41119 7124 41153 7158
rect 41153 7124 41162 7158
rect 41110 7115 41162 7124
rect 31030 7041 31082 7093
rect 31702 7084 31754 7093
rect 31702 7050 31711 7084
rect 31711 7050 31745 7084
rect 31745 7050 31754 7084
rect 31702 7041 31754 7050
rect 32662 7041 32714 7093
rect 33238 7084 33290 7093
rect 33238 7050 33247 7084
rect 33247 7050 33281 7084
rect 33281 7050 33290 7084
rect 33238 7041 33290 7050
rect 34774 7084 34826 7093
rect 34774 7050 34783 7084
rect 34783 7050 34817 7084
rect 34817 7050 34826 7084
rect 34774 7041 34826 7050
rect 36214 7084 36266 7093
rect 36214 7050 36223 7084
rect 36223 7050 36257 7084
rect 36257 7050 36266 7084
rect 36214 7041 36266 7050
rect 37750 7084 37802 7093
rect 37750 7050 37759 7084
rect 37759 7050 37793 7084
rect 37793 7050 37802 7084
rect 37750 7041 37802 7050
rect 38518 7084 38570 7093
rect 38518 7050 38527 7084
rect 38527 7050 38561 7084
rect 38561 7050 38570 7084
rect 38518 7041 38570 7050
rect 41494 7115 41546 7167
rect 43606 7115 43658 7167
rect 48790 7158 48842 7167
rect 48790 7124 48799 7158
rect 48799 7124 48833 7158
rect 48833 7124 48842 7158
rect 48790 7115 48842 7124
rect 43030 7084 43082 7093
rect 43030 7050 43039 7084
rect 43039 7050 43073 7084
rect 43073 7050 43082 7084
rect 43030 7041 43082 7050
rect 43798 7084 43850 7093
rect 43798 7050 43807 7084
rect 43807 7050 43841 7084
rect 43841 7050 43850 7084
rect 43798 7041 43850 7050
rect 44278 7041 44330 7093
rect 10582 6936 10634 6945
rect 10582 6902 10591 6936
rect 10591 6902 10625 6936
rect 10625 6902 10634 6936
rect 10582 6893 10634 6902
rect 13462 6893 13514 6945
rect 14614 6893 14666 6945
rect 15382 6893 15434 6945
rect 25174 6967 25226 7019
rect 17302 6936 17354 6945
rect 17302 6902 17311 6936
rect 17311 6902 17345 6936
rect 17345 6902 17354 6936
rect 17302 6893 17354 6902
rect 19510 6893 19562 6945
rect 20374 6893 20426 6945
rect 21142 6893 21194 6945
rect 21910 6893 21962 6945
rect 22678 6893 22730 6945
rect 23446 6893 23498 6945
rect 24502 6893 24554 6945
rect 25942 6967 25994 7019
rect 26998 6967 27050 7019
rect 28534 6967 28586 7019
rect 27958 6893 28010 6945
rect 30742 6967 30794 7019
rect 29974 6893 30026 6945
rect 32182 6967 32234 7019
rect 31702 6893 31754 6945
rect 34486 6967 34538 7019
rect 37366 6967 37418 7019
rect 33718 6893 33770 6945
rect 34102 6893 34154 6945
rect 35542 6893 35594 6945
rect 36502 6893 36554 6945
rect 37078 6893 37130 6945
rect 38518 6893 38570 6945
rect 44374 6967 44426 7019
rect 45142 7041 45194 7093
rect 47350 7041 47402 7093
rect 49942 7158 49994 7167
rect 49942 7124 49951 7158
rect 49951 7124 49985 7158
rect 49985 7124 49994 7158
rect 49942 7115 49994 7124
rect 52054 7084 52106 7093
rect 52054 7050 52063 7084
rect 52063 7050 52097 7084
rect 52097 7050 52106 7084
rect 52054 7041 52106 7050
rect 38134 6819 38186 6871
rect 38230 6819 38282 6871
rect 36406 6745 36458 6797
rect 42262 6936 42314 6945
rect 39862 6819 39914 6871
rect 42262 6902 42271 6936
rect 42271 6902 42305 6936
rect 42305 6902 42314 6936
rect 42262 6893 42314 6902
rect 41590 6819 41642 6871
rect 43030 6893 43082 6945
rect 52534 6967 52586 7019
rect 54742 7010 54794 7019
rect 43990 6819 44042 6871
rect 45718 6819 45770 6871
rect 47062 6893 47114 6945
rect 46870 6819 46922 6871
rect 48406 6893 48458 6945
rect 50134 6819 50186 6871
rect 50422 6893 50474 6945
rect 51190 6893 51242 6945
rect 51574 6893 51626 6945
rect 50230 6745 50282 6797
rect 54742 6976 54751 7010
rect 54751 6976 54785 7010
rect 54785 6976 54794 7010
rect 54742 6967 54794 6976
rect 55414 6967 55466 7019
rect 58486 6967 58538 7019
rect 52246 6819 52298 6871
rect 57046 6893 57098 6945
rect 4294 6634 4346 6686
rect 4358 6634 4410 6686
rect 4422 6634 4474 6686
rect 4486 6634 4538 6686
rect 35014 6634 35066 6686
rect 35078 6634 35130 6686
rect 35142 6634 35194 6686
rect 35206 6634 35258 6686
rect 5398 6566 5450 6575
rect 5398 6532 5407 6566
rect 5407 6532 5441 6566
rect 5441 6532 5450 6566
rect 5398 6523 5450 6532
rect 6646 6523 6698 6575
rect 10582 6523 10634 6575
rect 13078 6523 13130 6575
rect 14038 6523 14090 6575
rect 18838 6566 18890 6575
rect 18838 6532 18847 6566
rect 18847 6532 18881 6566
rect 18881 6532 18890 6566
rect 18838 6523 18890 6532
rect 20566 6523 20618 6575
rect 22582 6566 22634 6575
rect 22582 6532 22591 6566
rect 22591 6532 22625 6566
rect 22625 6532 22634 6566
rect 22582 6523 22634 6532
rect 24118 6566 24170 6575
rect 24118 6532 24127 6566
rect 24127 6532 24161 6566
rect 24161 6532 24170 6566
rect 24118 6523 24170 6532
rect 27862 6566 27914 6575
rect 27862 6532 27871 6566
rect 27871 6532 27905 6566
rect 27905 6532 27914 6566
rect 27862 6523 27914 6532
rect 31798 6566 31850 6575
rect 31798 6532 31807 6566
rect 31807 6532 31841 6566
rect 31841 6532 31850 6566
rect 31798 6523 31850 6532
rect 42262 6523 42314 6575
rect 46486 6566 46538 6575
rect 46486 6532 46495 6566
rect 46495 6532 46529 6566
rect 46529 6532 46538 6566
rect 46486 6523 46538 6532
rect 49654 6523 49706 6575
rect 51286 6566 51338 6575
rect 9238 6449 9290 6501
rect 9814 6449 9866 6501
rect 50422 6449 50474 6501
rect 6262 6375 6314 6427
rect 7126 6375 7178 6427
rect 13942 6418 13994 6427
rect 13942 6384 13951 6418
rect 13951 6384 13985 6418
rect 13985 6384 13994 6418
rect 13942 6375 13994 6384
rect 14710 6418 14762 6427
rect 14710 6384 14719 6418
rect 14719 6384 14753 6418
rect 14753 6384 14762 6418
rect 14710 6375 14762 6384
rect 15478 6418 15530 6427
rect 15478 6384 15487 6418
rect 15487 6384 15521 6418
rect 15521 6384 15530 6418
rect 15478 6375 15530 6384
rect 16246 6418 16298 6427
rect 16246 6384 16255 6418
rect 16255 6384 16289 6418
rect 16289 6384 16298 6418
rect 16246 6375 16298 6384
rect 17686 6418 17738 6427
rect 17686 6384 17695 6418
rect 17695 6384 17729 6418
rect 17729 6384 17738 6418
rect 17686 6375 17738 6384
rect 18454 6418 18506 6427
rect 18454 6384 18463 6418
rect 18463 6384 18497 6418
rect 18497 6384 18506 6418
rect 18454 6375 18506 6384
rect 18838 6375 18890 6427
rect 20566 6375 20618 6427
rect 1558 6344 1610 6353
rect 1558 6310 1567 6344
rect 1567 6310 1601 6344
rect 1601 6310 1610 6344
rect 1558 6301 1610 6310
rect 2038 6301 2090 6353
rect 3190 6344 3242 6353
rect 3190 6310 3199 6344
rect 3199 6310 3233 6344
rect 3233 6310 3242 6344
rect 3190 6301 3242 6310
rect 3862 6301 3914 6353
rect 4630 6301 4682 6353
rect 9430 6344 9482 6353
rect 9430 6310 9439 6344
rect 9439 6310 9473 6344
rect 9473 6310 9482 6344
rect 9430 6301 9482 6310
rect 10102 6301 10154 6353
rect 10870 6301 10922 6353
rect 11638 6301 11690 6353
rect 13078 6344 13130 6353
rect 13078 6310 13087 6344
rect 13087 6310 13121 6344
rect 13121 6310 13130 6344
rect 13078 6301 13130 6310
rect 15958 6301 16010 6353
rect 20086 6301 20138 6353
rect 22582 6375 22634 6427
rect 23734 6418 23786 6427
rect 23734 6384 23743 6418
rect 23743 6384 23777 6418
rect 23777 6384 23786 6418
rect 23734 6375 23786 6384
rect 24118 6375 24170 6427
rect 27862 6375 27914 6427
rect 29110 6375 29162 6427
rect 30646 6418 30698 6427
rect 30646 6384 30655 6418
rect 30655 6384 30689 6418
rect 30689 6384 30698 6418
rect 30646 6375 30698 6384
rect 31798 6375 31850 6427
rect 34294 6418 34346 6427
rect 34294 6384 34303 6418
rect 34303 6384 34337 6418
rect 34337 6384 34346 6418
rect 34294 6375 34346 6384
rect 34870 6375 34922 6427
rect 37270 6418 37322 6427
rect 37270 6384 37279 6418
rect 37279 6384 37313 6418
rect 37313 6384 37322 6418
rect 37270 6375 37322 6384
rect 41302 6418 41354 6427
rect 41302 6384 41311 6418
rect 41311 6384 41345 6418
rect 41345 6384 41354 6418
rect 41302 6375 41354 6384
rect 42838 6418 42890 6427
rect 42838 6384 42847 6418
rect 42847 6384 42881 6418
rect 42881 6384 42890 6418
rect 42838 6375 42890 6384
rect 44086 6418 44138 6427
rect 44086 6384 44095 6418
rect 44095 6384 44129 6418
rect 44129 6384 44138 6418
rect 44086 6375 44138 6384
rect 44950 6375 45002 6427
rect 49846 6375 49898 6427
rect 25366 6301 25418 6353
rect 25654 6344 25706 6353
rect 25654 6310 25663 6344
rect 25663 6310 25697 6344
rect 25697 6310 25706 6344
rect 25654 6301 25706 6310
rect 26806 6344 26858 6353
rect 26806 6310 26815 6344
rect 26815 6310 26849 6344
rect 26849 6310 26858 6344
rect 26806 6301 26858 6310
rect 29686 6344 29738 6353
rect 29686 6310 29695 6344
rect 29695 6310 29729 6344
rect 29729 6310 29738 6344
rect 29686 6301 29738 6310
rect 31222 6344 31274 6353
rect 31222 6310 31231 6344
rect 31231 6310 31265 6344
rect 31265 6310 31274 6344
rect 31222 6301 31274 6310
rect 32566 6301 32618 6353
rect 36310 6344 36362 6353
rect 36310 6310 36319 6344
rect 36319 6310 36353 6344
rect 36353 6310 36362 6344
rect 36310 6301 36362 6310
rect 38902 6344 38954 6353
rect 38902 6310 38911 6344
rect 38911 6310 38945 6344
rect 38945 6310 38954 6344
rect 38902 6301 38954 6310
rect 40342 6344 40394 6353
rect 40342 6310 40351 6344
rect 40351 6310 40385 6344
rect 40385 6310 40394 6344
rect 40342 6301 40394 6310
rect 41878 6344 41930 6353
rect 41878 6310 41887 6344
rect 41887 6310 41921 6344
rect 41921 6310 41930 6344
rect 41878 6301 41930 6310
rect 45526 6344 45578 6353
rect 45526 6310 45535 6344
rect 45535 6310 45569 6344
rect 45569 6310 45578 6344
rect 45526 6301 45578 6310
rect 46966 6344 47018 6353
rect 46966 6310 46975 6344
rect 46975 6310 47009 6344
rect 47009 6310 47018 6344
rect 46966 6301 47018 6310
rect 47734 6344 47786 6353
rect 47734 6310 47743 6344
rect 47743 6310 47777 6344
rect 47777 6310 47786 6344
rect 47734 6301 47786 6310
rect 48790 6301 48842 6353
rect 49558 6301 49610 6353
rect 51286 6532 51295 6566
rect 51295 6532 51329 6566
rect 51329 6532 51338 6566
rect 51286 6523 51338 6532
rect 51094 6301 51146 6353
rect 7126 6270 7178 6279
rect 7126 6236 7135 6270
rect 7135 6236 7169 6270
rect 7169 6236 7178 6270
rect 7126 6227 7178 6236
rect 14902 6227 14954 6279
rect 5206 6153 5258 6205
rect 5494 6079 5546 6131
rect 14230 6153 14282 6205
rect 13750 6079 13802 6131
rect 13942 6079 13994 6131
rect 19318 6227 19370 6279
rect 18070 6153 18122 6205
rect 16726 6079 16778 6131
rect 18358 6122 18410 6131
rect 18358 6088 18367 6122
rect 18367 6088 18401 6122
rect 18401 6088 18410 6122
rect 18358 6079 18410 6088
rect 18934 6153 18986 6205
rect 22966 6227 23018 6279
rect 33526 6270 33578 6279
rect 22294 6153 22346 6205
rect 22870 6122 22922 6131
rect 22870 6088 22879 6122
rect 22879 6088 22913 6122
rect 22913 6088 22922 6122
rect 22870 6079 22922 6088
rect 33526 6236 33535 6270
rect 33535 6236 33569 6270
rect 33569 6236 33578 6270
rect 33526 6227 33578 6236
rect 38134 6227 38186 6279
rect 46678 6227 46730 6279
rect 27478 6153 27530 6205
rect 26326 6079 26378 6131
rect 31798 6153 31850 6205
rect 29782 6079 29834 6131
rect 31510 6079 31562 6131
rect 40630 6153 40682 6205
rect 33814 6079 33866 6131
rect 35350 6079 35402 6131
rect 39190 6079 39242 6131
rect 42166 6153 42218 6205
rect 52438 6227 52490 6279
rect 51478 6153 51530 6205
rect 53974 6301 54026 6353
rect 54646 6301 54698 6353
rect 55030 6227 55082 6279
rect 58102 6301 58154 6353
rect 58870 6227 58922 6279
rect 44182 6079 44234 6131
rect 51094 6079 51146 6131
rect 56278 6153 56330 6205
rect 19654 5968 19706 6020
rect 19718 5968 19770 6020
rect 19782 5968 19834 6020
rect 19846 5968 19898 6020
rect 50374 5968 50426 6020
rect 50438 5968 50490 6020
rect 50502 5968 50554 6020
rect 50566 5968 50618 6020
rect 5110 5783 5162 5835
rect 42742 5783 42794 5835
rect 57046 5783 57098 5835
rect 57718 5783 57770 5835
rect 15958 5709 16010 5761
rect 21622 5709 21674 5761
rect 1078 5635 1130 5687
rect 2902 5678 2954 5687
rect 2902 5644 2911 5678
rect 2911 5644 2945 5678
rect 2945 5644 2954 5678
rect 2902 5635 2954 5644
rect 4918 5635 4970 5687
rect 5206 5678 5258 5687
rect 5206 5644 5215 5678
rect 5215 5644 5249 5678
rect 5249 5644 5258 5678
rect 5206 5635 5258 5644
rect 6838 5678 6890 5687
rect 6838 5644 6847 5678
rect 6847 5644 6881 5678
rect 6881 5644 6890 5678
rect 6838 5635 6890 5644
rect 7222 5635 7274 5687
rect 8758 5635 8810 5687
rect 10198 5635 10250 5687
rect 10486 5635 10538 5687
rect 12598 5678 12650 5687
rect 12598 5644 12607 5678
rect 12607 5644 12641 5678
rect 12641 5644 12650 5678
rect 12598 5635 12650 5644
rect 13654 5635 13706 5687
rect 14998 5678 15050 5687
rect 14998 5644 15007 5678
rect 15007 5644 15041 5678
rect 15041 5644 15050 5678
rect 14998 5635 15050 5644
rect 15862 5678 15914 5687
rect 15862 5644 15871 5678
rect 15871 5644 15905 5678
rect 15905 5644 15914 5678
rect 15862 5635 15914 5644
rect 16150 5635 16202 5687
rect 17302 5678 17354 5687
rect 17302 5644 17311 5678
rect 17311 5644 17345 5678
rect 17345 5644 17354 5678
rect 18742 5678 18794 5687
rect 17302 5635 17354 5644
rect 18742 5644 18751 5678
rect 18751 5644 18785 5678
rect 18785 5644 18794 5678
rect 18742 5635 18794 5644
rect 20182 5678 20234 5687
rect 20182 5644 20191 5678
rect 20191 5644 20225 5678
rect 20225 5644 20234 5678
rect 20182 5635 20234 5644
rect 20566 5635 20618 5687
rect 21718 5678 21770 5687
rect 21718 5644 21727 5678
rect 21727 5644 21761 5678
rect 21761 5644 21770 5678
rect 21718 5635 21770 5644
rect 26038 5709 26090 5761
rect 23158 5635 23210 5687
rect 23446 5635 23498 5687
rect 24598 5635 24650 5687
rect 26230 5678 26282 5687
rect 26230 5644 26239 5678
rect 26239 5644 26273 5678
rect 26273 5644 26282 5678
rect 26230 5635 26282 5644
rect 37462 5709 37514 5761
rect 27382 5635 27434 5687
rect 27862 5635 27914 5687
rect 28822 5635 28874 5687
rect 30262 5635 30314 5687
rect 30838 5635 30890 5687
rect 31702 5635 31754 5687
rect 33142 5678 33194 5687
rect 33142 5644 33151 5678
rect 33151 5644 33185 5678
rect 33185 5644 33194 5678
rect 33142 5635 33194 5644
rect 33238 5635 33290 5687
rect 34774 5635 34826 5687
rect 36118 5678 36170 5687
rect 36118 5644 36127 5678
rect 36127 5644 36161 5678
rect 36161 5644 36170 5678
rect 36118 5635 36170 5644
rect 36214 5635 36266 5687
rect 37558 5678 37610 5687
rect 37558 5644 37567 5678
rect 37567 5644 37601 5678
rect 37601 5644 37610 5678
rect 37558 5635 37610 5644
rect 39094 5678 39146 5687
rect 39094 5644 39103 5678
rect 39103 5644 39137 5678
rect 39137 5644 39146 5678
rect 39094 5635 39146 5644
rect 39286 5635 39338 5687
rect 40726 5635 40778 5687
rect 41782 5635 41834 5687
rect 42262 5635 42314 5687
rect 43222 5635 43274 5687
rect 43702 5635 43754 5687
rect 45142 5678 45194 5687
rect 45142 5644 45151 5678
rect 45151 5644 45185 5678
rect 45185 5644 45194 5678
rect 45142 5635 45194 5644
rect 46102 5635 46154 5687
rect 46678 5635 46730 5687
rect 47542 5635 47594 5687
rect 49078 5635 49130 5687
rect 49654 5678 49706 5687
rect 49654 5644 49663 5678
rect 49663 5644 49697 5678
rect 49697 5644 49706 5678
rect 49654 5635 49706 5644
rect 50710 5635 50762 5687
rect 52150 5678 52202 5687
rect 52150 5644 52159 5678
rect 52159 5644 52193 5678
rect 52193 5644 52202 5678
rect 52150 5635 52202 5644
rect 52534 5635 52586 5687
rect 53686 5678 53738 5687
rect 53686 5644 53695 5678
rect 53695 5644 53729 5678
rect 53729 5644 53738 5678
rect 53686 5635 53738 5644
rect 57430 5678 57482 5687
rect 5974 5604 6026 5613
rect 5974 5570 5983 5604
rect 5983 5570 6017 5604
rect 6017 5570 6026 5604
rect 5974 5561 6026 5570
rect 50806 5561 50858 5613
rect 53590 5561 53642 5613
rect 57430 5644 57439 5678
rect 57439 5644 57473 5678
rect 57473 5644 57482 5678
rect 57430 5635 57482 5644
rect 59638 5561 59690 5613
rect 7606 5487 7658 5539
rect 17590 5413 17642 5465
rect 17878 5413 17930 5465
rect 29494 5413 29546 5465
rect 33526 5413 33578 5465
rect 4294 5302 4346 5354
rect 4358 5302 4410 5354
rect 4422 5302 4474 5354
rect 4486 5302 4538 5354
rect 35014 5302 35066 5354
rect 35078 5302 35130 5354
rect 35142 5302 35194 5354
rect 35206 5302 35258 5354
rect 7126 5191 7178 5243
rect 38134 5191 38186 5243
rect 4726 5117 4778 5169
rect 11062 5117 11114 5169
rect 20470 5117 20522 5169
rect 3574 5043 3626 5095
rect 310 4969 362 5021
rect 1846 4969 1898 5021
rect 3094 5012 3146 5021
rect 3094 4978 3103 5012
rect 3103 4978 3137 5012
rect 3137 4978 3146 5012
rect 3094 4969 3146 4978
rect 4150 5012 4202 5021
rect 4150 4978 4159 5012
rect 4159 4978 4193 5012
rect 4193 4978 4202 5012
rect 4150 4969 4202 4978
rect 5398 5012 5450 5021
rect 5398 4978 5407 5012
rect 5407 4978 5441 5012
rect 5441 4978 5450 5012
rect 5398 4969 5450 4978
rect 6070 4969 6122 5021
rect 9238 5012 9290 5021
rect 9238 4978 9247 5012
rect 9247 4978 9281 5012
rect 9281 4978 9290 5012
rect 9238 4969 9290 4978
rect 10582 4969 10634 5021
rect 11062 4969 11114 5021
rect 11830 4969 11882 5021
rect 12982 5012 13034 5021
rect 12982 4978 12991 5012
rect 12991 4978 13025 5012
rect 13025 4978 13034 5012
rect 12982 4969 13034 4978
rect 13942 5012 13994 5021
rect 13942 4978 13951 5012
rect 13951 4978 13985 5012
rect 13985 4978 13994 5012
rect 13942 4969 13994 4978
rect 14422 4969 14474 5021
rect 14806 4969 14858 5021
rect 16438 4969 16490 5021
rect 17494 5012 17546 5021
rect 17494 4978 17503 5012
rect 17503 4978 17537 5012
rect 17537 4978 17546 5012
rect 17494 4969 17546 4978
rect 18262 5012 18314 5021
rect 18262 4978 18271 5012
rect 18271 4978 18305 5012
rect 18305 4978 18314 5012
rect 18262 4969 18314 4978
rect 19030 5012 19082 5021
rect 19030 4978 19039 5012
rect 19039 4978 19073 5012
rect 19073 4978 19082 5012
rect 19030 4969 19082 4978
rect 19126 4969 19178 5021
rect 20662 5012 20714 5021
rect 20662 4978 20671 5012
rect 20671 4978 20705 5012
rect 20705 4978 20714 5012
rect 20662 4969 20714 4978
rect 20854 4969 20906 5021
rect 22774 5012 22826 5021
rect 22774 4978 22783 5012
rect 22783 4978 22817 5012
rect 22817 4978 22826 5012
rect 22774 4969 22826 4978
rect 23542 5012 23594 5021
rect 23542 4978 23551 5012
rect 23551 4978 23585 5012
rect 23585 4978 23594 5012
rect 23542 4969 23594 4978
rect 25078 5012 25130 5021
rect 23062 4895 23114 4947
rect 25078 4978 25087 5012
rect 25087 4978 25121 5012
rect 25121 4978 25130 5012
rect 25078 4969 25130 4978
rect 25846 5012 25898 5021
rect 25846 4978 25855 5012
rect 25855 4978 25889 5012
rect 25889 4978 25898 5012
rect 25846 4969 25898 4978
rect 26614 5012 26666 5021
rect 26614 4978 26623 5012
rect 26623 4978 26657 5012
rect 26657 4978 26666 5012
rect 26614 4969 26666 4978
rect 28054 5012 28106 5021
rect 28054 4978 28063 5012
rect 28063 4978 28097 5012
rect 28097 4978 28106 5012
rect 28054 4969 28106 4978
rect 28918 5012 28970 5021
rect 28918 4978 28927 5012
rect 28927 4978 28961 5012
rect 28961 4978 28970 5012
rect 28918 4969 28970 4978
rect 29302 4969 29354 5021
rect 30358 5012 30410 5021
rect 30358 4978 30367 5012
rect 30367 4978 30401 5012
rect 30401 4978 30410 5012
rect 30358 4969 30410 4978
rect 30454 4969 30506 5021
rect 31894 5012 31946 5021
rect 31894 4978 31903 5012
rect 31903 4978 31937 5012
rect 31937 4978 31946 5012
rect 31894 4969 31946 4978
rect 33334 5012 33386 5021
rect 33334 4978 33343 5012
rect 33343 4978 33377 5012
rect 33377 4978 33386 5012
rect 33334 4969 33386 4978
rect 34102 5012 34154 5021
rect 34102 4978 34111 5012
rect 34111 4978 34145 5012
rect 34145 4978 34154 5012
rect 34102 4969 34154 4978
rect 34870 5012 34922 5021
rect 34870 4978 34879 5012
rect 34879 4978 34913 5012
rect 34913 4978 34922 5012
rect 34870 4969 34922 4978
rect 36406 5012 36458 5021
rect 34582 4895 34634 4947
rect 36406 4978 36415 5012
rect 36415 4978 36449 5012
rect 36449 4978 36458 5012
rect 36406 4969 36458 4978
rect 36694 4969 36746 5021
rect 38614 5012 38666 5021
rect 38614 4978 38623 5012
rect 38623 4978 38657 5012
rect 38657 4978 38666 5012
rect 38614 4969 38666 4978
rect 39382 5012 39434 5021
rect 39382 4978 39391 5012
rect 39391 4978 39425 5012
rect 39425 4978 39434 5012
rect 39382 4969 39434 4978
rect 40150 5012 40202 5021
rect 40150 4978 40159 5012
rect 40159 4978 40193 5012
rect 40193 4978 40202 5012
rect 40150 4969 40202 4978
rect 40918 5012 40970 5021
rect 40918 4978 40927 5012
rect 40927 4978 40961 5012
rect 40961 4978 40970 5012
rect 40918 4969 40970 4978
rect 41686 5012 41738 5021
rect 41686 4978 41695 5012
rect 41695 4978 41729 5012
rect 41729 4978 41738 5012
rect 41686 4969 41738 4978
rect 42070 4969 42122 5021
rect 43510 4969 43562 5021
rect 44758 5012 44810 5021
rect 44758 4978 44767 5012
rect 44767 4978 44801 5012
rect 44801 4978 44810 5012
rect 44758 4969 44810 4978
rect 45430 5012 45482 5021
rect 45430 4978 45439 5012
rect 45439 4978 45473 5012
rect 45473 4978 45482 5012
rect 45430 4969 45482 4978
rect 46198 5012 46250 5021
rect 46198 4978 46207 5012
rect 46207 4978 46241 5012
rect 46241 4978 46250 5012
rect 46198 4969 46250 4978
rect 46294 4969 46346 5021
rect 47638 4969 47690 5021
rect 49366 5012 49418 5021
rect 49366 4978 49375 5012
rect 49375 4978 49409 5012
rect 49409 4978 49418 5012
rect 49366 4969 49418 4978
rect 50422 5012 50474 5021
rect 50422 4978 50431 5012
rect 50431 4978 50465 5012
rect 50465 4978 50474 5012
rect 50422 4969 50474 4978
rect 50902 4969 50954 5021
rect 51862 5012 51914 5021
rect 51862 4978 51871 5012
rect 51871 4978 51905 5012
rect 51905 4978 51914 5012
rect 51862 4969 51914 4978
rect 51958 4969 52010 5021
rect 53302 4969 53354 5021
rect 57046 5012 57098 5021
rect 57046 4978 57055 5012
rect 57055 4978 57089 5012
rect 57089 4978 57098 5012
rect 57046 4969 57098 4978
rect 57814 4895 57866 4947
rect 2134 4747 2186 4799
rect 59254 4821 59306 4873
rect 19654 4636 19706 4688
rect 19718 4636 19770 4688
rect 19782 4636 19834 4688
rect 19846 4636 19898 4688
rect 50374 4636 50426 4688
rect 50438 4636 50490 4688
rect 50502 4636 50554 4688
rect 50566 4636 50618 4688
rect 11158 4525 11210 4577
rect 20470 4525 20522 4577
rect 38134 4568 38186 4577
rect 38134 4534 38143 4568
rect 38143 4534 38177 4568
rect 38177 4534 38186 4568
rect 38134 4525 38186 4534
rect 57334 4525 57386 4577
rect 10774 4451 10826 4503
rect 11446 4451 11498 4503
rect 790 4377 842 4429
rect 1174 4303 1226 4355
rect 1366 4229 1418 4281
rect 3766 4229 3818 4281
rect 4726 4303 4778 4355
rect 3478 4155 3530 4207
rect 4918 4155 4970 4207
rect 5110 4155 5162 4207
rect 7414 4346 7466 4355
rect 5686 4229 5738 4281
rect 7414 4312 7423 4346
rect 7423 4312 7457 4346
rect 7457 4312 7466 4346
rect 7414 4303 7466 4312
rect 9622 4346 9674 4355
rect 6454 4155 6506 4207
rect 9622 4312 9631 4346
rect 9631 4312 9665 4346
rect 9665 4312 9674 4346
rect 9622 4303 9674 4312
rect 10390 4346 10442 4355
rect 10390 4312 10399 4346
rect 10399 4312 10433 4346
rect 10433 4312 10442 4346
rect 10390 4303 10442 4312
rect 10774 4303 10826 4355
rect 9814 4229 9866 4281
rect 10198 4229 10250 4281
rect 11158 4155 11210 4207
rect 13558 4346 13610 4355
rect 11446 4229 11498 4281
rect 13558 4312 13567 4346
rect 13567 4312 13601 4346
rect 13601 4312 13610 4346
rect 13558 4303 13610 4312
rect 15478 4346 15530 4355
rect 15478 4312 15487 4346
rect 15487 4312 15521 4346
rect 15521 4312 15530 4346
rect 15478 4303 15530 4312
rect 15958 4303 16010 4355
rect 16246 4155 16298 4207
rect 982 4081 1034 4133
rect 2326 4081 2378 4133
rect 2422 4081 2474 4133
rect 5014 4081 5066 4133
rect 9046 4081 9098 4133
rect 11062 4081 11114 4133
rect 16918 4081 16970 4133
rect 20278 4346 20330 4355
rect 17686 4229 17738 4281
rect 20278 4312 20287 4346
rect 20287 4312 20321 4346
rect 20321 4312 20330 4346
rect 20278 4303 20330 4312
rect 21046 4346 21098 4355
rect 21046 4312 21055 4346
rect 21055 4312 21089 4346
rect 21089 4312 21098 4346
rect 21046 4303 21098 4312
rect 21814 4346 21866 4355
rect 21814 4312 21823 4346
rect 21823 4312 21857 4346
rect 21857 4312 21866 4346
rect 21814 4303 21866 4312
rect 23254 4346 23306 4355
rect 23254 4312 23263 4346
rect 23263 4312 23297 4346
rect 23297 4312 23306 4346
rect 23254 4303 23306 4312
rect 25462 4346 25514 4355
rect 22006 4229 22058 4281
rect 25462 4312 25471 4346
rect 25471 4312 25505 4346
rect 25505 4312 25514 4346
rect 25462 4303 25514 4312
rect 26134 4303 26186 4355
rect 26518 4303 26570 4355
rect 28342 4346 28394 4355
rect 28342 4312 28351 4346
rect 28351 4312 28385 4346
rect 28385 4312 28394 4346
rect 28342 4303 28394 4312
rect 29110 4346 29162 4355
rect 29110 4312 29119 4346
rect 29119 4312 29153 4346
rect 29153 4312 29162 4346
rect 29110 4303 29162 4312
rect 30934 4346 30986 4355
rect 30934 4312 30943 4346
rect 30943 4312 30977 4346
rect 30977 4312 30986 4346
rect 30934 4303 30986 4312
rect 31702 4346 31754 4355
rect 31702 4312 31711 4346
rect 31711 4312 31745 4346
rect 31745 4312 31754 4346
rect 31702 4303 31754 4312
rect 32758 4346 32810 4355
rect 32758 4312 32767 4346
rect 32767 4312 32801 4346
rect 32801 4312 32810 4346
rect 32758 4303 32810 4312
rect 33910 4346 33962 4355
rect 33910 4312 33919 4346
rect 33919 4312 33953 4346
rect 33953 4312 33962 4346
rect 33910 4303 33962 4312
rect 34582 4303 34634 4355
rect 34198 4229 34250 4281
rect 36790 4346 36842 4355
rect 36790 4312 36799 4346
rect 36799 4312 36833 4346
rect 36833 4312 36842 4346
rect 36790 4303 36842 4312
rect 37174 4229 37226 4281
rect 38998 4346 39050 4355
rect 38998 4312 39007 4346
rect 39007 4312 39041 4346
rect 39041 4312 39050 4346
rect 38998 4303 39050 4312
rect 39766 4346 39818 4355
rect 39766 4312 39775 4346
rect 39775 4312 39809 4346
rect 39809 4312 39818 4346
rect 39766 4303 39818 4312
rect 41974 4346 42026 4355
rect 41974 4312 41983 4346
rect 41983 4312 42017 4346
rect 42017 4312 42026 4346
rect 41974 4303 42026 4312
rect 42358 4303 42410 4355
rect 43414 4303 43466 4355
rect 44950 4346 45002 4355
rect 44950 4312 44959 4346
rect 44959 4312 44993 4346
rect 44993 4312 45002 4346
rect 44950 4303 45002 4312
rect 46774 4346 46826 4355
rect 46774 4312 46783 4346
rect 46783 4312 46817 4346
rect 46817 4312 46826 4346
rect 46774 4303 46826 4312
rect 44470 4229 44522 4281
rect 45142 4229 45194 4281
rect 47446 4229 47498 4281
rect 47830 4303 47882 4355
rect 52630 4346 52682 4355
rect 48598 4229 48650 4281
rect 43798 4155 43850 4207
rect 47158 4155 47210 4207
rect 48982 4155 49034 4207
rect 49942 4229 49994 4281
rect 50998 4229 51050 4281
rect 52630 4312 52639 4346
rect 52639 4312 52673 4346
rect 52673 4312 52682 4346
rect 52630 4303 52682 4312
rect 53014 4229 53066 4281
rect 54070 4303 54122 4355
rect 55606 4346 55658 4355
rect 55606 4312 55615 4346
rect 55615 4312 55649 4346
rect 55649 4312 55658 4346
rect 55606 4303 55658 4312
rect 56662 4303 56714 4355
rect 56854 4229 56906 4281
rect 59158 4229 59210 4281
rect 56374 4155 56426 4207
rect 58294 4155 58346 4207
rect 17878 4081 17930 4133
rect 20950 4081 21002 4133
rect 21526 4081 21578 4133
rect 22870 4081 22922 4133
rect 24982 4081 25034 4133
rect 26614 4081 26666 4133
rect 40054 4081 40106 4133
rect 41686 4081 41738 4133
rect 45334 4081 45386 4133
rect 46294 4081 46346 4133
rect 48118 4081 48170 4133
rect 49078 4081 49130 4133
rect 49174 4081 49226 4133
rect 50710 4081 50762 4133
rect 56278 4081 56330 4133
rect 58006 4081 58058 4133
rect 4294 3970 4346 4022
rect 4358 3970 4410 4022
rect 4422 3970 4474 4022
rect 4486 3970 4538 4022
rect 35014 3970 35066 4022
rect 35078 3970 35130 4022
rect 35142 3970 35194 4022
rect 35206 3970 35258 4022
rect 1942 3859 1994 3911
rect 2998 3859 3050 3911
rect 8278 3859 8330 3911
rect 10582 3859 10634 3911
rect 13174 3859 13226 3911
rect 14038 3859 14090 3911
rect 18166 3859 18218 3911
rect 18550 3902 18602 3911
rect 18550 3868 18559 3902
rect 18559 3868 18593 3902
rect 18593 3868 18602 3902
rect 18550 3859 18602 3868
rect 21238 3859 21290 3911
rect 22774 3859 22826 3911
rect 23926 3859 23978 3911
rect 25078 3859 25130 3911
rect 27478 3859 27530 3911
rect 28918 3859 28970 3911
rect 29014 3859 29066 3911
rect 30358 3859 30410 3911
rect 38518 3859 38570 3911
rect 40150 3859 40202 3911
rect 41302 3859 41354 3911
rect 41494 3859 41546 3911
rect 502 3785 554 3837
rect 1654 3785 1706 3837
rect 2326 3785 2378 3837
rect 3094 3785 3146 3837
rect 7894 3785 7946 3837
rect 9238 3785 9290 3837
rect 12022 3785 12074 3837
rect 13654 3785 13706 3837
rect 15286 3785 15338 3837
rect 16534 3785 16586 3837
rect 17302 3785 17354 3837
rect 19414 3785 19466 3837
rect 20662 3785 20714 3837
rect 24214 3785 24266 3837
rect 25846 3785 25898 3837
rect 26422 3785 26474 3837
rect 28054 3785 28106 3837
rect 29398 3785 29450 3837
rect 30454 3785 30506 3837
rect 33430 3785 33482 3837
rect 34870 3785 34922 3837
rect 35638 3785 35690 3837
rect 36406 3785 36458 3837
rect 37846 3785 37898 3837
rect 39382 3785 39434 3837
rect 2998 3711 3050 3763
rect 3286 3711 3338 3763
rect 3382 3711 3434 3763
rect 118 3637 170 3689
rect 1654 3637 1706 3689
rect 2710 3637 2762 3689
rect 28726 3711 28778 3763
rect 5590 3680 5642 3689
rect 3094 3489 3146 3541
rect 5590 3646 5599 3680
rect 5599 3646 5633 3680
rect 5633 3646 5642 3680
rect 5590 3637 5642 3646
rect 6358 3637 6410 3689
rect 7030 3637 7082 3689
rect 7798 3637 7850 3689
rect 8566 3637 8618 3689
rect 9334 3637 9386 3689
rect 8086 3563 8138 3615
rect 9718 3563 9770 3615
rect 5110 3489 5162 3541
rect 5974 3489 6026 3541
rect 10006 3489 10058 3541
rect 13174 3637 13226 3689
rect 13654 3680 13706 3689
rect 13654 3646 13663 3680
rect 13663 3646 13697 3680
rect 13697 3646 13706 3680
rect 13654 3637 13706 3646
rect 14038 3637 14090 3689
rect 14806 3637 14858 3689
rect 15286 3637 15338 3689
rect 17398 3637 17450 3689
rect 18070 3637 18122 3689
rect 18454 3637 18506 3689
rect 19222 3637 19274 3689
rect 20662 3637 20714 3689
rect 22102 3637 22154 3689
rect 22870 3637 22922 3689
rect 23638 3637 23690 3689
rect 24406 3637 24458 3689
rect 19990 3563 20042 3615
rect 24694 3563 24746 3615
rect 15094 3489 15146 3541
rect 598 3415 650 3467
rect 1462 3415 1514 3467
rect 3286 3415 3338 3467
rect 3958 3415 4010 3467
rect 17302 3415 17354 3467
rect 17494 3415 17546 3467
rect 25846 3489 25898 3541
rect 27286 3637 27338 3689
rect 37750 3711 37802 3763
rect 43798 3859 43850 3911
rect 43990 3859 44042 3911
rect 44758 3859 44810 3911
rect 46294 3859 46346 3911
rect 47638 3859 47690 3911
rect 48502 3859 48554 3911
rect 49654 3859 49706 3911
rect 51382 3859 51434 3911
rect 51862 3859 51914 3911
rect 55990 3859 56042 3911
rect 57910 3859 57962 3911
rect 44086 3785 44138 3837
rect 45430 3785 45482 3837
rect 46102 3785 46154 3837
rect 47062 3785 47114 3837
rect 49078 3785 49130 3837
rect 50038 3785 50090 3837
rect 45238 3711 45290 3763
rect 28054 3489 28106 3541
rect 29494 3563 29546 3615
rect 30454 3637 30506 3689
rect 31318 3637 31370 3689
rect 32470 3637 32522 3689
rect 33526 3637 33578 3689
rect 34294 3637 34346 3689
rect 34966 3637 35018 3689
rect 35734 3637 35786 3689
rect 36502 3637 36554 3689
rect 37942 3637 37994 3689
rect 38710 3637 38762 3689
rect 32854 3563 32906 3615
rect 33718 3563 33770 3615
rect 28918 3489 28970 3541
rect 29782 3489 29834 3541
rect 30454 3489 30506 3541
rect 31894 3489 31946 3541
rect 35926 3489 35978 3541
rect 36694 3489 36746 3541
rect 39382 3489 39434 3541
rect 36022 3415 36074 3467
rect 36214 3415 36266 3467
rect 37078 3415 37130 3467
rect 38614 3415 38666 3467
rect 40150 3415 40202 3467
rect 41014 3637 41066 3689
rect 41590 3563 41642 3615
rect 42742 3637 42794 3689
rect 43798 3563 43850 3615
rect 44566 3563 44618 3615
rect 46006 3563 46058 3615
rect 47158 3637 47210 3689
rect 48214 3637 48266 3689
rect 50710 3637 50762 3689
rect 50806 3637 50858 3689
rect 51286 3637 51338 3689
rect 52054 3637 52106 3689
rect 53398 3637 53450 3689
rect 47638 3563 47690 3615
rect 48406 3563 48458 3615
rect 54358 3563 54410 3615
rect 55318 3637 55370 3689
rect 55894 3563 55946 3615
rect 44758 3489 44810 3541
rect 46198 3489 46250 3541
rect 51286 3489 51338 3541
rect 51574 3489 51626 3541
rect 52054 3489 52106 3541
rect 52246 3489 52298 3541
rect 56278 3489 56330 3541
rect 42550 3415 42602 3467
rect 43510 3415 43562 3467
rect 19654 3304 19706 3356
rect 19718 3304 19770 3356
rect 19782 3304 19834 3356
rect 19846 3304 19898 3356
rect 50374 3304 50426 3356
rect 50438 3304 50490 3356
rect 50502 3304 50554 3356
rect 50566 3304 50618 3356
rect 1462 3193 1514 3245
rect 2230 3193 2282 3245
rect 3958 3193 4010 3245
rect 5206 3193 5258 3245
rect 12310 3193 12362 3245
rect 13078 3193 13130 3245
rect 13270 3236 13322 3245
rect 13270 3202 13279 3236
rect 13279 3202 13313 3236
rect 13313 3202 13322 3236
rect 13270 3193 13322 3202
rect 13366 3193 13418 3245
rect 14134 3193 14186 3245
rect 17590 3193 17642 3245
rect 20950 3193 21002 3245
rect 22774 3193 22826 3245
rect 23158 3193 23210 3245
rect 28246 3193 28298 3245
rect 29302 3193 29354 3245
rect 31894 3193 31946 3245
rect 33334 3193 33386 3245
rect 33814 3193 33866 3245
rect 35062 3193 35114 3245
rect 36694 3193 36746 3245
rect 37558 3193 37610 3245
rect 41494 3193 41546 3245
rect 41782 3193 41834 3245
rect 43318 3236 43370 3245
rect 43318 3202 43327 3236
rect 43327 3202 43361 3236
rect 43361 3202 43370 3236
rect 43318 3193 43370 3202
rect 214 3119 266 3171
rect 1750 3119 1802 3171
rect 12214 3119 12266 3171
rect 12982 3119 13034 3171
rect 13750 3119 13802 3171
rect 17782 3119 17834 3171
rect 19798 3119 19850 3171
rect 20182 3119 20234 3171
rect 22390 3119 22442 3171
rect 23542 3119 23594 3171
rect 25366 3119 25418 3171
rect 26230 3119 26282 3171
rect 32662 3119 32714 3171
rect 34102 3119 34154 3171
rect 34678 3119 34730 3171
rect 35350 3119 35402 3171
rect 36214 3119 36266 3171
rect 13078 3045 13130 3097
rect 17494 3045 17546 3097
rect 18358 3045 18410 3097
rect 19606 3045 19658 3097
rect 22 2971 74 3023
rect 694 2897 746 2949
rect 2134 2897 2186 2949
rect 4918 3014 4970 3023
rect 4918 2980 4927 3014
rect 4927 2980 4961 3014
rect 4961 2980 4970 3014
rect 4918 2971 4970 2980
rect 5206 2971 5258 3023
rect 5974 2971 6026 3023
rect 6742 2897 6794 2949
rect 8182 2971 8234 3023
rect 8950 2897 9002 2949
rect 11734 2971 11786 3023
rect 12406 2971 12458 3023
rect 12982 3014 13034 3023
rect 12982 2980 12991 3014
rect 12991 2980 13025 3014
rect 13025 2980 13034 3014
rect 12982 2971 13034 2980
rect 13366 2971 13418 3023
rect 14518 2971 14570 3023
rect 16630 3014 16682 3023
rect 16630 2980 16639 3014
rect 16639 2980 16673 3014
rect 16673 2980 16682 3014
rect 16630 2971 16682 2980
rect 17014 2971 17066 3023
rect 15382 2897 15434 2949
rect 16438 2897 16490 2949
rect 17686 2897 17738 2949
rect 18838 2971 18890 3023
rect 20950 3045 21002 3097
rect 21718 3045 21770 3097
rect 22486 3045 22538 3097
rect 21430 2971 21482 3023
rect 25078 3045 25130 3097
rect 24022 2971 24074 3023
rect 27670 3045 27722 3097
rect 26902 2971 26954 3023
rect 30550 3045 30602 3097
rect 29878 2971 29930 3023
rect 32086 3045 32138 3097
rect 32278 2971 32330 3023
rect 33142 2971 33194 3023
rect 33334 3045 33386 3097
rect 35446 3045 35498 3097
rect 35350 2971 35402 3023
rect 36118 2971 36170 3023
rect 39670 3119 39722 3171
rect 40918 3119 40970 3171
rect 41110 3119 41162 3171
rect 42070 3119 42122 3171
rect 38326 3045 38378 3097
rect 37558 2971 37610 3023
rect 41206 3045 41258 3097
rect 40534 2971 40586 3023
rect 17974 2897 18026 2949
rect 18262 2897 18314 2949
rect 18358 2897 18410 2949
rect 19030 2897 19082 2949
rect 37750 2897 37802 2949
rect 38134 2897 38186 2949
rect 39094 2897 39146 2949
rect 41782 2897 41834 2949
rect 43318 2971 43370 3023
rect 44182 3193 44234 3245
rect 55318 3193 55370 3245
rect 55510 3193 55562 3245
rect 44374 3119 44426 3171
rect 58198 3193 58250 3245
rect 57718 3119 57770 3171
rect 59446 3119 59498 3171
rect 44182 3045 44234 3097
rect 52438 3045 52490 3097
rect 44374 2897 44426 2949
rect 45622 2971 45674 3023
rect 46390 2897 46442 2949
rect 49654 2971 49706 3023
rect 51478 2971 51530 3023
rect 52246 2897 52298 2949
rect 53782 2971 53834 3023
rect 52918 2897 52970 2949
rect 53686 2897 53738 2949
rect 54838 2897 54890 2949
rect 16822 2749 16874 2801
rect 27766 2749 27818 2801
rect 27958 2749 28010 2801
rect 32950 2792 33002 2801
rect 32950 2758 32959 2792
rect 32959 2758 32993 2792
rect 32993 2758 33002 2792
rect 32950 2749 33002 2758
rect 50038 2823 50090 2875
rect 52822 2749 52874 2801
rect 54454 2792 54506 2801
rect 54454 2758 54463 2792
rect 54463 2758 54497 2792
rect 54497 2758 54506 2792
rect 54454 2749 54506 2758
rect 4294 2638 4346 2690
rect 4358 2638 4410 2690
rect 4422 2638 4474 2690
rect 4486 2638 4538 2690
rect 35014 2638 35066 2690
rect 35078 2638 35130 2690
rect 35142 2638 35194 2690
rect 35206 2638 35258 2690
rect 3958 2527 4010 2579
rect 4246 2527 4298 2579
rect 4342 2527 4394 2579
rect 4822 2527 4874 2579
rect 7990 2527 8042 2579
rect 32950 2527 33002 2579
rect 35158 2527 35210 2579
rect 35542 2527 35594 2579
rect 5782 2453 5834 2505
rect 54454 2453 54506 2505
rect 20182 2379 20234 2431
rect 20854 2379 20906 2431
rect 4726 2009 4778 2061
rect 5302 2009 5354 2061
rect 4534 1861 4586 1913
rect 4822 1861 4874 1913
rect 30358 1713 30410 1765
rect 31510 1713 31562 1765
rect 34870 1713 34922 1765
rect 35638 1713 35690 1765
rect 41014 1713 41066 1765
rect 41302 1713 41354 1765
rect 54358 1713 54410 1765
rect 54646 1713 54698 1765
rect 35638 1565 35690 1617
rect 35926 1565 35978 1617
rect 36310 1491 36362 1543
rect 50518 1491 50570 1543
rect 51094 1491 51146 1543
rect 33238 1417 33290 1469
rect 33718 1417 33770 1469
rect 34678 1417 34730 1469
rect 35446 1417 35498 1469
rect 45430 1417 45482 1469
rect 45718 1417 45770 1469
rect 50710 1417 50762 1469
rect 50902 1417 50954 1469
rect 43318 1269 43370 1321
rect 43990 1269 44042 1321
rect 50902 1269 50954 1321
rect 51574 1269 51626 1321
rect 36310 1121 36362 1173
rect 45142 1047 45194 1099
rect 45334 1047 45386 1099
rect 43030 899 43082 951
rect 44374 899 44426 951
<< metal2 >>
rect 212 59200 268 60000
rect 692 59200 748 60000
rect 1172 59200 1228 60000
rect 1748 59200 1804 60000
rect 2228 59200 2284 60000
rect 2804 59200 2860 60000
rect 3284 59200 3340 60000
rect 3860 59200 3916 60000
rect 4340 59200 4396 60000
rect 4916 59200 4972 60000
rect 5396 59200 5452 60000
rect 5972 59200 6028 60000
rect 6452 59200 6508 60000
rect 7028 59200 7084 60000
rect 7508 59200 7564 60000
rect 8084 59200 8140 60000
rect 8564 59200 8620 60000
rect 9140 59200 9196 60000
rect 9620 59200 9676 60000
rect 10196 59200 10252 60000
rect 10676 59200 10732 60000
rect 11252 59200 11308 60000
rect 11732 59200 11788 60000
rect 12308 59200 12364 60000
rect 12788 59200 12844 60000
rect 13364 59200 13420 60000
rect 13844 59200 13900 60000
rect 14420 59200 14476 60000
rect 14900 59200 14956 60000
rect 15380 59200 15436 60000
rect 15956 59200 16012 60000
rect 16436 59200 16492 60000
rect 17012 59200 17068 60000
rect 17492 59200 17548 60000
rect 18068 59200 18124 60000
rect 18548 59200 18604 60000
rect 19124 59200 19180 60000
rect 19604 59200 19660 60000
rect 20180 59200 20236 60000
rect 20660 59200 20716 60000
rect 21236 59200 21292 60000
rect 21716 59200 21772 60000
rect 22292 59200 22348 60000
rect 22772 59200 22828 60000
rect 23348 59200 23404 60000
rect 23828 59200 23884 60000
rect 24404 59200 24460 60000
rect 24884 59200 24940 60000
rect 25460 59200 25516 60000
rect 25940 59200 25996 60000
rect 26516 59200 26572 60000
rect 26996 59200 27052 60000
rect 27572 59200 27628 60000
rect 28052 59200 28108 60000
rect 28628 59200 28684 60000
rect 29108 59200 29164 60000
rect 29684 59200 29740 60000
rect 30164 59200 30220 60000
rect 30644 59200 30700 60000
rect 31220 59200 31276 60000
rect 31700 59200 31756 60000
rect 32276 59200 32332 60000
rect 32756 59200 32812 60000
rect 33332 59200 33388 60000
rect 33812 59200 33868 60000
rect 34388 59200 34444 60000
rect 34868 59200 34924 60000
rect 35444 59200 35500 60000
rect 35924 59200 35980 60000
rect 36500 59200 36556 60000
rect 36980 59200 37036 60000
rect 37556 59200 37612 60000
rect 38036 59200 38092 60000
rect 38612 59200 38668 60000
rect 39092 59200 39148 60000
rect 39668 59200 39724 60000
rect 40148 59200 40204 60000
rect 40724 59200 40780 60000
rect 41204 59200 41260 60000
rect 41780 59200 41836 60000
rect 42260 59200 42316 60000
rect 42836 59200 42892 60000
rect 43316 59200 43372 60000
rect 43892 59200 43948 60000
rect 44372 59200 44428 60000
rect 44948 59200 45004 60000
rect 45428 59200 45484 60000
rect 45908 59200 45964 60000
rect 46484 59200 46540 60000
rect 46964 59200 47020 60000
rect 47540 59200 47596 60000
rect 48020 59200 48076 60000
rect 48596 59200 48652 60000
rect 49076 59200 49132 60000
rect 49652 59200 49708 60000
rect 50132 59200 50188 60000
rect 50708 59200 50764 60000
rect 51188 59200 51244 60000
rect 51764 59200 51820 60000
rect 52244 59200 52300 60000
rect 52820 59200 52876 60000
rect 53300 59200 53356 60000
rect 53876 59200 53932 60000
rect 54356 59200 54412 60000
rect 54932 59200 54988 60000
rect 55412 59200 55468 60000
rect 55988 59200 56044 60000
rect 56468 59200 56524 60000
rect 57044 59200 57100 60000
rect 57524 59200 57580 60000
rect 58100 59200 58156 60000
rect 58580 59200 58636 60000
rect 59156 59200 59212 60000
rect 59636 59200 59692 60000
rect 226 56975 254 59200
rect 214 56969 266 56975
rect 214 56911 266 56917
rect 706 56531 734 59200
rect 694 56525 746 56531
rect 694 56467 746 56473
rect 1186 55717 1214 59200
rect 1762 57049 1790 59200
rect 1750 57043 1802 57049
rect 1750 56985 1802 56991
rect 2038 56895 2090 56901
rect 2038 56837 2090 56843
rect 1750 56229 1802 56235
rect 1750 56171 1802 56177
rect 1174 55711 1226 55717
rect 1174 55653 1226 55659
rect 1762 50907 1790 56171
rect 1846 55415 1898 55421
rect 1846 55357 1898 55363
rect 1750 50901 1802 50907
rect 1750 50843 1802 50849
rect 1858 28115 1886 55357
rect 1846 28109 1898 28115
rect 1846 28051 1898 28057
rect 1750 16269 1802 16275
rect 1750 16211 1802 16217
rect 1762 8431 1790 16211
rect 1750 8425 1802 8431
rect 1750 8367 1802 8373
rect 1654 8277 1706 8283
rect 1654 8219 1706 8225
rect 1462 7685 1514 7691
rect 1462 7627 1514 7633
rect 1078 5687 1130 5693
rect 1078 5629 1130 5635
rect 310 5021 362 5027
rect 310 4963 362 4969
rect 118 3689 170 3695
rect 118 3631 170 3637
rect 22 3023 74 3029
rect 22 2965 74 2971
rect 34 800 62 2965
rect 130 800 158 3631
rect 214 3171 266 3177
rect 214 3113 266 3119
rect 226 800 254 3113
rect 322 800 350 4963
rect 790 4429 842 4435
rect 790 4371 842 4377
rect 502 3837 554 3843
rect 502 3779 554 3785
rect 514 800 542 3779
rect 598 3467 650 3473
rect 598 3409 650 3415
rect 610 800 638 3409
rect 694 2949 746 2955
rect 694 2891 746 2897
rect 706 800 734 2891
rect 802 800 830 4371
rect 982 4133 1034 4139
rect 982 4075 1034 4081
rect 994 800 1022 4075
rect 1090 800 1118 5629
rect 1174 4355 1226 4361
rect 1174 4297 1226 4303
rect 1186 800 1214 4297
rect 1366 4281 1418 4287
rect 1366 4223 1418 4229
rect 1378 800 1406 4223
rect 1474 3473 1502 7627
rect 1666 7214 1694 8219
rect 2050 7214 2078 56837
rect 2242 56531 2270 59200
rect 2818 56531 2846 59200
rect 3298 57049 3326 59200
rect 3286 57043 3338 57049
rect 3286 56985 3338 56991
rect 3574 56895 3626 56901
rect 3574 56837 3626 56843
rect 2230 56525 2282 56531
rect 2230 56467 2282 56473
rect 2806 56525 2858 56531
rect 2806 56467 2858 56473
rect 2518 56229 2570 56235
rect 2518 56171 2570 56177
rect 3382 56229 3434 56235
rect 3382 56171 3434 56177
rect 2134 54157 2186 54163
rect 2134 54099 2186 54105
rect 2146 7913 2174 54099
rect 2422 37433 2474 37439
rect 2422 37375 2474 37381
rect 2326 32105 2378 32111
rect 2326 32047 2378 32053
rect 2338 11835 2366 32047
rect 2326 11829 2378 11835
rect 2326 11771 2378 11777
rect 2434 8431 2462 37375
rect 2530 37069 2558 56171
rect 3286 52899 3338 52905
rect 3286 52841 3338 52847
rect 2710 48089 2762 48095
rect 2710 48031 2762 48037
rect 2722 47873 2750 48031
rect 2710 47867 2762 47873
rect 2710 47809 2762 47815
rect 2518 37063 2570 37069
rect 2518 37005 2570 37011
rect 2614 22263 2666 22269
rect 2614 22205 2666 22211
rect 2626 21751 2654 22205
rect 2614 21745 2666 21751
rect 2614 21687 2666 21693
rect 3298 8431 3326 52841
rect 3394 20567 3422 56171
rect 3382 20561 3434 20567
rect 3382 20503 3434 20509
rect 2422 8425 2474 8431
rect 2422 8367 2474 8373
rect 3286 8425 3338 8431
rect 3286 8367 3338 8373
rect 3286 8277 3338 8283
rect 3286 8219 3338 8225
rect 2230 8203 2282 8209
rect 2230 8145 2282 8151
rect 2134 7907 2186 7913
rect 2134 7849 2186 7855
rect 1666 7186 1790 7214
rect 2050 7186 2174 7214
rect 1654 7019 1706 7025
rect 1654 6961 1706 6967
rect 1558 6353 1610 6359
rect 1558 6295 1610 6301
rect 1462 3467 1514 3473
rect 1462 3409 1514 3415
rect 1462 3245 1514 3251
rect 1462 3187 1514 3193
rect 1474 800 1502 3187
rect 1570 800 1598 6295
rect 1666 3843 1694 6961
rect 1654 3837 1706 3843
rect 1654 3779 1706 3785
rect 1654 3689 1706 3695
rect 1654 3631 1706 3637
rect 1666 800 1694 3631
rect 1762 3177 1790 7186
rect 2038 6353 2090 6359
rect 2038 6295 2090 6301
rect 1846 5021 1898 5027
rect 1846 4963 1898 4969
rect 1750 3171 1802 3177
rect 1750 3113 1802 3119
rect 1858 800 1886 4963
rect 1942 3911 1994 3917
rect 1942 3853 1994 3859
rect 1954 800 1982 3853
rect 2050 800 2078 6295
rect 2146 4805 2174 7186
rect 2134 4799 2186 4805
rect 2134 4741 2186 4747
rect 2242 3251 2270 8145
rect 2326 7463 2378 7469
rect 2326 7405 2378 7411
rect 2998 7463 3050 7469
rect 2998 7405 3050 7411
rect 2338 4139 2366 7405
rect 2518 7019 2570 7025
rect 2518 6961 2570 6967
rect 2326 4133 2378 4139
rect 2326 4075 2378 4081
rect 2422 4133 2474 4139
rect 2422 4075 2474 4081
rect 2326 3837 2378 3843
rect 2326 3779 2378 3785
rect 2230 3245 2282 3251
rect 2230 3187 2282 3193
rect 2134 2949 2186 2955
rect 2134 2891 2186 2897
rect 2146 800 2174 2891
rect 2338 800 2366 3779
rect 2434 800 2462 4075
rect 2530 800 2558 6961
rect 2902 5687 2954 5693
rect 2902 5629 2954 5635
rect 2710 3689 2762 3695
rect 2710 3631 2762 3637
rect 2722 800 2750 3631
rect 2914 2900 2942 5629
rect 3010 3917 3038 7405
rect 3190 6353 3242 6359
rect 3190 6295 3242 6301
rect 3094 5021 3146 5027
rect 3094 4963 3146 4969
rect 2998 3911 3050 3917
rect 2998 3853 3050 3859
rect 3106 3843 3134 4963
rect 3094 3837 3146 3843
rect 3094 3779 3146 3785
rect 2998 3763 3050 3769
rect 2998 3705 3050 3711
rect 2818 2872 2942 2900
rect 2818 800 2846 2872
rect 3010 2752 3038 3705
rect 3094 3541 3146 3547
rect 3094 3483 3146 3489
rect 2914 2724 3038 2752
rect 2914 800 2942 2724
rect 3106 1864 3134 3483
rect 3010 1836 3134 1864
rect 3010 800 3038 1836
rect 3202 800 3230 6295
rect 3298 3769 3326 8219
rect 3586 5101 3614 56837
rect 3874 56531 3902 59200
rect 4354 57614 4382 59200
rect 4354 57586 4670 57614
rect 4268 57304 4564 57324
rect 4324 57302 4348 57304
rect 4404 57302 4428 57304
rect 4484 57302 4508 57304
rect 4346 57250 4348 57302
rect 4410 57250 4422 57302
rect 4484 57250 4486 57302
rect 4324 57248 4348 57250
rect 4404 57248 4428 57250
rect 4484 57248 4508 57250
rect 4268 57228 4564 57248
rect 3862 56525 3914 56531
rect 3862 56467 3914 56473
rect 3766 56303 3818 56309
rect 3766 56245 3818 56251
rect 3670 42095 3722 42101
rect 3670 42037 3722 42043
rect 3682 7913 3710 42037
rect 3778 16571 3806 56245
rect 4268 55972 4564 55992
rect 4324 55970 4348 55972
rect 4404 55970 4428 55972
rect 4484 55970 4508 55972
rect 4346 55918 4348 55970
rect 4410 55918 4422 55970
rect 4484 55918 4486 55970
rect 4324 55916 4348 55918
rect 4404 55916 4428 55918
rect 4484 55916 4508 55918
rect 4268 55896 4564 55916
rect 4642 55717 4670 57586
rect 4930 56975 4958 59200
rect 4918 56969 4970 56975
rect 4918 56911 4970 56917
rect 5110 56895 5162 56901
rect 5110 56837 5162 56843
rect 4630 55711 4682 55717
rect 4630 55653 4682 55659
rect 4630 55563 4682 55569
rect 4630 55505 4682 55511
rect 4268 54640 4564 54660
rect 4324 54638 4348 54640
rect 4404 54638 4428 54640
rect 4484 54638 4508 54640
rect 4346 54586 4348 54638
rect 4410 54586 4422 54638
rect 4484 54586 4486 54638
rect 4324 54584 4348 54586
rect 4404 54584 4428 54586
rect 4484 54584 4508 54586
rect 4268 54564 4564 54584
rect 4268 53308 4564 53328
rect 4324 53306 4348 53308
rect 4404 53306 4428 53308
rect 4484 53306 4508 53308
rect 4346 53254 4348 53306
rect 4410 53254 4422 53306
rect 4484 53254 4486 53306
rect 4324 53252 4348 53254
rect 4404 53252 4428 53254
rect 4484 53252 4508 53254
rect 4268 53232 4564 53252
rect 4268 51976 4564 51996
rect 4324 51974 4348 51976
rect 4404 51974 4428 51976
rect 4484 51974 4508 51976
rect 4346 51922 4348 51974
rect 4410 51922 4422 51974
rect 4484 51922 4486 51974
rect 4324 51920 4348 51922
rect 4404 51920 4428 51922
rect 4484 51920 4508 51922
rect 4268 51900 4564 51920
rect 4268 50644 4564 50664
rect 4324 50642 4348 50644
rect 4404 50642 4428 50644
rect 4484 50642 4508 50644
rect 4346 50590 4348 50642
rect 4410 50590 4422 50642
rect 4484 50590 4486 50642
rect 4324 50588 4348 50590
rect 4404 50588 4428 50590
rect 4484 50588 4508 50590
rect 4268 50568 4564 50588
rect 4268 49312 4564 49332
rect 4324 49310 4348 49312
rect 4404 49310 4428 49312
rect 4484 49310 4508 49312
rect 4346 49258 4348 49310
rect 4410 49258 4422 49310
rect 4484 49258 4486 49310
rect 4324 49256 4348 49258
rect 4404 49256 4428 49258
rect 4484 49256 4508 49258
rect 4268 49236 4564 49256
rect 4268 47980 4564 48000
rect 4324 47978 4348 47980
rect 4404 47978 4428 47980
rect 4484 47978 4508 47980
rect 4346 47926 4348 47978
rect 4410 47926 4422 47978
rect 4484 47926 4486 47978
rect 4324 47924 4348 47926
rect 4404 47924 4428 47926
rect 4484 47924 4508 47926
rect 4268 47904 4564 47924
rect 4268 46648 4564 46668
rect 4324 46646 4348 46648
rect 4404 46646 4428 46648
rect 4484 46646 4508 46648
rect 4346 46594 4348 46646
rect 4410 46594 4422 46646
rect 4484 46594 4486 46646
rect 4324 46592 4348 46594
rect 4404 46592 4428 46594
rect 4484 46592 4508 46594
rect 4268 46572 4564 46592
rect 4268 45316 4564 45336
rect 4324 45314 4348 45316
rect 4404 45314 4428 45316
rect 4484 45314 4508 45316
rect 4346 45262 4348 45314
rect 4410 45262 4422 45314
rect 4484 45262 4486 45314
rect 4324 45260 4348 45262
rect 4404 45260 4428 45262
rect 4484 45260 4508 45262
rect 4268 45240 4564 45260
rect 4268 43984 4564 44004
rect 4324 43982 4348 43984
rect 4404 43982 4428 43984
rect 4484 43982 4508 43984
rect 4346 43930 4348 43982
rect 4410 43930 4422 43982
rect 4484 43930 4486 43982
rect 4324 43928 4348 43930
rect 4404 43928 4428 43930
rect 4484 43928 4508 43930
rect 4268 43908 4564 43928
rect 4268 42652 4564 42672
rect 4324 42650 4348 42652
rect 4404 42650 4428 42652
rect 4484 42650 4508 42652
rect 4346 42598 4348 42650
rect 4410 42598 4422 42650
rect 4484 42598 4486 42650
rect 4324 42596 4348 42598
rect 4404 42596 4428 42598
rect 4484 42596 4508 42598
rect 4268 42576 4564 42596
rect 4268 41320 4564 41340
rect 4324 41318 4348 41320
rect 4404 41318 4428 41320
rect 4484 41318 4508 41320
rect 4346 41266 4348 41318
rect 4410 41266 4422 41318
rect 4484 41266 4486 41318
rect 4324 41264 4348 41266
rect 4404 41264 4428 41266
rect 4484 41264 4508 41266
rect 4268 41244 4564 41264
rect 4268 39988 4564 40008
rect 4324 39986 4348 39988
rect 4404 39986 4428 39988
rect 4484 39986 4508 39988
rect 4346 39934 4348 39986
rect 4410 39934 4422 39986
rect 4484 39934 4486 39986
rect 4324 39932 4348 39934
rect 4404 39932 4428 39934
rect 4484 39932 4508 39934
rect 4268 39912 4564 39932
rect 4268 38656 4564 38676
rect 4324 38654 4348 38656
rect 4404 38654 4428 38656
rect 4484 38654 4508 38656
rect 4346 38602 4348 38654
rect 4410 38602 4422 38654
rect 4484 38602 4486 38654
rect 4324 38600 4348 38602
rect 4404 38600 4428 38602
rect 4484 38600 4508 38602
rect 4268 38580 4564 38600
rect 4268 37324 4564 37344
rect 4324 37322 4348 37324
rect 4404 37322 4428 37324
rect 4484 37322 4508 37324
rect 4346 37270 4348 37322
rect 4410 37270 4422 37322
rect 4484 37270 4486 37322
rect 4324 37268 4348 37270
rect 4404 37268 4428 37270
rect 4484 37268 4508 37270
rect 4268 37248 4564 37268
rect 4268 35992 4564 36012
rect 4324 35990 4348 35992
rect 4404 35990 4428 35992
rect 4484 35990 4508 35992
rect 4346 35938 4348 35990
rect 4410 35938 4422 35990
rect 4484 35938 4486 35990
rect 4324 35936 4348 35938
rect 4404 35936 4428 35938
rect 4484 35936 4508 35938
rect 4268 35916 4564 35936
rect 4268 34660 4564 34680
rect 4324 34658 4348 34660
rect 4404 34658 4428 34660
rect 4484 34658 4508 34660
rect 4346 34606 4348 34658
rect 4410 34606 4422 34658
rect 4484 34606 4486 34658
rect 4324 34604 4348 34606
rect 4404 34604 4428 34606
rect 4484 34604 4508 34606
rect 4268 34584 4564 34604
rect 4268 33328 4564 33348
rect 4324 33326 4348 33328
rect 4404 33326 4428 33328
rect 4484 33326 4508 33328
rect 4346 33274 4348 33326
rect 4410 33274 4422 33326
rect 4484 33274 4486 33326
rect 4324 33272 4348 33274
rect 4404 33272 4428 33274
rect 4484 33272 4508 33274
rect 4268 33252 4564 33272
rect 4642 33134 4670 55505
rect 4642 33106 4862 33134
rect 4268 31996 4564 32016
rect 4324 31994 4348 31996
rect 4404 31994 4428 31996
rect 4484 31994 4508 31996
rect 4346 31942 4348 31994
rect 4410 31942 4422 31994
rect 4484 31942 4486 31994
rect 4324 31940 4348 31942
rect 4404 31940 4428 31942
rect 4484 31940 4508 31942
rect 4268 31920 4564 31940
rect 4268 30664 4564 30684
rect 4324 30662 4348 30664
rect 4404 30662 4428 30664
rect 4484 30662 4508 30664
rect 4346 30610 4348 30662
rect 4410 30610 4422 30662
rect 4484 30610 4486 30662
rect 4324 30608 4348 30610
rect 4404 30608 4428 30610
rect 4484 30608 4508 30610
rect 4268 30588 4564 30608
rect 4268 29332 4564 29352
rect 4324 29330 4348 29332
rect 4404 29330 4428 29332
rect 4484 29330 4508 29332
rect 4346 29278 4348 29330
rect 4410 29278 4422 29330
rect 4484 29278 4486 29330
rect 4324 29276 4348 29278
rect 4404 29276 4428 29278
rect 4484 29276 4508 29278
rect 4268 29256 4564 29276
rect 4268 28000 4564 28020
rect 4324 27998 4348 28000
rect 4404 27998 4428 28000
rect 4484 27998 4508 28000
rect 4346 27946 4348 27998
rect 4410 27946 4422 27998
rect 4484 27946 4486 27998
rect 4324 27944 4348 27946
rect 4404 27944 4428 27946
rect 4484 27944 4508 27946
rect 4268 27924 4564 27944
rect 4268 26668 4564 26688
rect 4324 26666 4348 26668
rect 4404 26666 4428 26668
rect 4484 26666 4508 26668
rect 4346 26614 4348 26666
rect 4410 26614 4422 26666
rect 4484 26614 4486 26666
rect 4324 26612 4348 26614
rect 4404 26612 4428 26614
rect 4484 26612 4508 26614
rect 4268 26592 4564 26612
rect 4268 25336 4564 25356
rect 4324 25334 4348 25336
rect 4404 25334 4428 25336
rect 4484 25334 4508 25336
rect 4346 25282 4348 25334
rect 4410 25282 4422 25334
rect 4484 25282 4486 25334
rect 4324 25280 4348 25282
rect 4404 25280 4428 25282
rect 4484 25280 4508 25282
rect 4268 25260 4564 25280
rect 4268 24004 4564 24024
rect 4324 24002 4348 24004
rect 4404 24002 4428 24004
rect 4484 24002 4508 24004
rect 4346 23950 4348 24002
rect 4410 23950 4422 24002
rect 4484 23950 4486 24002
rect 4324 23948 4348 23950
rect 4404 23948 4428 23950
rect 4484 23948 4508 23950
rect 4268 23928 4564 23948
rect 4268 22672 4564 22692
rect 4324 22670 4348 22672
rect 4404 22670 4428 22672
rect 4484 22670 4508 22672
rect 4346 22618 4348 22670
rect 4410 22618 4422 22670
rect 4484 22618 4486 22670
rect 4324 22616 4348 22618
rect 4404 22616 4428 22618
rect 4484 22616 4508 22618
rect 4268 22596 4564 22616
rect 4268 21340 4564 21360
rect 4324 21338 4348 21340
rect 4404 21338 4428 21340
rect 4484 21338 4508 21340
rect 4346 21286 4348 21338
rect 4410 21286 4422 21338
rect 4484 21286 4486 21338
rect 4324 21284 4348 21286
rect 4404 21284 4428 21286
rect 4484 21284 4508 21286
rect 4268 21264 4564 21284
rect 4268 20008 4564 20028
rect 4324 20006 4348 20008
rect 4404 20006 4428 20008
rect 4484 20006 4508 20008
rect 4346 19954 4348 20006
rect 4410 19954 4422 20006
rect 4484 19954 4486 20006
rect 4324 19952 4348 19954
rect 4404 19952 4428 19954
rect 4484 19952 4508 19954
rect 4268 19932 4564 19952
rect 4268 18676 4564 18696
rect 4324 18674 4348 18676
rect 4404 18674 4428 18676
rect 4484 18674 4508 18676
rect 4346 18622 4348 18674
rect 4410 18622 4422 18674
rect 4484 18622 4486 18674
rect 4324 18620 4348 18622
rect 4404 18620 4428 18622
rect 4484 18620 4508 18622
rect 4268 18600 4564 18620
rect 4268 17344 4564 17364
rect 4324 17342 4348 17344
rect 4404 17342 4428 17344
rect 4484 17342 4508 17344
rect 4346 17290 4348 17342
rect 4410 17290 4422 17342
rect 4484 17290 4486 17342
rect 4324 17288 4348 17290
rect 4404 17288 4428 17290
rect 4484 17288 4508 17290
rect 4268 17268 4564 17288
rect 3766 16565 3818 16571
rect 3766 16507 3818 16513
rect 3862 16195 3914 16201
rect 3862 16137 3914 16143
rect 3874 15905 3902 16137
rect 4268 16012 4564 16032
rect 4324 16010 4348 16012
rect 4404 16010 4428 16012
rect 4484 16010 4508 16012
rect 4346 15958 4348 16010
rect 4410 15958 4422 16010
rect 4484 15958 4486 16010
rect 4324 15956 4348 15958
rect 4404 15956 4428 15958
rect 4484 15956 4508 15958
rect 4268 15936 4564 15956
rect 3862 15899 3914 15905
rect 3862 15841 3914 15847
rect 4268 14680 4564 14700
rect 4324 14678 4348 14680
rect 4404 14678 4428 14680
rect 4484 14678 4508 14680
rect 4346 14626 4348 14678
rect 4410 14626 4422 14678
rect 4484 14626 4486 14678
rect 4324 14624 4348 14626
rect 4404 14624 4428 14626
rect 4484 14624 4508 14626
rect 4268 14604 4564 14624
rect 4268 13348 4564 13368
rect 4324 13346 4348 13348
rect 4404 13346 4428 13348
rect 4484 13346 4508 13348
rect 4346 13294 4348 13346
rect 4410 13294 4422 13346
rect 4484 13294 4486 13346
rect 4324 13292 4348 13294
rect 4404 13292 4428 13294
rect 4484 13292 4508 13294
rect 4268 13272 4564 13292
rect 4834 12974 4862 33106
rect 4738 12946 4862 12974
rect 4268 12016 4564 12036
rect 4324 12014 4348 12016
rect 4404 12014 4428 12016
rect 4484 12014 4508 12016
rect 4346 11962 4348 12014
rect 4410 11962 4422 12014
rect 4484 11962 4486 12014
rect 4324 11960 4348 11962
rect 4404 11960 4428 11962
rect 4484 11960 4508 11962
rect 4268 11940 4564 11960
rect 4268 10684 4564 10704
rect 4324 10682 4348 10684
rect 4404 10682 4428 10684
rect 4484 10682 4508 10684
rect 4346 10630 4348 10682
rect 4410 10630 4422 10682
rect 4484 10630 4486 10682
rect 4324 10628 4348 10630
rect 4404 10628 4428 10630
rect 4484 10628 4508 10630
rect 4268 10608 4564 10628
rect 4268 9352 4564 9372
rect 4324 9350 4348 9352
rect 4404 9350 4428 9352
rect 4484 9350 4508 9352
rect 4346 9298 4348 9350
rect 4410 9298 4422 9350
rect 4484 9298 4486 9350
rect 4324 9296 4348 9298
rect 4404 9296 4428 9298
rect 4484 9296 4508 9298
rect 4268 9276 4564 9296
rect 4268 8020 4564 8040
rect 4324 8018 4348 8020
rect 4404 8018 4428 8020
rect 4484 8018 4508 8020
rect 4346 7966 4348 8018
rect 4410 7966 4422 8018
rect 4484 7966 4486 8018
rect 4324 7964 4348 7966
rect 4404 7964 4428 7966
rect 4484 7964 4508 7966
rect 4268 7944 4564 7964
rect 3670 7907 3722 7913
rect 3670 7849 3722 7855
rect 3958 7463 4010 7469
rect 3958 7405 4010 7411
rect 4054 7463 4106 7469
rect 4054 7405 4106 7411
rect 3670 6797 3722 6803
rect 3670 6739 3722 6745
rect 3574 5095 3626 5101
rect 3574 5037 3626 5043
rect 3478 4207 3530 4213
rect 3478 4149 3530 4155
rect 3286 3763 3338 3769
rect 3286 3705 3338 3711
rect 3382 3763 3434 3769
rect 3382 3705 3434 3711
rect 3286 3467 3338 3473
rect 3286 3409 3338 3415
rect 3298 800 3326 3409
rect 3394 800 3422 3705
rect 3490 800 3518 4149
rect 3682 800 3710 6739
rect 3862 6353 3914 6359
rect 3862 6295 3914 6301
rect 3766 4281 3818 4287
rect 3766 4223 3818 4229
rect 3778 800 3806 4223
rect 3874 800 3902 6295
rect 3970 3473 3998 7405
rect 3958 3467 4010 3473
rect 3958 3409 4010 3415
rect 3958 3245 4010 3251
rect 3958 3187 4010 3193
rect 3970 2585 3998 3187
rect 3958 2579 4010 2585
rect 3958 2521 4010 2527
rect 4066 800 4094 7405
rect 4268 6688 4564 6708
rect 4324 6686 4348 6688
rect 4404 6686 4428 6688
rect 4484 6686 4508 6688
rect 4346 6634 4348 6686
rect 4410 6634 4422 6686
rect 4484 6634 4486 6686
rect 4324 6632 4348 6634
rect 4404 6632 4428 6634
rect 4484 6632 4508 6634
rect 4268 6612 4564 6632
rect 4630 6353 4682 6359
rect 4630 6295 4682 6301
rect 4268 5356 4564 5376
rect 4324 5354 4348 5356
rect 4404 5354 4428 5356
rect 4484 5354 4508 5356
rect 4346 5302 4348 5354
rect 4410 5302 4422 5354
rect 4484 5302 4486 5354
rect 4324 5300 4348 5302
rect 4404 5300 4428 5302
rect 4484 5300 4508 5302
rect 4268 5280 4564 5300
rect 4150 5021 4202 5027
rect 4150 4963 4202 4969
rect 4162 800 4190 4963
rect 4268 4024 4564 4044
rect 4324 4022 4348 4024
rect 4404 4022 4428 4024
rect 4484 4022 4508 4024
rect 4346 3970 4348 4022
rect 4410 3970 4422 4022
rect 4484 3970 4486 4022
rect 4324 3968 4348 3970
rect 4404 3968 4428 3970
rect 4484 3968 4508 3970
rect 4268 3948 4564 3968
rect 4268 2692 4564 2712
rect 4324 2690 4348 2692
rect 4404 2690 4428 2692
rect 4484 2690 4508 2692
rect 4346 2638 4348 2690
rect 4410 2638 4422 2690
rect 4484 2638 4486 2690
rect 4324 2636 4348 2638
rect 4404 2636 4428 2638
rect 4484 2636 4508 2638
rect 4268 2616 4564 2636
rect 4246 2579 4298 2585
rect 4246 2521 4298 2527
rect 4342 2579 4394 2585
rect 4342 2521 4394 2527
rect 4258 800 4286 2521
rect 4354 800 4382 2521
rect 4642 2456 4670 6295
rect 4738 5175 4766 12946
rect 4822 8203 4874 8209
rect 4822 8145 4874 8151
rect 4726 5169 4778 5175
rect 4726 5111 4778 5117
rect 4726 4355 4778 4361
rect 4726 4297 4778 4303
rect 4450 2428 4670 2456
rect 4450 2012 4478 2428
rect 4738 2160 4766 4297
rect 4834 2585 4862 8145
rect 5122 7007 5150 56837
rect 5410 56531 5438 59200
rect 5986 56531 6014 59200
rect 6466 56975 6494 59200
rect 6454 56969 6506 56975
rect 6454 56911 6506 56917
rect 7042 56531 7070 59200
rect 7222 56895 7274 56901
rect 7222 56837 7274 56843
rect 5398 56525 5450 56531
rect 5398 56467 5450 56473
rect 5974 56525 6026 56531
rect 5974 56467 6026 56473
rect 7030 56525 7082 56531
rect 7030 56467 7082 56473
rect 5206 56229 5258 56235
rect 5206 56171 5258 56177
rect 5590 56229 5642 56235
rect 5590 56171 5642 56177
rect 6358 56229 6410 56235
rect 6358 56171 6410 56177
rect 6454 56229 6506 56235
rect 6454 56171 6506 56177
rect 5218 11243 5246 56171
rect 5302 54971 5354 54977
rect 5302 54913 5354 54919
rect 5314 12974 5342 54913
rect 5602 36255 5630 56171
rect 6370 38253 6398 56171
rect 6358 38247 6410 38253
rect 6358 38189 6410 38195
rect 6466 37439 6494 56171
rect 6454 37433 6506 37439
rect 6454 37375 6506 37381
rect 5590 36249 5642 36255
rect 5590 36191 5642 36197
rect 6742 32105 6794 32111
rect 6742 32047 6794 32053
rect 6646 30773 6698 30779
rect 6646 30715 6698 30721
rect 6070 17453 6122 17459
rect 6070 17395 6122 17401
rect 5314 12946 5438 12974
rect 5206 11237 5258 11243
rect 5206 11179 5258 11185
rect 5302 7463 5354 7469
rect 5302 7405 5354 7411
rect 5122 6979 5246 7007
rect 5110 6945 5162 6951
rect 5110 6887 5162 6893
rect 5014 6871 5066 6877
rect 5014 6813 5066 6819
rect 4918 5687 4970 5693
rect 4918 5629 4970 5635
rect 4930 4213 4958 5629
rect 4918 4207 4970 4213
rect 4918 4149 4970 4155
rect 5026 4139 5054 6813
rect 5122 5841 5150 6887
rect 5218 6211 5246 6979
rect 5206 6205 5258 6211
rect 5206 6147 5258 6153
rect 5110 5835 5162 5841
rect 5110 5777 5162 5783
rect 5206 5687 5258 5693
rect 5206 5629 5258 5635
rect 5110 4207 5162 4213
rect 5110 4149 5162 4155
rect 5014 4133 5066 4139
rect 5014 4075 5066 4081
rect 5122 3640 5150 4149
rect 5026 3612 5150 3640
rect 4918 3023 4970 3029
rect 4918 2965 4970 2971
rect 4822 2579 4874 2585
rect 4822 2521 4874 2527
rect 4738 2132 4862 2160
rect 4726 2061 4778 2067
rect 4450 1984 4670 2012
rect 4726 2003 4778 2009
rect 4534 1913 4586 1919
rect 4534 1855 4586 1861
rect 4546 800 4574 1855
rect 4642 800 4670 1984
rect 4738 800 4766 2003
rect 4834 1919 4862 2132
rect 4822 1913 4874 1919
rect 4822 1855 4874 1861
rect 4930 800 4958 2965
rect 5026 800 5054 3612
rect 5110 3541 5162 3547
rect 5110 3483 5162 3489
rect 5122 800 5150 3483
rect 5218 3251 5246 5629
rect 5206 3245 5258 3251
rect 5206 3187 5258 3193
rect 5206 3023 5258 3029
rect 5206 2965 5258 2971
rect 5218 800 5246 2965
rect 5314 2067 5342 7405
rect 5410 6581 5438 12946
rect 5686 7759 5738 7765
rect 5686 7701 5738 7707
rect 5590 7611 5642 7617
rect 5590 7553 5642 7559
rect 5602 7247 5630 7553
rect 5590 7241 5642 7247
rect 5590 7183 5642 7189
rect 5398 6575 5450 6581
rect 5398 6517 5450 6523
rect 5494 6131 5546 6137
rect 5494 6073 5546 6079
rect 5398 5021 5450 5027
rect 5398 4963 5450 4969
rect 5302 2061 5354 2067
rect 5302 2003 5354 2009
rect 5410 800 5438 4963
rect 5506 800 5534 6073
rect 5698 4380 5726 7701
rect 6082 7099 6110 17395
rect 6070 7093 6122 7099
rect 6070 7035 6122 7041
rect 5878 6945 5930 6951
rect 5878 6887 5930 6893
rect 6550 6945 6602 6951
rect 6550 6887 6602 6893
rect 5698 4352 5822 4380
rect 5686 4281 5738 4287
rect 5686 4223 5738 4229
rect 5590 3689 5642 3695
rect 5590 3631 5642 3637
rect 5602 800 5630 3631
rect 5698 800 5726 4223
rect 5794 2511 5822 4352
rect 5782 2505 5834 2511
rect 5782 2447 5834 2453
rect 5890 800 5918 6887
rect 6262 6427 6314 6433
rect 6262 6369 6314 6375
rect 5974 5613 6026 5619
rect 5974 5555 6026 5561
rect 5986 3547 6014 5555
rect 6070 5021 6122 5027
rect 6070 4963 6122 4969
rect 5974 3541 6026 3547
rect 5974 3483 6026 3489
rect 5974 3023 6026 3029
rect 5974 2965 6026 2971
rect 5986 800 6014 2965
rect 6082 800 6110 4963
rect 6274 800 6302 6369
rect 6454 4207 6506 4213
rect 6454 4149 6506 4155
rect 6358 3689 6410 3695
rect 6358 3631 6410 3637
rect 6370 800 6398 3631
rect 6466 800 6494 4149
rect 6562 800 6590 6887
rect 6658 6581 6686 30715
rect 6754 10799 6782 32047
rect 7234 25840 7262 56837
rect 7522 55717 7550 59200
rect 8098 56975 8126 59200
rect 8086 56969 8138 56975
rect 8086 56911 8138 56917
rect 8578 56531 8606 59200
rect 8566 56525 8618 56531
rect 8566 56467 8618 56473
rect 9154 55717 9182 59200
rect 9634 57049 9662 59200
rect 9622 57043 9674 57049
rect 9622 56985 9674 56991
rect 9814 56747 9866 56753
rect 9814 56689 9866 56695
rect 7510 55711 7562 55717
rect 7510 55653 7562 55659
rect 9142 55711 9194 55717
rect 9142 55653 9194 55659
rect 7702 55563 7754 55569
rect 7702 55505 7754 55511
rect 8470 55563 8522 55569
rect 8470 55505 8522 55511
rect 9238 55563 9290 55569
rect 9238 55505 9290 55511
rect 7714 45505 7742 55505
rect 8482 54829 8510 55505
rect 8470 54823 8522 54829
rect 8470 54765 8522 54771
rect 9046 49199 9098 49205
rect 9046 49141 9098 49147
rect 7702 45499 7754 45505
rect 7702 45441 7754 45447
rect 7318 30995 7370 31001
rect 7318 30937 7370 30943
rect 7330 30261 7358 30937
rect 7318 30255 7370 30261
rect 7318 30197 7370 30203
rect 8566 26777 8618 26783
rect 8566 26719 8618 26725
rect 8230 26555 8282 26561
rect 8230 26497 8282 26503
rect 8242 26376 8270 26497
rect 8578 26432 8606 26719
rect 8530 26404 8606 26432
rect 8530 26376 8558 26404
rect 8230 26370 8282 26376
rect 8230 26312 8282 26318
rect 8518 26370 8570 26376
rect 8518 26312 8570 26318
rect 6946 25812 7262 25840
rect 6946 12974 6974 25812
rect 8086 24853 8138 24859
rect 8086 24795 8138 24801
rect 8098 24563 8126 24795
rect 8086 24557 8138 24563
rect 8086 24499 8138 24505
rect 8086 23521 8138 23527
rect 8086 23463 8138 23469
rect 8098 23231 8126 23463
rect 8086 23225 8138 23231
rect 8086 23167 8138 23173
rect 7894 22781 7946 22787
rect 7894 22723 7946 22729
rect 7126 20931 7178 20937
rect 7126 20873 7178 20879
rect 7138 20419 7166 20873
rect 7126 20413 7178 20419
rect 7126 20355 7178 20361
rect 6946 12946 7166 12974
rect 6742 10793 6794 10799
rect 6742 10735 6794 10741
rect 6934 6945 6986 6951
rect 6934 6887 6986 6893
rect 6646 6575 6698 6581
rect 6646 6517 6698 6523
rect 6838 5687 6890 5693
rect 6838 5629 6890 5635
rect 6742 2949 6794 2955
rect 6742 2891 6794 2897
rect 6754 800 6782 2891
rect 6850 800 6878 5629
rect 6946 800 6974 6887
rect 7138 6433 7166 12946
rect 7798 12199 7850 12205
rect 7798 12141 7850 12147
rect 7810 11835 7838 12141
rect 7798 11829 7850 11835
rect 7798 11771 7850 11777
rect 7906 10300 7934 22723
rect 8086 22189 8138 22195
rect 8086 22131 8138 22137
rect 8098 21899 8126 22131
rect 8086 21893 8138 21899
rect 8086 21835 8138 21841
rect 8086 21523 8138 21529
rect 8086 21465 8138 21471
rect 8098 20863 8126 21465
rect 8086 20857 8138 20863
rect 8086 20799 8138 20805
rect 8758 19451 8810 19457
rect 8758 19393 8810 19399
rect 8770 19235 8798 19393
rect 8758 19229 8810 19235
rect 8758 19171 8810 19177
rect 8086 11015 8138 11021
rect 8086 10957 8138 10963
rect 8098 10355 8126 10957
rect 8278 10867 8330 10873
rect 8278 10809 8330 10815
rect 7810 10272 7934 10300
rect 8086 10349 8138 10355
rect 8086 10291 8138 10297
rect 7810 8431 7838 10272
rect 8182 9905 8234 9911
rect 8182 9847 8234 9853
rect 8086 9683 8138 9689
rect 8086 9625 8138 9631
rect 8098 9097 8126 9625
rect 8194 9171 8222 9847
rect 8182 9165 8234 9171
rect 8182 9107 8234 9113
rect 8086 9091 8138 9097
rect 8086 9033 8138 9039
rect 8194 8968 8222 9107
rect 8098 8940 8222 8968
rect 8098 8801 8126 8940
rect 8086 8795 8138 8801
rect 8086 8737 8138 8743
rect 7798 8425 7850 8431
rect 7798 8367 7850 8373
rect 8290 8357 8318 10809
rect 8374 9757 8426 9763
rect 8374 9699 8426 9705
rect 8386 9097 8414 9699
rect 8662 9609 8714 9615
rect 8662 9551 8714 9557
rect 8374 9091 8426 9097
rect 8374 9033 8426 9039
rect 7606 8351 7658 8357
rect 7606 8293 7658 8299
rect 8278 8351 8330 8357
rect 8278 8293 8330 8299
rect 7618 7913 7646 8293
rect 7702 8277 7754 8283
rect 7702 8219 7754 8225
rect 7606 7907 7658 7913
rect 7606 7849 7658 7855
rect 7318 6871 7370 6877
rect 7318 6813 7370 6819
rect 7126 6427 7178 6433
rect 7126 6369 7178 6375
rect 7126 6279 7178 6285
rect 7126 6221 7178 6227
rect 7138 5249 7166 6221
rect 7222 5687 7274 5693
rect 7222 5629 7274 5635
rect 7126 5243 7178 5249
rect 7126 5185 7178 5191
rect 7030 3689 7082 3695
rect 7030 3631 7082 3637
rect 7042 800 7070 3631
rect 7234 800 7262 5629
rect 7330 800 7358 6813
rect 7606 5539 7658 5545
rect 7606 5481 7658 5487
rect 7414 4355 7466 4361
rect 7414 4297 7466 4303
rect 7426 800 7454 4297
rect 7618 800 7646 5481
rect 7714 800 7742 8219
rect 8086 8129 8138 8135
rect 8086 8071 8138 8077
rect 8098 7765 8126 8071
rect 8086 7759 8138 7765
rect 8086 7701 8138 7707
rect 8290 7636 8318 8293
rect 8674 7784 8702 9551
rect 9058 7913 9086 49141
rect 9142 29441 9194 29447
rect 9142 29383 9194 29389
rect 9154 29151 9182 29383
rect 9142 29145 9194 29151
rect 9142 29087 9194 29093
rect 9142 28775 9194 28781
rect 9142 28717 9194 28723
rect 9154 28559 9182 28717
rect 9142 28553 9194 28559
rect 9142 28495 9194 28501
rect 9046 7907 9098 7913
rect 9046 7849 9098 7855
rect 8386 7765 8702 7784
rect 9058 7765 9086 7849
rect 8374 7759 8702 7765
rect 8426 7756 8702 7759
rect 9046 7759 9098 7765
rect 8374 7701 8426 7707
rect 9046 7701 9098 7707
rect 9142 7685 9194 7691
rect 8290 7608 8414 7636
rect 9142 7627 9194 7633
rect 8386 7469 8414 7608
rect 8374 7463 8426 7469
rect 8374 7405 8426 7411
rect 8758 7463 8810 7469
rect 8758 7405 8810 7411
rect 8770 7340 8798 7405
rect 8482 7312 8798 7340
rect 7798 6945 7850 6951
rect 7798 6887 7850 6893
rect 7810 4676 7838 6887
rect 7810 4648 8030 4676
rect 7894 3837 7946 3843
rect 7894 3779 7946 3785
rect 7798 3689 7850 3695
rect 7798 3631 7850 3637
rect 7810 800 7838 3631
rect 7906 800 7934 3779
rect 8002 2585 8030 4648
rect 8278 3911 8330 3917
rect 8278 3853 8330 3859
rect 8086 3615 8138 3621
rect 8086 3557 8138 3563
rect 7990 2579 8042 2585
rect 7990 2521 8042 2527
rect 8098 800 8126 3557
rect 8182 3023 8234 3029
rect 8182 2965 8234 2971
rect 8194 800 8222 2965
rect 8290 800 8318 3853
rect 8482 800 8510 7312
rect 8854 7167 8906 7173
rect 8854 7109 8906 7115
rect 8758 5687 8810 5693
rect 8758 5629 8810 5635
rect 8770 4232 8798 5629
rect 8674 4204 8798 4232
rect 8566 3689 8618 3695
rect 8566 3631 8618 3637
rect 8578 800 8606 3631
rect 8674 800 8702 4204
rect 8866 2894 8894 7109
rect 9046 4133 9098 4139
rect 9046 4075 9098 4081
rect 8770 2866 8894 2894
rect 8950 2949 9002 2955
rect 8950 2891 9002 2897
rect 8770 800 8798 2866
rect 8962 800 8990 2891
rect 9058 800 9086 4075
rect 9154 800 9182 7627
rect 9250 6507 9278 55505
rect 9430 50753 9482 50759
rect 9430 50695 9482 50701
rect 9334 19451 9386 19457
rect 9334 19393 9386 19399
rect 9346 19235 9374 19393
rect 9334 19229 9386 19235
rect 9334 19171 9386 19177
rect 9442 12974 9470 50695
rect 9622 20561 9674 20567
rect 9622 20503 9674 20509
rect 9634 20345 9662 20503
rect 9622 20339 9674 20345
rect 9622 20281 9674 20287
rect 9622 14937 9674 14943
rect 9622 14879 9674 14885
rect 9634 14573 9662 14879
rect 9622 14567 9674 14573
rect 9622 14509 9674 14515
rect 9442 12946 9662 12974
rect 9526 12125 9578 12131
rect 9526 12067 9578 12073
rect 9538 11761 9566 12067
rect 9526 11755 9578 11761
rect 9526 11697 9578 11703
rect 9526 11459 9578 11465
rect 9526 11401 9578 11407
rect 9538 11243 9566 11401
rect 9526 11237 9578 11243
rect 9526 11179 9578 11185
rect 9526 8277 9578 8283
rect 9526 8219 9578 8225
rect 9238 6501 9290 6507
rect 9238 6443 9290 6449
rect 9430 6353 9482 6359
rect 9430 6295 9482 6301
rect 9238 5021 9290 5027
rect 9238 4963 9290 4969
rect 9250 3843 9278 4963
rect 9238 3837 9290 3843
rect 9238 3779 9290 3785
rect 9334 3689 9386 3695
rect 9334 3631 9386 3637
rect 9346 2894 9374 3631
rect 9250 2866 9374 2894
rect 9250 800 9278 2866
rect 9442 800 9470 6295
rect 9538 800 9566 8219
rect 9634 7839 9662 12946
rect 9826 8135 9854 56689
rect 10210 56531 10238 59200
rect 10690 56531 10718 59200
rect 11266 57049 11294 59200
rect 11254 57043 11306 57049
rect 11254 56985 11306 56991
rect 11254 56895 11306 56901
rect 11254 56837 11306 56843
rect 10198 56525 10250 56531
rect 10198 56467 10250 56473
rect 10678 56525 10730 56531
rect 10678 56467 10730 56473
rect 10774 56229 10826 56235
rect 10774 56171 10826 56177
rect 10294 50457 10346 50463
rect 10294 50399 10346 50405
rect 10306 49723 10334 50399
rect 10294 49717 10346 49723
rect 10294 49659 10346 49665
rect 9910 34251 9962 34257
rect 9910 34193 9962 34199
rect 9922 8579 9950 34193
rect 10786 33134 10814 56171
rect 10786 33106 11006 33134
rect 10870 28553 10922 28559
rect 10870 28495 10922 28501
rect 10774 24779 10826 24785
rect 10774 24721 10826 24727
rect 10582 20117 10634 20123
rect 10582 20059 10634 20065
rect 10594 19827 10622 20059
rect 10582 19821 10634 19827
rect 10582 19763 10634 19769
rect 10486 11829 10538 11835
rect 10538 11789 10670 11817
rect 10486 11771 10538 11777
rect 10642 11687 10670 11789
rect 10630 11681 10682 11687
rect 10630 11623 10682 11629
rect 10678 10793 10730 10799
rect 10678 10735 10730 10741
rect 10690 10577 10718 10735
rect 10198 10571 10250 10577
rect 10198 10513 10250 10519
rect 10678 10571 10730 10577
rect 10678 10513 10730 10519
rect 9910 8573 9962 8579
rect 9910 8515 9962 8521
rect 9814 8129 9866 8135
rect 9814 8071 9866 8077
rect 9622 7833 9674 7839
rect 9622 7775 9674 7781
rect 10210 7691 10238 10513
rect 10678 9461 10730 9467
rect 10678 9403 10730 9409
rect 10690 9245 10718 9403
rect 10678 9239 10730 9245
rect 10678 9181 10730 9187
rect 10294 8425 10346 8431
rect 10294 8367 10346 8373
rect 10198 7685 10250 7691
rect 10198 7627 10250 7633
rect 9910 7463 9962 7469
rect 9910 7405 9962 7411
rect 9718 6945 9770 6951
rect 9718 6887 9770 6893
rect 9814 6945 9866 6951
rect 9814 6887 9866 6893
rect 9622 4355 9674 4361
rect 9622 4297 9674 4303
rect 9634 800 9662 4297
rect 9730 3621 9758 6887
rect 9826 6507 9854 6887
rect 9814 6501 9866 6507
rect 9814 6443 9866 6449
rect 9814 4281 9866 4287
rect 9814 4223 9866 4229
rect 9718 3615 9770 3621
rect 9718 3557 9770 3563
rect 9826 800 9854 4223
rect 9922 800 9950 7405
rect 10102 6353 10154 6359
rect 10102 6295 10154 6301
rect 10006 3541 10058 3547
rect 10006 3483 10058 3489
rect 10018 800 10046 3483
rect 10114 800 10142 6295
rect 10198 5687 10250 5693
rect 10198 5629 10250 5635
rect 10210 4287 10238 5629
rect 10198 4281 10250 4287
rect 10198 4223 10250 4229
rect 10306 800 10334 8367
rect 10582 8277 10634 8283
rect 10582 8219 10634 8225
rect 10678 8277 10730 8283
rect 10678 8219 10730 8225
rect 10594 8135 10622 8219
rect 10582 8129 10634 8135
rect 10582 8071 10634 8077
rect 10582 6945 10634 6951
rect 10582 6887 10634 6893
rect 10594 6581 10622 6887
rect 10582 6575 10634 6581
rect 10582 6517 10634 6523
rect 10486 5687 10538 5693
rect 10486 5629 10538 5635
rect 10390 4355 10442 4361
rect 10390 4297 10442 4303
rect 10402 800 10430 4297
rect 10498 800 10526 5629
rect 10582 5021 10634 5027
rect 10582 4963 10634 4969
rect 10594 3917 10622 4963
rect 10582 3911 10634 3917
rect 10582 3853 10634 3859
rect 10690 2894 10718 8219
rect 10786 4509 10814 24721
rect 10882 12974 10910 28495
rect 10978 24193 11006 33106
rect 11158 29441 11210 29447
rect 11158 29383 11210 29389
rect 11170 29151 11198 29383
rect 11158 29145 11210 29151
rect 11158 29087 11210 29093
rect 11158 24557 11210 24563
rect 11158 24499 11210 24505
rect 10966 24187 11018 24193
rect 10966 24129 11018 24135
rect 10882 12946 11102 12974
rect 10870 12199 10922 12205
rect 10870 12141 10922 12147
rect 10882 11835 10910 12141
rect 10870 11829 10922 11835
rect 10870 11771 10922 11777
rect 10966 7463 11018 7469
rect 10966 7405 11018 7411
rect 10870 6353 10922 6359
rect 10870 6295 10922 6301
rect 10774 4503 10826 4509
rect 10774 4445 10826 4451
rect 10774 4355 10826 4361
rect 10774 4297 10826 4303
rect 10594 2866 10718 2894
rect 10594 800 10622 2866
rect 10786 800 10814 4297
rect 10882 800 10910 6295
rect 10978 800 11006 7405
rect 11074 5175 11102 12946
rect 11062 5169 11114 5175
rect 11062 5111 11114 5117
rect 11062 5021 11114 5027
rect 11062 4963 11114 4969
rect 11074 4139 11102 4963
rect 11170 4583 11198 24499
rect 11266 7617 11294 56837
rect 11746 56531 11774 59200
rect 12322 56531 12350 59200
rect 12802 56975 12830 59200
rect 12790 56969 12842 56975
rect 12790 56911 12842 56917
rect 12982 56895 13034 56901
rect 12982 56837 13034 56843
rect 11734 56525 11786 56531
rect 11734 56467 11786 56473
rect 12310 56525 12362 56531
rect 12310 56467 12362 56473
rect 11926 56229 11978 56235
rect 11926 56171 11978 56177
rect 12694 56229 12746 56235
rect 12694 56171 12746 56177
rect 11938 52239 11966 56171
rect 12022 55193 12074 55199
rect 12022 55135 12074 55141
rect 11926 52233 11978 52239
rect 11926 52175 11978 52181
rect 11350 34769 11402 34775
rect 11350 34711 11402 34717
rect 11362 8431 11390 34711
rect 11446 24853 11498 24859
rect 11446 24795 11498 24801
rect 11350 8425 11402 8431
rect 11350 8367 11402 8373
rect 11350 8277 11402 8283
rect 11350 8219 11402 8225
rect 11254 7611 11306 7617
rect 11254 7553 11306 7559
rect 11254 7019 11306 7025
rect 11254 6961 11306 6967
rect 11158 4577 11210 4583
rect 11158 4519 11210 4525
rect 11158 4207 11210 4213
rect 11158 4149 11210 4155
rect 11062 4133 11114 4139
rect 11062 4075 11114 4081
rect 11170 800 11198 4149
rect 11266 800 11294 6961
rect 11362 800 11390 8219
rect 11458 4509 11486 24795
rect 11542 9535 11594 9541
rect 11542 9477 11594 9483
rect 11554 7173 11582 9477
rect 12034 9245 12062 55135
rect 12598 45425 12650 45431
rect 12598 45367 12650 45373
rect 12022 9239 12074 9245
rect 12022 9181 12074 9187
rect 12214 8573 12266 8579
rect 11746 8505 11966 8524
rect 12214 8515 12266 8521
rect 11734 8499 11978 8505
rect 11786 8496 11926 8499
rect 11734 8441 11786 8447
rect 11926 8441 11978 8447
rect 11542 7167 11594 7173
rect 11542 7109 11594 7115
rect 11638 6353 11690 6359
rect 11638 6295 11690 6301
rect 11446 4503 11498 4509
rect 11446 4445 11498 4451
rect 11446 4281 11498 4287
rect 11446 4223 11498 4229
rect 11458 800 11486 4223
rect 11650 800 11678 6295
rect 12226 5564 12254 8515
rect 12310 8277 12362 8283
rect 12310 8219 12362 8225
rect 12322 7691 12350 8219
rect 12610 7765 12638 45367
rect 12706 20567 12734 56171
rect 12994 30254 13022 56837
rect 13378 56531 13406 59200
rect 13366 56525 13418 56531
rect 13366 56467 13418 56473
rect 13750 56377 13802 56383
rect 13750 56319 13802 56325
rect 12994 30226 13310 30254
rect 12982 23891 13034 23897
rect 12982 23833 13034 23839
rect 12694 20561 12746 20567
rect 12694 20503 12746 20509
rect 12994 20174 13022 23833
rect 13282 23768 13310 30226
rect 13366 24113 13418 24119
rect 13366 24055 13418 24061
rect 13378 23897 13406 24055
rect 13366 23891 13418 23897
rect 13366 23833 13418 23839
rect 13282 23740 13406 23768
rect 13174 22189 13226 22195
rect 13174 22131 13226 22137
rect 12994 20146 13118 20174
rect 12982 15899 13034 15905
rect 12982 15841 13034 15847
rect 12994 9023 13022 15841
rect 12982 9017 13034 9023
rect 12982 8959 13034 8965
rect 12886 8277 12938 8283
rect 12886 8219 12938 8225
rect 12898 7784 12926 8219
rect 12598 7759 12650 7765
rect 12598 7701 12650 7707
rect 12694 7759 12746 7765
rect 12898 7756 13022 7784
rect 12694 7701 12746 7707
rect 12310 7685 12362 7691
rect 12310 7627 12362 7633
rect 12502 7611 12554 7617
rect 12502 7553 12554 7559
rect 12406 7463 12458 7469
rect 12406 7405 12458 7411
rect 12130 5536 12254 5564
rect 11830 5021 11882 5027
rect 11830 4963 11882 4969
rect 11734 3023 11786 3029
rect 11734 2965 11786 2971
rect 11746 800 11774 2965
rect 11842 800 11870 4963
rect 12022 3837 12074 3843
rect 12022 3779 12074 3785
rect 12034 800 12062 3779
rect 12130 800 12158 5536
rect 12310 3245 12362 3251
rect 12310 3187 12362 3193
rect 12214 3171 12266 3177
rect 12214 3113 12266 3119
rect 12226 800 12254 3113
rect 12322 800 12350 3187
rect 12418 3029 12446 7405
rect 12514 7247 12542 7553
rect 12502 7241 12554 7247
rect 12706 7192 12734 7701
rect 12994 7247 13022 7756
rect 12502 7183 12554 7189
rect 12610 7164 12734 7192
rect 12790 7241 12842 7247
rect 12790 7183 12842 7189
rect 12982 7241 13034 7247
rect 12982 7183 13034 7189
rect 12610 5860 12638 7164
rect 12694 7019 12746 7025
rect 12694 6961 12746 6967
rect 12514 5832 12638 5860
rect 12406 3023 12458 3029
rect 12406 2965 12458 2971
rect 12514 800 12542 5832
rect 12598 5687 12650 5693
rect 12598 5629 12650 5635
rect 12610 800 12638 5629
rect 12706 800 12734 6961
rect 12802 800 12830 7183
rect 13090 6581 13118 20146
rect 13078 6575 13130 6581
rect 13078 6517 13130 6523
rect 13078 6353 13130 6359
rect 13078 6295 13130 6301
rect 12982 5021 13034 5027
rect 12982 4963 13034 4969
rect 12994 3177 13022 4963
rect 13090 3251 13118 6295
rect 13186 3917 13214 22131
rect 13270 21893 13322 21899
rect 13270 21835 13322 21841
rect 13174 3911 13226 3917
rect 13174 3853 13226 3859
rect 13174 3689 13226 3695
rect 13174 3631 13226 3637
rect 13078 3245 13130 3251
rect 13078 3187 13130 3193
rect 12982 3171 13034 3177
rect 12982 3113 13034 3119
rect 13078 3097 13130 3103
rect 13078 3039 13130 3045
rect 12982 3023 13034 3029
rect 12982 2965 13034 2971
rect 12994 800 13022 2965
rect 13090 800 13118 3039
rect 13186 800 13214 3631
rect 13282 3251 13310 21835
rect 13378 9615 13406 23740
rect 13462 22115 13514 22121
rect 13462 22057 13514 22063
rect 13366 9609 13418 9615
rect 13366 9551 13418 9557
rect 13474 7214 13502 22057
rect 13654 20117 13706 20123
rect 13654 20059 13706 20065
rect 13666 8431 13694 20059
rect 13762 8949 13790 56319
rect 13858 55717 13886 59200
rect 14434 56975 14462 59200
rect 14422 56969 14474 56975
rect 14422 56911 14474 56917
rect 14914 56531 14942 59200
rect 14902 56525 14954 56531
rect 14902 56467 14954 56473
rect 15190 56303 15242 56309
rect 15190 56245 15242 56251
rect 15094 56229 15146 56235
rect 15094 56171 15146 56177
rect 13846 55711 13898 55717
rect 13846 55653 13898 55659
rect 14038 55563 14090 55569
rect 14038 55505 14090 55511
rect 13942 36323 13994 36329
rect 13942 36265 13994 36271
rect 13750 8943 13802 8949
rect 13750 8885 13802 8891
rect 13654 8425 13706 8431
rect 13654 8367 13706 8373
rect 13750 8203 13802 8209
rect 13750 8145 13802 8151
rect 13762 7839 13790 8145
rect 13750 7833 13802 7839
rect 13750 7775 13802 7781
rect 13378 7186 13502 7214
rect 13378 3251 13406 7186
rect 13462 6945 13514 6951
rect 13462 6887 13514 6893
rect 13270 3245 13322 3251
rect 13270 3187 13322 3193
rect 13366 3245 13418 3251
rect 13366 3187 13418 3193
rect 13366 3023 13418 3029
rect 13366 2965 13418 2971
rect 13378 800 13406 2965
rect 13474 800 13502 6887
rect 13954 6433 13982 36265
rect 14050 18125 14078 55505
rect 14134 23225 14186 23231
rect 14134 23167 14186 23173
rect 14038 18119 14090 18125
rect 14038 18061 14090 18067
rect 14038 6575 14090 6581
rect 14038 6517 14090 6523
rect 13942 6427 13994 6433
rect 13942 6369 13994 6375
rect 13750 6131 13802 6137
rect 13750 6073 13802 6079
rect 13942 6131 13994 6137
rect 13942 6073 13994 6079
rect 13654 5687 13706 5693
rect 13654 5629 13706 5635
rect 13558 4355 13610 4361
rect 13558 4297 13610 4303
rect 13570 800 13598 4297
rect 13666 3843 13694 5629
rect 13654 3837 13706 3843
rect 13654 3779 13706 3785
rect 13654 3689 13706 3695
rect 13654 3631 13706 3637
rect 13666 800 13694 3631
rect 13762 3177 13790 6073
rect 13954 5120 13982 6073
rect 13858 5092 13982 5120
rect 13750 3171 13802 3177
rect 13750 3113 13802 3119
rect 13858 800 13886 5092
rect 13942 5021 13994 5027
rect 13942 4963 13994 4969
rect 13954 800 13982 4963
rect 14050 3917 14078 6517
rect 14038 3911 14090 3917
rect 14038 3853 14090 3859
rect 14038 3689 14090 3695
rect 14038 3631 14090 3637
rect 14050 800 14078 3631
rect 14146 3251 14174 23167
rect 14710 16195 14762 16201
rect 14710 16137 14762 16143
rect 14614 6945 14666 6951
rect 14614 6887 14666 6893
rect 14230 6205 14282 6211
rect 14230 6147 14282 6153
rect 14134 3245 14186 3251
rect 14134 3187 14186 3193
rect 14242 3085 14270 6147
rect 14422 5021 14474 5027
rect 14422 4963 14474 4969
rect 14146 3057 14270 3085
rect 14146 800 14174 3057
rect 14434 2900 14462 4963
rect 14518 3023 14570 3029
rect 14518 2965 14570 2971
rect 14338 2872 14462 2900
rect 14338 800 14366 2872
rect 14530 1568 14558 2965
rect 14434 1540 14558 1568
rect 14434 800 14462 1540
rect 14626 1420 14654 6887
rect 14722 6433 14750 16137
rect 15106 14499 15134 56171
rect 15202 40547 15230 56245
rect 15394 56161 15422 59200
rect 15970 56975 15998 59200
rect 16450 57049 16478 59200
rect 16438 57043 16490 57049
rect 16438 56985 16490 56991
rect 15958 56969 16010 56975
rect 15958 56911 16010 56917
rect 16150 56895 16202 56901
rect 16150 56837 16202 56843
rect 15766 56229 15818 56235
rect 15766 56171 15818 56177
rect 15382 56155 15434 56161
rect 15382 56097 15434 56103
rect 15190 40541 15242 40547
rect 15190 40483 15242 40489
rect 15286 29071 15338 29077
rect 15286 29013 15338 29019
rect 15094 14493 15146 14499
rect 15094 14435 15146 14441
rect 15094 10793 15146 10799
rect 15094 10735 15146 10741
rect 15106 7099 15134 10735
rect 15298 7214 15326 29013
rect 15382 27665 15434 27671
rect 15382 27607 15434 27613
rect 15202 7186 15326 7214
rect 15094 7093 15146 7099
rect 15094 7035 15146 7041
rect 14710 6427 14762 6433
rect 14710 6369 14762 6375
rect 14902 6279 14954 6285
rect 14902 6221 14954 6227
rect 14806 5021 14858 5027
rect 14530 1392 14654 1420
rect 14722 4981 14806 5009
rect 14530 800 14558 1392
rect 14722 800 14750 4981
rect 14806 4963 14858 4969
rect 14806 3689 14858 3695
rect 14806 3631 14858 3637
rect 14818 800 14846 3631
rect 14914 800 14942 6221
rect 14998 5687 15050 5693
rect 14998 5629 15050 5635
rect 15010 800 15038 5629
rect 15202 3788 15230 7186
rect 15394 7007 15422 27607
rect 15478 22485 15530 22491
rect 15478 22427 15530 22433
rect 15298 6979 15422 7007
rect 15298 3843 15326 6979
rect 15382 6945 15434 6951
rect 15382 6887 15434 6893
rect 15106 3760 15230 3788
rect 15286 3837 15338 3843
rect 15286 3779 15338 3785
rect 15106 3547 15134 3760
rect 15286 3689 15338 3695
rect 15202 3649 15286 3677
rect 15094 3541 15146 3547
rect 15094 3483 15146 3489
rect 15202 800 15230 3649
rect 15286 3631 15338 3637
rect 15394 3492 15422 6887
rect 15490 6433 15518 22427
rect 15778 10873 15806 56171
rect 15958 40097 16010 40103
rect 15958 40039 16010 40045
rect 15862 39875 15914 39881
rect 15862 39817 15914 39823
rect 15766 10867 15818 10873
rect 15766 10809 15818 10815
rect 15874 7765 15902 39817
rect 15970 12372 15998 40039
rect 16054 23447 16106 23453
rect 16054 23389 16106 23395
rect 16066 12501 16094 23389
rect 16162 23054 16190 56837
rect 17026 56531 17054 59200
rect 17506 56975 17534 59200
rect 17494 56969 17546 56975
rect 17494 56911 17546 56917
rect 17974 56895 18026 56901
rect 17974 56837 18026 56843
rect 17014 56525 17066 56531
rect 17014 56467 17066 56473
rect 16534 56451 16586 56457
rect 16534 56393 16586 56399
rect 16438 42761 16490 42767
rect 16438 42703 16490 42709
rect 16450 42545 16478 42703
rect 16438 42539 16490 42545
rect 16438 42481 16490 42487
rect 16162 23026 16382 23054
rect 16246 20413 16298 20419
rect 16246 20355 16298 20361
rect 16150 16121 16202 16127
rect 16150 16063 16202 16069
rect 16162 15905 16190 16063
rect 16150 15899 16202 15905
rect 16150 15841 16202 15847
rect 16054 12495 16106 12501
rect 16054 12437 16106 12443
rect 15970 12344 16094 12372
rect 15958 12273 16010 12279
rect 15958 12215 16010 12221
rect 15862 7759 15914 7765
rect 15862 7701 15914 7707
rect 15670 7463 15722 7469
rect 15670 7405 15722 7411
rect 15478 6427 15530 6433
rect 15478 6369 15530 6375
rect 15478 4355 15530 4361
rect 15478 4297 15530 4303
rect 15298 3464 15422 3492
rect 15298 800 15326 3464
rect 15382 2949 15434 2955
rect 15382 2891 15434 2897
rect 15394 800 15422 2891
rect 15490 800 15518 4297
rect 15682 800 15710 7405
rect 15970 7099 15998 12215
rect 16066 8579 16094 12344
rect 16054 8573 16106 8579
rect 16054 8515 16106 8521
rect 16066 8431 16094 8515
rect 16054 8425 16106 8431
rect 16054 8367 16106 8373
rect 16054 8277 16106 8283
rect 16054 8219 16106 8225
rect 15958 7093 16010 7099
rect 15958 7035 16010 7041
rect 15958 6353 16010 6359
rect 15958 6295 16010 6301
rect 15970 5767 15998 6295
rect 15958 5761 16010 5767
rect 15958 5703 16010 5709
rect 15862 5687 15914 5693
rect 15862 5629 15914 5635
rect 15874 2900 15902 5629
rect 15958 4355 16010 4361
rect 15958 4297 16010 4303
rect 15778 2872 15902 2900
rect 15778 800 15806 2872
rect 15970 2160 15998 4297
rect 15874 2132 15998 2160
rect 15874 800 15902 2132
rect 16066 800 16094 8219
rect 16258 6433 16286 20355
rect 16354 9097 16382 23026
rect 16546 20863 16574 56393
rect 16630 56229 16682 56235
rect 16630 56171 16682 56177
rect 16534 20857 16586 20863
rect 16534 20799 16586 20805
rect 16342 9091 16394 9097
rect 16342 9033 16394 9039
rect 16342 8277 16394 8283
rect 16342 8219 16394 8225
rect 16246 6427 16298 6433
rect 16246 6369 16298 6375
rect 16150 5687 16202 5693
rect 16150 5629 16202 5635
rect 16162 800 16190 5629
rect 16246 4207 16298 4213
rect 16246 4149 16298 4155
rect 16258 800 16286 4149
rect 16354 800 16382 8219
rect 16642 7025 16670 56171
rect 16726 42243 16778 42249
rect 16726 42185 16778 42191
rect 16738 8875 16766 42185
rect 17590 27887 17642 27893
rect 17590 27829 17642 27835
rect 17398 26185 17450 26191
rect 17398 26127 17450 26133
rect 16822 25149 16874 25155
rect 16822 25091 16874 25097
rect 16726 8869 16778 8875
rect 16726 8811 16778 8817
rect 16834 8801 16862 25091
rect 17410 23054 17438 26127
rect 17410 23026 17534 23054
rect 17302 9609 17354 9615
rect 17302 9551 17354 9557
rect 16822 8795 16874 8801
rect 16822 8737 16874 8743
rect 16822 8351 16874 8357
rect 16822 8293 16874 8299
rect 16630 7019 16682 7025
rect 16630 6961 16682 6967
rect 16726 6131 16778 6137
rect 16726 6073 16778 6079
rect 16438 5021 16490 5027
rect 16438 4963 16490 4969
rect 16450 2955 16478 4963
rect 16534 3837 16586 3843
rect 16534 3779 16586 3785
rect 16438 2949 16490 2955
rect 16438 2891 16490 2897
rect 16546 800 16574 3779
rect 16630 3023 16682 3029
rect 16630 2965 16682 2971
rect 16642 800 16670 2965
rect 16738 800 16766 6073
rect 16834 2807 16862 8293
rect 17110 8203 17162 8209
rect 17110 8145 17162 8151
rect 17122 7617 17150 8145
rect 17110 7611 17162 7617
rect 17110 7553 17162 7559
rect 17110 7241 17162 7247
rect 17110 7183 17162 7189
rect 16918 4133 16970 4139
rect 16918 4075 16970 4081
rect 16822 2801 16874 2807
rect 16822 2743 16874 2749
rect 16930 800 16958 4075
rect 17014 3023 17066 3029
rect 17014 2965 17066 2971
rect 17026 800 17054 2965
rect 17122 800 17150 7183
rect 17314 7173 17342 9551
rect 17302 7167 17354 7173
rect 17302 7109 17354 7115
rect 17314 6951 17342 7109
rect 17302 6945 17354 6951
rect 17302 6887 17354 6893
rect 17302 5687 17354 5693
rect 17302 5629 17354 5635
rect 17314 3843 17342 5629
rect 17506 5120 17534 23026
rect 17602 5471 17630 27829
rect 17878 26111 17930 26117
rect 17878 26053 17930 26059
rect 17686 8795 17738 8801
rect 17686 8737 17738 8743
rect 17698 6433 17726 8737
rect 17890 7214 17918 26053
rect 17986 9467 18014 56837
rect 18082 56531 18110 59200
rect 18562 57614 18590 59200
rect 18562 57586 18782 57614
rect 18754 56531 18782 57586
rect 19138 56975 19166 59200
rect 19618 57614 19646 59200
rect 19522 57586 19646 57614
rect 19126 56969 19178 56975
rect 19126 56911 19178 56917
rect 19318 56895 19370 56901
rect 19318 56837 19370 56843
rect 18070 56525 18122 56531
rect 18070 56467 18122 56473
rect 18742 56525 18794 56531
rect 18742 56467 18794 56473
rect 18262 56229 18314 56235
rect 18262 56171 18314 56177
rect 18742 56229 18794 56235
rect 18742 56171 18794 56177
rect 18166 26777 18218 26783
rect 18166 26719 18218 26725
rect 17974 9461 18026 9467
rect 17974 9403 18026 9409
rect 18070 8869 18122 8875
rect 18070 8811 18122 8817
rect 17794 7186 17918 7214
rect 17974 7241 18026 7247
rect 17686 6427 17738 6433
rect 17686 6369 17738 6375
rect 17590 5465 17642 5471
rect 17590 5407 17642 5413
rect 17506 5092 17630 5120
rect 17494 5021 17546 5027
rect 17494 4963 17546 4969
rect 17302 3837 17354 3843
rect 17302 3779 17354 3785
rect 17398 3689 17450 3695
rect 17398 3631 17450 3637
rect 17302 3467 17354 3473
rect 17302 3409 17354 3415
rect 17314 2900 17342 3409
rect 17218 2872 17342 2900
rect 17218 800 17246 2872
rect 17410 800 17438 3631
rect 17506 3473 17534 4963
rect 17494 3467 17546 3473
rect 17494 3409 17546 3415
rect 17602 3251 17630 5092
rect 17686 4281 17738 4287
rect 17686 4223 17738 4229
rect 17590 3245 17642 3251
rect 17590 3187 17642 3193
rect 17494 3097 17546 3103
rect 17494 3039 17546 3045
rect 17506 800 17534 3039
rect 17698 3011 17726 4223
rect 17794 3177 17822 7186
rect 17974 7183 18026 7189
rect 17878 5465 17930 5471
rect 17878 5407 17930 5413
rect 17890 4139 17918 5407
rect 17878 4133 17930 4139
rect 17878 4075 17930 4081
rect 17986 3640 18014 7183
rect 18082 7099 18110 8811
rect 18070 7093 18122 7099
rect 18070 7035 18122 7041
rect 18070 6205 18122 6211
rect 18070 6147 18122 6153
rect 18082 3788 18110 6147
rect 18178 3917 18206 26719
rect 18274 14277 18302 56171
rect 18550 26555 18602 26561
rect 18550 26497 18602 26503
rect 18454 17453 18506 17459
rect 18454 17395 18506 17401
rect 18262 14271 18314 14277
rect 18262 14213 18314 14219
rect 18466 6433 18494 17395
rect 18454 6427 18506 6433
rect 18454 6369 18506 6375
rect 18358 6131 18410 6137
rect 18358 6073 18410 6079
rect 18262 5021 18314 5027
rect 18262 4963 18314 4969
rect 18166 3911 18218 3917
rect 18166 3853 18218 3859
rect 18082 3760 18206 3788
rect 17890 3612 18014 3640
rect 18070 3689 18122 3695
rect 18070 3631 18122 3637
rect 17782 3171 17834 3177
rect 17782 3113 17834 3119
rect 17602 2983 17726 3011
rect 17602 800 17630 2983
rect 17686 2949 17738 2955
rect 17686 2891 17738 2897
rect 17698 800 17726 2891
rect 17890 800 17918 3612
rect 17974 2949 18026 2955
rect 17974 2891 18026 2897
rect 17986 800 18014 2891
rect 18082 800 18110 3631
rect 18178 2752 18206 3760
rect 18274 2955 18302 4963
rect 18370 3103 18398 6073
rect 18562 3917 18590 26497
rect 18754 24267 18782 56171
rect 18838 40837 18890 40843
rect 18838 40779 18890 40785
rect 18742 24261 18794 24267
rect 18742 24203 18794 24209
rect 18646 7241 18698 7247
rect 18646 7183 18698 7189
rect 18550 3911 18602 3917
rect 18550 3853 18602 3859
rect 18454 3689 18506 3695
rect 18658 3640 18686 7183
rect 18850 6581 18878 40779
rect 18934 26481 18986 26487
rect 18934 26423 18986 26429
rect 18946 7099 18974 26423
rect 19330 9689 19358 56837
rect 19522 56161 19550 57586
rect 19628 56638 19924 56658
rect 19684 56636 19708 56638
rect 19764 56636 19788 56638
rect 19844 56636 19868 56638
rect 19706 56584 19708 56636
rect 19770 56584 19782 56636
rect 19844 56584 19846 56636
rect 19684 56582 19708 56584
rect 19764 56582 19788 56584
rect 19844 56582 19868 56584
rect 19628 56562 19924 56582
rect 19990 56229 20042 56235
rect 19990 56171 20042 56177
rect 19510 56155 19562 56161
rect 19510 56097 19562 56103
rect 19628 55306 19924 55326
rect 19684 55304 19708 55306
rect 19764 55304 19788 55306
rect 19844 55304 19868 55306
rect 19706 55252 19708 55304
rect 19770 55252 19782 55304
rect 19844 55252 19846 55304
rect 19684 55250 19708 55252
rect 19764 55250 19788 55252
rect 19844 55250 19868 55252
rect 19628 55230 19924 55250
rect 19628 53974 19924 53994
rect 19684 53972 19708 53974
rect 19764 53972 19788 53974
rect 19844 53972 19868 53974
rect 19706 53920 19708 53972
rect 19770 53920 19782 53972
rect 19844 53920 19846 53972
rect 19684 53918 19708 53920
rect 19764 53918 19788 53920
rect 19844 53918 19868 53920
rect 19628 53898 19924 53918
rect 19628 52642 19924 52662
rect 19684 52640 19708 52642
rect 19764 52640 19788 52642
rect 19844 52640 19868 52642
rect 19706 52588 19708 52640
rect 19770 52588 19782 52640
rect 19844 52588 19846 52640
rect 19684 52586 19708 52588
rect 19764 52586 19788 52588
rect 19844 52586 19868 52588
rect 19628 52566 19924 52586
rect 19628 51310 19924 51330
rect 19684 51308 19708 51310
rect 19764 51308 19788 51310
rect 19844 51308 19868 51310
rect 19706 51256 19708 51308
rect 19770 51256 19782 51308
rect 19844 51256 19846 51308
rect 19684 51254 19708 51256
rect 19764 51254 19788 51256
rect 19844 51254 19868 51256
rect 19628 51234 19924 51254
rect 19628 49978 19924 49998
rect 19684 49976 19708 49978
rect 19764 49976 19788 49978
rect 19844 49976 19868 49978
rect 19706 49924 19708 49976
rect 19770 49924 19782 49976
rect 19844 49924 19846 49976
rect 19684 49922 19708 49924
rect 19764 49922 19788 49924
rect 19844 49922 19868 49924
rect 19628 49902 19924 49922
rect 19628 48646 19924 48666
rect 19684 48644 19708 48646
rect 19764 48644 19788 48646
rect 19844 48644 19868 48646
rect 19706 48592 19708 48644
rect 19770 48592 19782 48644
rect 19844 48592 19846 48644
rect 19684 48590 19708 48592
rect 19764 48590 19788 48592
rect 19844 48590 19868 48592
rect 19628 48570 19924 48590
rect 19628 47314 19924 47334
rect 19684 47312 19708 47314
rect 19764 47312 19788 47314
rect 19844 47312 19868 47314
rect 19706 47260 19708 47312
rect 19770 47260 19782 47312
rect 19844 47260 19846 47312
rect 19684 47258 19708 47260
rect 19764 47258 19788 47260
rect 19844 47258 19868 47260
rect 19628 47238 19924 47258
rect 19628 45982 19924 46002
rect 19684 45980 19708 45982
rect 19764 45980 19788 45982
rect 19844 45980 19868 45982
rect 19706 45928 19708 45980
rect 19770 45928 19782 45980
rect 19844 45928 19846 45980
rect 19684 45926 19708 45928
rect 19764 45926 19788 45928
rect 19844 45926 19868 45928
rect 19628 45906 19924 45926
rect 19628 44650 19924 44670
rect 19684 44648 19708 44650
rect 19764 44648 19788 44650
rect 19844 44648 19868 44650
rect 19706 44596 19708 44648
rect 19770 44596 19782 44648
rect 19844 44596 19846 44648
rect 19684 44594 19708 44596
rect 19764 44594 19788 44596
rect 19844 44594 19868 44596
rect 19628 44574 19924 44594
rect 19628 43318 19924 43338
rect 19684 43316 19708 43318
rect 19764 43316 19788 43318
rect 19844 43316 19868 43318
rect 19706 43264 19708 43316
rect 19770 43264 19782 43316
rect 19844 43264 19846 43316
rect 19684 43262 19708 43264
rect 19764 43262 19788 43264
rect 19844 43262 19868 43264
rect 19628 43242 19924 43262
rect 19628 41986 19924 42006
rect 19684 41984 19708 41986
rect 19764 41984 19788 41986
rect 19844 41984 19868 41986
rect 19706 41932 19708 41984
rect 19770 41932 19782 41984
rect 19844 41932 19846 41984
rect 19684 41930 19708 41932
rect 19764 41930 19788 41932
rect 19844 41930 19868 41932
rect 19628 41910 19924 41930
rect 19628 40654 19924 40674
rect 19684 40652 19708 40654
rect 19764 40652 19788 40654
rect 19844 40652 19868 40654
rect 19706 40600 19708 40652
rect 19770 40600 19782 40652
rect 19844 40600 19846 40652
rect 19684 40598 19708 40600
rect 19764 40598 19788 40600
rect 19844 40598 19868 40600
rect 19628 40578 19924 40598
rect 19628 39322 19924 39342
rect 19684 39320 19708 39322
rect 19764 39320 19788 39322
rect 19844 39320 19868 39322
rect 19706 39268 19708 39320
rect 19770 39268 19782 39320
rect 19844 39268 19846 39320
rect 19684 39266 19708 39268
rect 19764 39266 19788 39268
rect 19844 39266 19868 39268
rect 19628 39246 19924 39266
rect 19628 37990 19924 38010
rect 19684 37988 19708 37990
rect 19764 37988 19788 37990
rect 19844 37988 19868 37990
rect 19706 37936 19708 37988
rect 19770 37936 19782 37988
rect 19844 37936 19846 37988
rect 19684 37934 19708 37936
rect 19764 37934 19788 37936
rect 19844 37934 19868 37936
rect 19628 37914 19924 37934
rect 19628 36658 19924 36678
rect 19684 36656 19708 36658
rect 19764 36656 19788 36658
rect 19844 36656 19868 36658
rect 19706 36604 19708 36656
rect 19770 36604 19782 36656
rect 19844 36604 19846 36656
rect 19684 36602 19708 36604
rect 19764 36602 19788 36604
rect 19844 36602 19868 36604
rect 19628 36582 19924 36602
rect 19628 35326 19924 35346
rect 19684 35324 19708 35326
rect 19764 35324 19788 35326
rect 19844 35324 19868 35326
rect 19706 35272 19708 35324
rect 19770 35272 19782 35324
rect 19844 35272 19846 35324
rect 19684 35270 19708 35272
rect 19764 35270 19788 35272
rect 19844 35270 19868 35272
rect 19628 35250 19924 35270
rect 19628 33994 19924 34014
rect 19684 33992 19708 33994
rect 19764 33992 19788 33994
rect 19844 33992 19868 33994
rect 19706 33940 19708 33992
rect 19770 33940 19782 33992
rect 19844 33940 19846 33992
rect 19684 33938 19708 33940
rect 19764 33938 19788 33940
rect 19844 33938 19868 33940
rect 19628 33918 19924 33938
rect 19628 32662 19924 32682
rect 19684 32660 19708 32662
rect 19764 32660 19788 32662
rect 19844 32660 19868 32662
rect 19706 32608 19708 32660
rect 19770 32608 19782 32660
rect 19844 32608 19846 32660
rect 19684 32606 19708 32608
rect 19764 32606 19788 32608
rect 19844 32606 19868 32608
rect 19628 32586 19924 32606
rect 19628 31330 19924 31350
rect 19684 31328 19708 31330
rect 19764 31328 19788 31330
rect 19844 31328 19868 31330
rect 19706 31276 19708 31328
rect 19770 31276 19782 31328
rect 19844 31276 19846 31328
rect 19684 31274 19708 31276
rect 19764 31274 19788 31276
rect 19844 31274 19868 31276
rect 19628 31254 19924 31274
rect 19628 29998 19924 30018
rect 19684 29996 19708 29998
rect 19764 29996 19788 29998
rect 19844 29996 19868 29998
rect 19706 29944 19708 29996
rect 19770 29944 19782 29996
rect 19844 29944 19846 29996
rect 19684 29942 19708 29944
rect 19764 29942 19788 29944
rect 19844 29942 19868 29944
rect 19628 29922 19924 29942
rect 19628 28666 19924 28686
rect 19684 28664 19708 28666
rect 19764 28664 19788 28666
rect 19844 28664 19868 28666
rect 19706 28612 19708 28664
rect 19770 28612 19782 28664
rect 19844 28612 19846 28664
rect 19684 28610 19708 28612
rect 19764 28610 19788 28612
rect 19844 28610 19868 28612
rect 19628 28590 19924 28610
rect 19628 27334 19924 27354
rect 19684 27332 19708 27334
rect 19764 27332 19788 27334
rect 19844 27332 19868 27334
rect 19706 27280 19708 27332
rect 19770 27280 19782 27332
rect 19844 27280 19846 27332
rect 19684 27278 19708 27280
rect 19764 27278 19788 27280
rect 19844 27278 19868 27280
rect 19628 27258 19924 27278
rect 19628 26002 19924 26022
rect 19684 26000 19708 26002
rect 19764 26000 19788 26002
rect 19844 26000 19868 26002
rect 19706 25948 19708 26000
rect 19770 25948 19782 26000
rect 19844 25948 19846 26000
rect 19684 25946 19708 25948
rect 19764 25946 19788 25948
rect 19844 25946 19868 25948
rect 19628 25926 19924 25946
rect 19628 24670 19924 24690
rect 19684 24668 19708 24670
rect 19764 24668 19788 24670
rect 19844 24668 19868 24670
rect 19706 24616 19708 24668
rect 19770 24616 19782 24668
rect 19844 24616 19846 24668
rect 19684 24614 19708 24616
rect 19764 24614 19788 24616
rect 19844 24614 19868 24616
rect 19628 24594 19924 24614
rect 19628 23338 19924 23358
rect 19684 23336 19708 23338
rect 19764 23336 19788 23338
rect 19844 23336 19868 23338
rect 19706 23284 19708 23336
rect 19770 23284 19782 23336
rect 19844 23284 19846 23336
rect 19684 23282 19708 23284
rect 19764 23282 19788 23284
rect 19844 23282 19868 23284
rect 19628 23262 19924 23282
rect 19628 22006 19924 22026
rect 19684 22004 19708 22006
rect 19764 22004 19788 22006
rect 19844 22004 19868 22006
rect 19706 21952 19708 22004
rect 19770 21952 19782 22004
rect 19844 21952 19846 22004
rect 19684 21950 19708 21952
rect 19764 21950 19788 21952
rect 19844 21950 19868 21952
rect 19628 21930 19924 21950
rect 19628 20674 19924 20694
rect 19684 20672 19708 20674
rect 19764 20672 19788 20674
rect 19844 20672 19868 20674
rect 19706 20620 19708 20672
rect 19770 20620 19782 20672
rect 19844 20620 19846 20672
rect 19684 20618 19708 20620
rect 19764 20618 19788 20620
rect 19844 20618 19868 20620
rect 19628 20598 19924 20618
rect 19628 19342 19924 19362
rect 19684 19340 19708 19342
rect 19764 19340 19788 19342
rect 19844 19340 19868 19342
rect 19706 19288 19708 19340
rect 19770 19288 19782 19340
rect 19844 19288 19846 19340
rect 19684 19286 19708 19288
rect 19764 19286 19788 19288
rect 19844 19286 19868 19288
rect 19628 19266 19924 19286
rect 20002 18199 20030 56171
rect 20194 55717 20222 59200
rect 20674 56975 20702 59200
rect 20662 56969 20714 56975
rect 20662 56911 20714 56917
rect 20854 56895 20906 56901
rect 20854 56837 20906 56843
rect 20182 55711 20234 55717
rect 20182 55653 20234 55659
rect 20470 55563 20522 55569
rect 20470 55505 20522 55511
rect 20086 42761 20138 42767
rect 20086 42703 20138 42709
rect 19990 18193 20042 18199
rect 19990 18135 20042 18141
rect 19628 18010 19924 18030
rect 19684 18008 19708 18010
rect 19764 18008 19788 18010
rect 19844 18008 19868 18010
rect 19706 17956 19708 18008
rect 19770 17956 19782 18008
rect 19844 17956 19846 18008
rect 19684 17954 19708 17956
rect 19764 17954 19788 17956
rect 19844 17954 19868 17956
rect 19628 17934 19924 17954
rect 19628 16678 19924 16698
rect 19684 16676 19708 16678
rect 19764 16676 19788 16678
rect 19844 16676 19868 16678
rect 19706 16624 19708 16676
rect 19770 16624 19782 16676
rect 19844 16624 19846 16676
rect 19684 16622 19708 16624
rect 19764 16622 19788 16624
rect 19844 16622 19868 16624
rect 19628 16602 19924 16622
rect 19628 15346 19924 15366
rect 19684 15344 19708 15346
rect 19764 15344 19788 15346
rect 19844 15344 19868 15346
rect 19706 15292 19708 15344
rect 19770 15292 19782 15344
rect 19844 15292 19846 15344
rect 19684 15290 19708 15292
rect 19764 15290 19788 15292
rect 19844 15290 19868 15292
rect 19628 15270 19924 15290
rect 19628 14014 19924 14034
rect 19684 14012 19708 14014
rect 19764 14012 19788 14014
rect 19844 14012 19868 14014
rect 19706 13960 19708 14012
rect 19770 13960 19782 14012
rect 19844 13960 19846 14012
rect 19684 13958 19708 13960
rect 19764 13958 19788 13960
rect 19844 13958 19868 13960
rect 19628 13938 19924 13958
rect 19628 12682 19924 12702
rect 19684 12680 19708 12682
rect 19764 12680 19788 12682
rect 19844 12680 19868 12682
rect 19706 12628 19708 12680
rect 19770 12628 19782 12680
rect 19844 12628 19846 12680
rect 19684 12626 19708 12628
rect 19764 12626 19788 12628
rect 19844 12626 19868 12628
rect 19628 12606 19924 12626
rect 19628 11350 19924 11370
rect 19684 11348 19708 11350
rect 19764 11348 19788 11350
rect 19844 11348 19868 11350
rect 19706 11296 19708 11348
rect 19770 11296 19782 11348
rect 19844 11296 19846 11348
rect 19684 11294 19708 11296
rect 19764 11294 19788 11296
rect 19844 11294 19868 11296
rect 19628 11274 19924 11294
rect 19628 10018 19924 10038
rect 19684 10016 19708 10018
rect 19764 10016 19788 10018
rect 19844 10016 19868 10018
rect 19706 9964 19708 10016
rect 19770 9964 19782 10016
rect 19844 9964 19846 10016
rect 19684 9962 19708 9964
rect 19764 9962 19788 9964
rect 19844 9962 19868 9964
rect 19628 9942 19924 9962
rect 19318 9683 19370 9689
rect 19318 9625 19370 9631
rect 19628 8686 19924 8706
rect 19684 8684 19708 8686
rect 19764 8684 19788 8686
rect 19844 8684 19868 8686
rect 19706 8632 19708 8684
rect 19770 8632 19782 8684
rect 19844 8632 19846 8684
rect 19684 8630 19708 8632
rect 19764 8630 19788 8632
rect 19844 8630 19868 8632
rect 19628 8610 19924 8630
rect 20098 8431 20126 42703
rect 20482 38253 20510 55505
rect 20566 55045 20618 55051
rect 20566 54987 20618 54993
rect 20470 38247 20522 38253
rect 20470 38189 20522 38195
rect 20374 27443 20426 27449
rect 20374 27385 20426 27391
rect 20086 8425 20138 8431
rect 20086 8367 20138 8373
rect 19628 7354 19924 7374
rect 19684 7352 19708 7354
rect 19764 7352 19788 7354
rect 19844 7352 19868 7354
rect 19706 7300 19708 7352
rect 19770 7300 19782 7352
rect 19844 7300 19846 7352
rect 19684 7298 19708 7300
rect 19764 7298 19788 7300
rect 19844 7298 19868 7300
rect 19628 7278 19924 7298
rect 20386 7099 20414 27385
rect 18934 7093 18986 7099
rect 18934 7035 18986 7041
rect 20374 7093 20426 7099
rect 20374 7035 20426 7041
rect 19510 6945 19562 6951
rect 19510 6887 19562 6893
rect 20374 6945 20426 6951
rect 20374 6887 20426 6893
rect 18838 6575 18890 6581
rect 18838 6517 18890 6523
rect 18850 6433 18878 6517
rect 18838 6427 18890 6433
rect 18838 6369 18890 6375
rect 19318 6279 19370 6285
rect 19318 6221 19370 6227
rect 18934 6205 18986 6211
rect 18934 6147 18986 6153
rect 18742 5687 18794 5693
rect 18742 5629 18794 5635
rect 18454 3631 18506 3637
rect 18358 3097 18410 3103
rect 18358 3039 18410 3045
rect 18262 2949 18314 2955
rect 18262 2891 18314 2897
rect 18358 2949 18410 2955
rect 18358 2891 18410 2897
rect 18178 2724 18302 2752
rect 18274 800 18302 2724
rect 18370 800 18398 2891
rect 18466 800 18494 3631
rect 18562 3612 18686 3640
rect 18562 800 18590 3612
rect 18754 800 18782 5629
rect 18838 3023 18890 3029
rect 18838 2965 18890 2971
rect 18850 800 18878 2965
rect 18946 800 18974 6147
rect 19030 5021 19082 5027
rect 19030 4963 19082 4969
rect 19126 5021 19178 5027
rect 19126 4963 19178 4969
rect 19042 2955 19070 4963
rect 19030 2949 19082 2955
rect 19030 2891 19082 2897
rect 19138 2604 19166 4963
rect 19222 3689 19274 3695
rect 19222 3631 19274 3637
rect 19042 2576 19166 2604
rect 19042 800 19070 2576
rect 19234 800 19262 3631
rect 19330 800 19358 6221
rect 19414 3837 19466 3843
rect 19414 3779 19466 3785
rect 19426 800 19454 3779
rect 19522 3196 19550 6887
rect 20086 6353 20138 6359
rect 20086 6295 20138 6301
rect 19628 6022 19924 6042
rect 19684 6020 19708 6022
rect 19764 6020 19788 6022
rect 19844 6020 19868 6022
rect 19706 5968 19708 6020
rect 19770 5968 19782 6020
rect 19844 5968 19846 6020
rect 19684 5966 19708 5968
rect 19764 5966 19788 5968
rect 19844 5966 19868 5968
rect 19628 5946 19924 5966
rect 19628 4690 19924 4710
rect 19684 4688 19708 4690
rect 19764 4688 19788 4690
rect 19844 4688 19868 4690
rect 19706 4636 19708 4688
rect 19770 4636 19782 4688
rect 19844 4636 19846 4688
rect 19684 4634 19708 4636
rect 19764 4634 19788 4636
rect 19844 4634 19868 4636
rect 19628 4614 19924 4634
rect 19990 3615 20042 3621
rect 19990 3557 20042 3563
rect 19628 3358 19924 3378
rect 19684 3356 19708 3358
rect 19764 3356 19788 3358
rect 19844 3356 19868 3358
rect 19706 3304 19708 3356
rect 19770 3304 19782 3356
rect 19844 3304 19846 3356
rect 19684 3302 19708 3304
rect 19764 3302 19788 3304
rect 19844 3302 19868 3304
rect 19628 3282 19924 3302
rect 19522 3168 19742 3196
rect 19606 3097 19658 3103
rect 19606 3039 19658 3045
rect 19618 800 19646 3039
rect 19714 800 19742 3168
rect 19798 3171 19850 3177
rect 19798 3113 19850 3119
rect 19810 800 19838 3113
rect 20002 1864 20030 3557
rect 19906 1836 20030 1864
rect 19906 800 19934 1836
rect 20098 800 20126 6295
rect 20182 5687 20234 5693
rect 20182 5629 20234 5635
rect 20194 3177 20222 5629
rect 20278 4355 20330 4361
rect 20278 4297 20330 4303
rect 20182 3171 20234 3177
rect 20182 3113 20234 3119
rect 20182 2431 20234 2437
rect 20182 2373 20234 2379
rect 20194 800 20222 2373
rect 20290 800 20318 4297
rect 20386 3492 20414 6887
rect 20578 6581 20606 54987
rect 20866 9763 20894 56837
rect 21250 56531 21278 59200
rect 21730 56531 21758 59200
rect 22306 56975 22334 59200
rect 22294 56969 22346 56975
rect 22294 56911 22346 56917
rect 22786 56531 22814 59200
rect 21238 56525 21290 56531
rect 21238 56467 21290 56473
rect 21718 56525 21770 56531
rect 21718 56467 21770 56473
rect 22774 56525 22826 56531
rect 22774 56467 22826 56473
rect 21046 56229 21098 56235
rect 21046 56171 21098 56177
rect 21814 56229 21866 56235
rect 21814 56171 21866 56177
rect 22966 56229 23018 56235
rect 22966 56171 23018 56177
rect 20950 29145 21002 29151
rect 20950 29087 21002 29093
rect 20854 9757 20906 9763
rect 20854 9699 20906 9705
rect 20962 7765 20990 29087
rect 21058 18939 21086 56171
rect 21142 42761 21194 42767
rect 21142 42703 21194 42709
rect 21046 18933 21098 18939
rect 21046 18875 21098 18881
rect 20950 7759 21002 7765
rect 20950 7701 21002 7707
rect 20758 7463 20810 7469
rect 20758 7405 20810 7411
rect 20566 6575 20618 6581
rect 20566 6517 20618 6523
rect 20578 6433 20606 6517
rect 20566 6427 20618 6433
rect 20566 6369 20618 6375
rect 20566 5687 20618 5693
rect 20566 5629 20618 5635
rect 20470 5169 20522 5175
rect 20470 5111 20522 5117
rect 20482 4583 20510 5111
rect 20470 4577 20522 4583
rect 20470 4519 20522 4525
rect 20386 3464 20510 3492
rect 20482 800 20510 3464
rect 20578 800 20606 5629
rect 20662 5021 20714 5027
rect 20662 4963 20714 4969
rect 20674 3843 20702 4963
rect 20662 3837 20714 3843
rect 20662 3779 20714 3785
rect 20662 3689 20714 3695
rect 20662 3631 20714 3637
rect 20674 800 20702 3631
rect 20770 800 20798 7405
rect 21154 7099 21182 42703
rect 21826 13907 21854 56171
rect 22978 38771 23006 56171
rect 23362 55717 23390 59200
rect 23842 56975 23870 59200
rect 23830 56969 23882 56975
rect 23830 56911 23882 56917
rect 24022 56895 24074 56901
rect 24022 56837 24074 56843
rect 23350 55711 23402 55717
rect 23350 55653 23402 55659
rect 23446 55563 23498 55569
rect 23446 55505 23498 55511
rect 23062 51567 23114 51573
rect 23062 51509 23114 51515
rect 22966 38765 23018 38771
rect 22966 38707 23018 38713
rect 22582 32771 22634 32777
rect 22582 32713 22634 32719
rect 21910 18859 21962 18865
rect 21910 18801 21962 18807
rect 21814 13901 21866 13907
rect 21814 13843 21866 13849
rect 21922 7099 21950 18801
rect 21142 7093 21194 7099
rect 21142 7035 21194 7041
rect 21910 7093 21962 7099
rect 21910 7035 21962 7041
rect 21142 6945 21194 6951
rect 21142 6887 21194 6893
rect 21910 6945 21962 6951
rect 21910 6887 21962 6893
rect 20854 5021 20906 5027
rect 20854 4963 20906 4969
rect 20866 2437 20894 4963
rect 21046 4355 21098 4361
rect 21046 4297 21098 4303
rect 20950 4133 21002 4139
rect 20950 4075 21002 4081
rect 20962 3251 20990 4075
rect 20950 3245 21002 3251
rect 20950 3187 21002 3193
rect 20950 3097 21002 3103
rect 20950 3039 21002 3045
rect 20854 2431 20906 2437
rect 20854 2373 20906 2379
rect 20962 800 20990 3039
rect 21058 800 21086 4297
rect 21154 800 21182 6887
rect 21622 5761 21674 5767
rect 21622 5703 21674 5709
rect 21526 4133 21578 4139
rect 21526 4075 21578 4081
rect 21238 3911 21290 3917
rect 21238 3853 21290 3859
rect 21250 800 21278 3853
rect 21430 3023 21482 3029
rect 21430 2965 21482 2971
rect 21442 800 21470 2965
rect 21538 800 21566 4075
rect 21634 800 21662 5703
rect 21718 5687 21770 5693
rect 21718 5629 21770 5635
rect 21730 3103 21758 5629
rect 21814 4355 21866 4361
rect 21814 4297 21866 4303
rect 21718 3097 21770 3103
rect 21718 3039 21770 3045
rect 21826 800 21854 4297
rect 21922 800 21950 6887
rect 22594 6581 22622 32713
rect 22966 27591 23018 27597
rect 22966 27533 23018 27539
rect 22678 23891 22730 23897
rect 22678 23833 22730 23839
rect 22690 7099 22718 23833
rect 22978 9097 23006 27533
rect 22966 9091 23018 9097
rect 22966 9033 23018 9039
rect 23074 7173 23102 51509
rect 23350 40097 23402 40103
rect 23350 40039 23402 40045
rect 23062 7167 23114 7173
rect 23062 7109 23114 7115
rect 23362 7099 23390 40039
rect 23458 9911 23486 55505
rect 23542 52751 23594 52757
rect 23542 52693 23594 52699
rect 23446 9905 23498 9911
rect 23446 9847 23498 9853
rect 23554 8357 23582 52693
rect 23926 43501 23978 43507
rect 23926 43443 23978 43449
rect 23734 37063 23786 37069
rect 23734 37005 23786 37011
rect 23542 8351 23594 8357
rect 23542 8293 23594 8299
rect 22678 7093 22730 7099
rect 22678 7035 22730 7041
rect 23350 7093 23402 7099
rect 23350 7035 23402 7041
rect 22678 6945 22730 6951
rect 23446 6945 23498 6951
rect 22678 6887 22730 6893
rect 23362 6905 23446 6933
rect 22582 6575 22634 6581
rect 22582 6517 22634 6523
rect 22594 6433 22622 6517
rect 22582 6427 22634 6433
rect 22582 6369 22634 6375
rect 22294 6205 22346 6211
rect 22294 6147 22346 6153
rect 22006 4281 22058 4287
rect 22006 4223 22058 4229
rect 22018 800 22046 4223
rect 22102 3689 22154 3695
rect 22102 3631 22154 3637
rect 22114 800 22142 3631
rect 22306 800 22334 6147
rect 22690 3492 22718 6887
rect 22966 6279 23018 6285
rect 22966 6221 23018 6227
rect 22870 6131 22922 6137
rect 22870 6073 22922 6079
rect 22774 5021 22826 5027
rect 22774 4963 22826 4969
rect 22786 3917 22814 4963
rect 22882 4139 22910 6073
rect 22870 4133 22922 4139
rect 22870 4075 22922 4081
rect 22774 3911 22826 3917
rect 22774 3853 22826 3859
rect 22870 3689 22922 3695
rect 22870 3631 22922 3637
rect 22594 3464 22718 3492
rect 22390 3171 22442 3177
rect 22390 3113 22442 3119
rect 22402 800 22430 3113
rect 22486 3097 22538 3103
rect 22486 3039 22538 3045
rect 22498 800 22526 3039
rect 22594 800 22622 3464
rect 22774 3245 22826 3251
rect 22774 3187 22826 3193
rect 22786 800 22814 3187
rect 22882 800 22910 3631
rect 22978 800 23006 6221
rect 23158 5687 23210 5693
rect 23158 5629 23210 5635
rect 23062 4947 23114 4953
rect 23062 4889 23114 4895
rect 23074 2894 23102 4889
rect 23170 3251 23198 5629
rect 23254 4355 23306 4361
rect 23254 4297 23306 4303
rect 23158 3245 23210 3251
rect 23158 3187 23210 3193
rect 23074 2866 23198 2894
rect 23170 800 23198 2866
rect 23266 800 23294 4297
rect 23362 800 23390 6905
rect 23446 6887 23498 6893
rect 23746 6433 23774 37005
rect 23938 7765 23966 43443
rect 24034 11021 24062 56837
rect 24418 56531 24446 59200
rect 24406 56525 24458 56531
rect 24406 56467 24458 56473
rect 24310 56229 24362 56235
rect 24310 56171 24362 56177
rect 24118 36101 24170 36107
rect 24118 36043 24170 36049
rect 24022 11015 24074 11021
rect 24022 10957 24074 10963
rect 23926 7759 23978 7765
rect 23926 7701 23978 7707
rect 23830 7463 23882 7469
rect 23830 7405 23882 7411
rect 23734 6427 23786 6433
rect 23734 6369 23786 6375
rect 23446 5687 23498 5693
rect 23446 5629 23498 5635
rect 23458 800 23486 5629
rect 23542 5021 23594 5027
rect 23542 4963 23594 4969
rect 23554 3177 23582 4963
rect 23638 3689 23690 3695
rect 23638 3631 23690 3637
rect 23542 3171 23594 3177
rect 23542 3113 23594 3119
rect 23650 800 23678 3631
rect 23842 1568 23870 7405
rect 24130 6581 24158 36043
rect 24322 29225 24350 56171
rect 24898 55717 24926 59200
rect 25474 56975 25502 59200
rect 25462 56969 25514 56975
rect 25462 56911 25514 56917
rect 25954 56531 25982 59200
rect 26530 56531 26558 59200
rect 27010 56975 27038 59200
rect 26998 56969 27050 56975
rect 26998 56911 27050 56917
rect 27190 56895 27242 56901
rect 27190 56837 27242 56843
rect 26710 56821 26762 56827
rect 26710 56763 26762 56769
rect 25942 56525 25994 56531
rect 25942 56467 25994 56473
rect 26518 56525 26570 56531
rect 26518 56467 26570 56473
rect 26422 56303 26474 56309
rect 26422 56245 26474 56251
rect 26326 55785 26378 55791
rect 26326 55727 26378 55733
rect 24886 55711 24938 55717
rect 24886 55653 24938 55659
rect 24694 55415 24746 55421
rect 24694 55357 24746 55363
rect 24706 55199 24734 55357
rect 24694 55193 24746 55199
rect 24694 55135 24746 55141
rect 26134 53491 26186 53497
rect 26134 53433 26186 53439
rect 25078 52899 25130 52905
rect 25078 52841 25130 52847
rect 24310 29219 24362 29225
rect 24310 29161 24362 29167
rect 24694 10349 24746 10355
rect 24694 10291 24746 10297
rect 24310 9535 24362 9541
rect 24310 9477 24362 9483
rect 24214 7463 24266 7469
rect 24214 7405 24266 7411
rect 24118 6575 24170 6581
rect 24118 6517 24170 6523
rect 24130 6433 24158 6517
rect 24118 6427 24170 6433
rect 24118 6369 24170 6375
rect 24226 5120 24254 7405
rect 24322 7099 24350 9477
rect 24706 7765 24734 10291
rect 25090 7839 25118 52841
rect 25462 18785 25514 18791
rect 25462 18727 25514 18733
rect 25366 9461 25418 9467
rect 25366 9403 25418 9409
rect 25078 7833 25130 7839
rect 25078 7775 25130 7781
rect 24694 7759 24746 7765
rect 24694 7701 24746 7707
rect 24790 7463 24842 7469
rect 24790 7405 24842 7411
rect 24310 7093 24362 7099
rect 24310 7035 24362 7041
rect 24502 6945 24554 6951
rect 24502 6887 24554 6893
rect 24130 5092 24254 5120
rect 23926 3911 23978 3917
rect 23926 3853 23978 3859
rect 23746 1540 23870 1568
rect 23746 800 23774 1540
rect 23938 1420 23966 3853
rect 24022 3023 24074 3029
rect 24022 2965 24074 2971
rect 23842 1392 23966 1420
rect 23842 800 23870 1392
rect 24034 800 24062 2965
rect 24130 800 24158 5092
rect 24214 3837 24266 3843
rect 24214 3779 24266 3785
rect 24226 800 24254 3779
rect 24406 3689 24458 3695
rect 24406 3631 24458 3637
rect 24418 1864 24446 3631
rect 24322 1836 24446 1864
rect 24322 800 24350 1836
rect 24514 800 24542 6887
rect 24598 5687 24650 5693
rect 24598 5629 24650 5635
rect 24610 800 24638 5629
rect 24694 3615 24746 3621
rect 24694 3557 24746 3563
rect 24706 800 24734 3557
rect 24802 800 24830 7405
rect 25174 7019 25226 7025
rect 25174 6961 25226 6967
rect 25078 5021 25130 5027
rect 25078 4963 25130 4969
rect 24982 4133 25034 4139
rect 24982 4075 25034 4081
rect 24994 800 25022 4075
rect 25090 3917 25118 4963
rect 25078 3911 25130 3917
rect 25078 3853 25130 3859
rect 25078 3097 25130 3103
rect 25078 3039 25130 3045
rect 25090 800 25118 3039
rect 25186 800 25214 6961
rect 25378 6359 25406 9403
rect 25474 7099 25502 18727
rect 25654 10423 25706 10429
rect 25654 10365 25706 10371
rect 25666 8431 25694 10365
rect 25654 8425 25706 8431
rect 25654 8367 25706 8373
rect 26146 7765 26174 53433
rect 26134 7759 26186 7765
rect 26134 7701 26186 7707
rect 25558 7463 25610 7469
rect 25558 7405 25610 7411
rect 25462 7093 25514 7099
rect 25462 7035 25514 7041
rect 25366 6353 25418 6359
rect 25366 6295 25418 6301
rect 25462 4355 25514 4361
rect 25462 4297 25514 4303
rect 25366 3171 25418 3177
rect 25366 3113 25418 3119
rect 25378 800 25406 3113
rect 25474 800 25502 4297
rect 25570 800 25598 7405
rect 26338 7099 26366 55727
rect 26434 21085 26462 56245
rect 26518 56229 26570 56235
rect 26518 56171 26570 56177
rect 26422 21079 26474 21085
rect 26422 21021 26474 21027
rect 26530 10133 26558 56171
rect 26722 55199 26750 56763
rect 26710 55193 26762 55199
rect 26710 55135 26762 55141
rect 26998 34399 27050 34405
rect 26998 34341 27050 34347
rect 26806 16195 26858 16201
rect 26806 16137 26858 16143
rect 26818 15905 26846 16137
rect 26806 15899 26858 15905
rect 26806 15841 26858 15847
rect 26518 10127 26570 10133
rect 26518 10069 26570 10075
rect 27010 7765 27038 34341
rect 27202 11243 27230 56837
rect 27586 56531 27614 59200
rect 28066 56531 28094 59200
rect 28642 56975 28670 59200
rect 29122 57049 29150 59200
rect 29110 57043 29162 57049
rect 29110 56985 29162 56991
rect 28630 56969 28682 56975
rect 28630 56911 28682 56917
rect 28822 56895 28874 56901
rect 28822 56837 28874 56843
rect 27574 56525 27626 56531
rect 27574 56467 27626 56473
rect 28054 56525 28106 56531
rect 28054 56467 28106 56473
rect 27670 56229 27722 56235
rect 27670 56171 27722 56177
rect 28150 56229 28202 56235
rect 28150 56171 28202 56177
rect 27286 49125 27338 49131
rect 27286 49067 27338 49073
rect 27190 11237 27242 11243
rect 27190 11179 27242 11185
rect 26998 7759 27050 7765
rect 26998 7701 27050 7707
rect 26710 7463 26762 7469
rect 26710 7405 26762 7411
rect 26326 7093 26378 7099
rect 26326 7035 26378 7041
rect 25942 7019 25994 7025
rect 25942 6961 25994 6967
rect 25654 6353 25706 6359
rect 25654 6295 25706 6301
rect 25666 800 25694 6295
rect 25846 5021 25898 5027
rect 25846 4963 25898 4969
rect 25858 3843 25886 4963
rect 25846 3837 25898 3843
rect 25846 3779 25898 3785
rect 25846 3541 25898 3547
rect 25846 3483 25898 3489
rect 25858 800 25886 3483
rect 25954 800 25982 6961
rect 26326 6131 26378 6137
rect 26326 6073 26378 6079
rect 26038 5761 26090 5767
rect 26038 5703 26090 5709
rect 26050 800 26078 5703
rect 26230 5687 26282 5693
rect 26230 5629 26282 5635
rect 26134 4355 26186 4361
rect 26134 4297 26186 4303
rect 26146 800 26174 4297
rect 26242 3177 26270 5629
rect 26230 3171 26282 3177
rect 26230 3113 26282 3119
rect 26338 800 26366 6073
rect 26614 5021 26666 5027
rect 26614 4963 26666 4969
rect 26518 4355 26570 4361
rect 26518 4297 26570 4303
rect 26422 3837 26474 3843
rect 26422 3779 26474 3785
rect 26434 800 26462 3779
rect 26530 800 26558 4297
rect 26626 4139 26654 4963
rect 26614 4133 26666 4139
rect 26614 4075 26666 4081
rect 26722 800 26750 7405
rect 27298 7099 27326 49067
rect 27682 14869 27710 56171
rect 27766 42539 27818 42545
rect 27766 42481 27818 42487
rect 27670 14863 27722 14869
rect 27670 14805 27722 14811
rect 27778 7839 27806 42481
rect 27862 33437 27914 33443
rect 27862 33379 27914 33385
rect 27766 7833 27818 7839
rect 27766 7775 27818 7781
rect 27286 7093 27338 7099
rect 27286 7035 27338 7041
rect 26998 7019 27050 7025
rect 26998 6961 27050 6967
rect 26806 6353 26858 6359
rect 26806 6295 26858 6301
rect 26818 800 26846 6295
rect 26902 3023 26954 3029
rect 26902 2965 26954 2971
rect 26914 800 26942 2965
rect 27010 800 27038 6961
rect 27874 6581 27902 33379
rect 28162 29521 28190 56171
rect 28630 55415 28682 55421
rect 28630 55357 28682 55363
rect 28642 54977 28670 55357
rect 28630 54971 28682 54977
rect 28630 54913 28682 54919
rect 28342 47571 28394 47577
rect 28342 47513 28394 47519
rect 28246 36915 28298 36921
rect 28246 36857 28298 36863
rect 28258 36551 28286 36857
rect 28246 36545 28298 36551
rect 28246 36487 28298 36493
rect 28150 29515 28202 29521
rect 28150 29457 28202 29463
rect 27958 14789 28010 14795
rect 27958 14731 28010 14737
rect 27970 7099 27998 14731
rect 28054 8129 28106 8135
rect 28054 8071 28106 8077
rect 28066 7913 28094 8071
rect 28054 7907 28106 7913
rect 28054 7849 28106 7855
rect 28150 7463 28202 7469
rect 28150 7405 28202 7411
rect 27958 7093 28010 7099
rect 27958 7035 28010 7041
rect 27958 6945 28010 6951
rect 27958 6887 28010 6893
rect 27862 6575 27914 6581
rect 27862 6517 27914 6523
rect 27874 6433 27902 6517
rect 27862 6427 27914 6433
rect 27862 6369 27914 6375
rect 27478 6205 27530 6211
rect 27478 6147 27530 6153
rect 27382 5687 27434 5693
rect 27382 5629 27434 5635
rect 27394 4232 27422 5629
rect 27202 4204 27422 4232
rect 27202 800 27230 4204
rect 27490 4121 27518 6147
rect 27862 5687 27914 5693
rect 27862 5629 27914 5635
rect 27394 4093 27518 4121
rect 27286 3689 27338 3695
rect 27286 3631 27338 3637
rect 27298 800 27326 3631
rect 27394 800 27422 4093
rect 27478 3911 27530 3917
rect 27478 3853 27530 3859
rect 27490 800 27518 3853
rect 27670 3097 27722 3103
rect 27670 3039 27722 3045
rect 27682 800 27710 3039
rect 27766 2801 27818 2807
rect 27766 2743 27818 2749
rect 27778 800 27806 2743
rect 27874 800 27902 5629
rect 27970 2807 27998 6887
rect 28054 5021 28106 5027
rect 28054 4963 28106 4969
rect 28066 3843 28094 4963
rect 28054 3837 28106 3843
rect 28054 3779 28106 3785
rect 28054 3541 28106 3547
rect 28054 3483 28106 3489
rect 27958 2801 28010 2807
rect 27958 2743 28010 2749
rect 28066 800 28094 3483
rect 28162 800 28190 7405
rect 28354 7173 28382 47513
rect 28834 12131 28862 56837
rect 29698 56531 29726 59200
rect 30178 56975 30206 59200
rect 30166 56969 30218 56975
rect 30166 56911 30218 56917
rect 30658 56531 30686 59200
rect 29686 56525 29738 56531
rect 29686 56467 29738 56473
rect 30646 56525 30698 56531
rect 30646 56467 30698 56473
rect 29590 56229 29642 56235
rect 29590 56171 29642 56177
rect 30934 56229 30986 56235
rect 30934 56171 30986 56177
rect 29110 49717 29162 49723
rect 29110 49659 29162 49665
rect 29014 44759 29066 44765
rect 29014 44701 29066 44707
rect 28822 12125 28874 12131
rect 28822 12067 28874 12073
rect 29026 7913 29054 44701
rect 29014 7907 29066 7913
rect 29014 7849 29066 7855
rect 29122 7747 29150 49659
rect 29206 20931 29258 20937
rect 29206 20873 29258 20879
rect 29026 7719 29150 7747
rect 29026 7173 29054 7719
rect 29218 7636 29246 20873
rect 29602 17294 29630 56171
rect 29782 55415 29834 55421
rect 29782 55357 29834 55363
rect 29122 7608 29246 7636
rect 29506 17266 29630 17294
rect 28342 7167 28394 7173
rect 28342 7109 28394 7115
rect 29014 7167 29066 7173
rect 29014 7109 29066 7115
rect 28534 7019 28586 7025
rect 28534 6961 28586 6967
rect 28342 4355 28394 4361
rect 28342 4297 28394 4303
rect 28246 3245 28298 3251
rect 28246 3187 28298 3193
rect 28258 800 28286 3187
rect 28354 800 28382 4297
rect 28546 800 28574 6961
rect 29122 6433 29150 7608
rect 29206 7463 29258 7469
rect 29206 7405 29258 7411
rect 29110 6427 29162 6433
rect 29110 6369 29162 6375
rect 28822 5687 28874 5693
rect 28822 5629 28874 5635
rect 28834 4232 28862 5629
rect 28918 5021 28970 5027
rect 28918 4963 28970 4969
rect 28642 4204 28862 4232
rect 28642 800 28670 4204
rect 28930 3917 28958 4963
rect 29110 4355 29162 4361
rect 29110 4297 29162 4303
rect 28918 3911 28970 3917
rect 28918 3853 28970 3859
rect 29014 3911 29066 3917
rect 29014 3853 29066 3859
rect 28726 3763 28778 3769
rect 28726 3705 28778 3711
rect 28738 800 28766 3705
rect 28918 3541 28970 3547
rect 28918 3483 28970 3489
rect 28930 800 28958 3483
rect 29026 800 29054 3853
rect 29122 800 29150 4297
rect 29218 800 29246 7405
rect 29506 5471 29534 17266
rect 29794 10207 29822 55357
rect 30166 55119 30218 55125
rect 30166 55061 30218 55067
rect 29782 10201 29834 10207
rect 29782 10143 29834 10149
rect 30178 7765 30206 55061
rect 30946 21011 30974 56171
rect 31234 56161 31262 59200
rect 31714 56975 31742 59200
rect 31702 56969 31754 56975
rect 31702 56911 31754 56917
rect 32290 56531 32318 59200
rect 32566 56895 32618 56901
rect 32566 56837 32618 56843
rect 32278 56525 32330 56531
rect 32278 56467 32330 56473
rect 31318 56229 31370 56235
rect 31318 56171 31370 56177
rect 32470 56229 32522 56235
rect 32470 56171 32522 56177
rect 31222 56155 31274 56161
rect 31222 56097 31274 56103
rect 31030 36249 31082 36255
rect 31030 36191 31082 36197
rect 30934 21005 30986 21011
rect 30934 20947 30986 20953
rect 30646 19821 30698 19827
rect 30646 19763 30698 19769
rect 30166 7759 30218 7765
rect 30166 7701 30218 7707
rect 29590 7463 29642 7469
rect 29590 7405 29642 7411
rect 29494 5465 29546 5471
rect 29494 5407 29546 5413
rect 29302 5021 29354 5027
rect 29302 4963 29354 4969
rect 29314 3251 29342 4963
rect 29398 3837 29450 3843
rect 29398 3779 29450 3785
rect 29302 3245 29354 3251
rect 29302 3187 29354 3193
rect 29410 800 29438 3779
rect 29494 3615 29546 3621
rect 29494 3557 29546 3563
rect 29506 800 29534 3557
rect 29602 800 29630 7405
rect 29974 6945 30026 6951
rect 29974 6887 30026 6893
rect 29686 6353 29738 6359
rect 29686 6295 29738 6301
rect 29698 800 29726 6295
rect 29782 6131 29834 6137
rect 29782 6073 29834 6079
rect 29794 3547 29822 6073
rect 29782 3541 29834 3547
rect 29782 3483 29834 3489
rect 29878 3023 29930 3029
rect 29878 2965 29930 2971
rect 29890 800 29918 2965
rect 29986 800 30014 6887
rect 30658 6433 30686 19763
rect 31042 7099 31070 36191
rect 31330 11761 31358 56171
rect 32374 55489 32426 55495
rect 32374 55431 32426 55437
rect 32386 55051 32414 55431
rect 32374 55045 32426 55051
rect 32374 54987 32426 54993
rect 31798 45203 31850 45209
rect 31798 45145 31850 45151
rect 31702 33659 31754 33665
rect 31702 33601 31754 33607
rect 31318 11755 31370 11761
rect 31318 11697 31370 11703
rect 31126 7463 31178 7469
rect 31126 7405 31178 7411
rect 31030 7093 31082 7099
rect 31030 7035 31082 7041
rect 30742 7019 30794 7025
rect 30742 6961 30794 6967
rect 30646 6427 30698 6433
rect 30646 6369 30698 6375
rect 30262 5687 30314 5693
rect 30262 5629 30314 5635
rect 30274 2894 30302 5629
rect 30358 5021 30410 5027
rect 30358 4963 30410 4969
rect 30454 5021 30506 5027
rect 30454 4963 30506 4969
rect 30370 3917 30398 4963
rect 30358 3911 30410 3917
rect 30358 3853 30410 3859
rect 30466 3843 30494 4963
rect 30454 3837 30506 3843
rect 30454 3779 30506 3785
rect 30454 3689 30506 3695
rect 30082 2866 30302 2894
rect 30370 3649 30454 3677
rect 30082 800 30110 2866
rect 30370 1864 30398 3649
rect 30454 3631 30506 3637
rect 30454 3541 30506 3547
rect 30454 3483 30506 3489
rect 30274 1836 30398 1864
rect 30274 800 30302 1836
rect 30358 1765 30410 1771
rect 30358 1707 30410 1713
rect 30370 800 30398 1707
rect 30466 800 30494 3483
rect 30550 3097 30602 3103
rect 30550 3039 30602 3045
rect 30562 800 30590 3039
rect 30754 800 30782 6961
rect 30838 5687 30890 5693
rect 30838 5629 30890 5635
rect 30850 800 30878 5629
rect 30934 4355 30986 4361
rect 30934 4297 30986 4303
rect 30946 800 30974 4297
rect 31138 2894 31166 7405
rect 31714 7099 31742 33601
rect 31702 7093 31754 7099
rect 31702 7035 31754 7041
rect 31702 6945 31754 6951
rect 31426 6905 31702 6933
rect 31222 6353 31274 6359
rect 31222 6295 31274 6301
rect 31042 2866 31166 2894
rect 31042 800 31070 2866
rect 31234 800 31262 6295
rect 31318 3689 31370 3695
rect 31318 3631 31370 3637
rect 31330 800 31358 3631
rect 31426 800 31454 6905
rect 31702 6887 31754 6893
rect 31810 6581 31838 45145
rect 32182 30329 32234 30335
rect 32182 30271 32234 30277
rect 32194 7173 32222 30271
rect 32278 21449 32330 21455
rect 32278 21391 32330 21397
rect 32290 21233 32318 21391
rect 32278 21227 32330 21233
rect 32278 21169 32330 21175
rect 32482 17607 32510 56171
rect 32578 21899 32606 56837
rect 32770 56161 32798 59200
rect 33346 56975 33374 59200
rect 33334 56969 33386 56975
rect 33334 56911 33386 56917
rect 33826 56531 33854 59200
rect 34102 56895 34154 56901
rect 34102 56837 34154 56843
rect 33814 56525 33866 56531
rect 33814 56467 33866 56473
rect 32854 56229 32906 56235
rect 32854 56171 32906 56177
rect 34006 56229 34058 56235
rect 34006 56171 34058 56177
rect 32758 56155 32810 56161
rect 32758 56097 32810 56103
rect 32662 28849 32714 28855
rect 32662 28791 32714 28797
rect 32566 21893 32618 21899
rect 32566 21835 32618 21841
rect 32470 17601 32522 17607
rect 32470 17543 32522 17549
rect 32182 7167 32234 7173
rect 32182 7109 32234 7115
rect 32674 7099 32702 28791
rect 32866 11835 32894 56171
rect 33622 54231 33674 54237
rect 33622 54173 33674 54179
rect 33238 49421 33290 49427
rect 33238 49363 33290 49369
rect 33250 49131 33278 49363
rect 33238 49125 33290 49131
rect 33238 49067 33290 49073
rect 33334 40911 33386 40917
rect 33334 40853 33386 40859
rect 33346 40769 33374 40853
rect 33334 40763 33386 40769
rect 33334 40705 33386 40711
rect 33238 13457 33290 13463
rect 33238 13399 33290 13405
rect 32854 11829 32906 11835
rect 32854 11771 32906 11777
rect 33250 7099 33278 13399
rect 33346 7765 33374 40705
rect 33526 26259 33578 26265
rect 33526 26201 33578 26207
rect 33538 8135 33566 26201
rect 33634 12224 33662 54173
rect 34018 54089 34046 56171
rect 34006 54083 34058 54089
rect 34006 54025 34058 54031
rect 33718 34843 33770 34849
rect 33718 34785 33770 34791
rect 33730 17294 33758 34785
rect 33730 17266 33854 17294
rect 33634 12196 33758 12224
rect 33526 8129 33578 8135
rect 33526 8071 33578 8077
rect 33334 7759 33386 7765
rect 33334 7701 33386 7707
rect 33622 7463 33674 7469
rect 33622 7405 33674 7411
rect 32662 7093 32714 7099
rect 32662 7035 32714 7041
rect 33238 7093 33290 7099
rect 33238 7035 33290 7041
rect 32182 7019 32234 7025
rect 32182 6961 32234 6967
rect 31798 6575 31850 6581
rect 31798 6517 31850 6523
rect 31810 6433 31838 6517
rect 31798 6427 31850 6433
rect 31798 6369 31850 6375
rect 31798 6205 31850 6211
rect 31798 6147 31850 6153
rect 31510 6131 31562 6137
rect 31510 6073 31562 6079
rect 31522 1771 31550 6073
rect 31702 5687 31754 5693
rect 31702 5629 31754 5635
rect 31714 4528 31742 5629
rect 31618 4500 31742 4528
rect 31510 1765 31562 1771
rect 31510 1707 31562 1713
rect 31618 800 31646 4500
rect 31702 4355 31754 4361
rect 31702 4297 31754 4303
rect 31714 800 31742 4297
rect 31810 800 31838 6147
rect 31894 5021 31946 5027
rect 31894 4963 31946 4969
rect 31906 3547 31934 4963
rect 31894 3541 31946 3547
rect 31894 3483 31946 3489
rect 31894 3245 31946 3251
rect 31894 3187 31946 3193
rect 31906 800 31934 3187
rect 32086 3097 32138 3103
rect 32086 3039 32138 3045
rect 32098 800 32126 3039
rect 32194 800 32222 6961
rect 32566 6353 32618 6359
rect 32566 6295 32618 6301
rect 32470 3689 32522 3695
rect 32470 3631 32522 3637
rect 32278 3023 32330 3029
rect 32278 2965 32330 2971
rect 32290 800 32318 2965
rect 32482 800 32510 3631
rect 32578 800 32606 6295
rect 33526 6279 33578 6285
rect 33526 6221 33578 6227
rect 33142 5687 33194 5693
rect 33142 5629 33194 5635
rect 33238 5687 33290 5693
rect 33238 5629 33290 5635
rect 32758 4355 32810 4361
rect 32758 4297 32810 4303
rect 32662 3171 32714 3177
rect 32662 3113 32714 3119
rect 32674 800 32702 3113
rect 32770 800 32798 4297
rect 32854 3615 32906 3621
rect 32854 3557 32906 3563
rect 32866 2456 32894 3557
rect 33154 3029 33182 5629
rect 33142 3023 33194 3029
rect 33142 2965 33194 2971
rect 33250 2900 33278 5629
rect 33538 5471 33566 6221
rect 33526 5465 33578 5471
rect 33526 5407 33578 5413
rect 33334 5021 33386 5027
rect 33334 4963 33386 4969
rect 33346 3251 33374 4963
rect 33430 3837 33482 3843
rect 33430 3779 33482 3785
rect 33334 3245 33386 3251
rect 33334 3187 33386 3193
rect 33334 3097 33386 3103
rect 33334 3039 33386 3045
rect 33058 2872 33278 2900
rect 32950 2801 33002 2807
rect 32950 2743 33002 2749
rect 32962 2585 32990 2743
rect 32950 2579 33002 2585
rect 32950 2521 33002 2527
rect 32866 2428 32990 2456
rect 32962 800 32990 2428
rect 33058 800 33086 2872
rect 33346 1568 33374 3039
rect 33154 1540 33374 1568
rect 33154 800 33182 1540
rect 33238 1469 33290 1475
rect 33238 1411 33290 1417
rect 33250 800 33278 1411
rect 33442 800 33470 3779
rect 33526 3689 33578 3695
rect 33526 3631 33578 3637
rect 33538 800 33566 3631
rect 33634 800 33662 7405
rect 33730 7173 33758 12196
rect 33826 7765 33854 17266
rect 34114 12871 34142 56837
rect 34402 56531 34430 59200
rect 34882 56975 34910 59200
rect 34988 57304 35284 57324
rect 35044 57302 35068 57304
rect 35124 57302 35148 57304
rect 35204 57302 35228 57304
rect 35066 57250 35068 57302
rect 35130 57250 35142 57302
rect 35204 57250 35206 57302
rect 35044 57248 35068 57250
rect 35124 57248 35148 57250
rect 35204 57248 35228 57250
rect 34988 57228 35284 57248
rect 34870 56969 34922 56975
rect 34870 56911 34922 56917
rect 34390 56525 34442 56531
rect 34390 56467 34442 56473
rect 34774 56229 34826 56235
rect 34774 56171 34826 56177
rect 34582 43723 34634 43729
rect 34582 43665 34634 43671
rect 34294 18193 34346 18199
rect 34294 18135 34346 18141
rect 34102 12865 34154 12871
rect 34102 12807 34154 12813
rect 33814 7759 33866 7765
rect 33814 7701 33866 7707
rect 33718 7167 33770 7173
rect 33718 7109 33770 7115
rect 33718 6945 33770 6951
rect 34102 6945 34154 6951
rect 33718 6887 33770 6893
rect 34018 6905 34102 6933
rect 33730 3621 33758 6887
rect 33814 6131 33866 6137
rect 33814 6073 33866 6079
rect 33718 3615 33770 3621
rect 33718 3557 33770 3563
rect 33826 3492 33854 6073
rect 33910 4355 33962 4361
rect 33910 4297 33962 4303
rect 33730 3464 33854 3492
rect 33730 1475 33758 3464
rect 33814 3245 33866 3251
rect 33814 3187 33866 3193
rect 33718 1469 33770 1475
rect 33718 1411 33770 1417
rect 33826 800 33854 3187
rect 33922 800 33950 4297
rect 34018 800 34046 6905
rect 34102 6887 34154 6893
rect 34306 6433 34334 18135
rect 34594 7765 34622 43665
rect 34786 33591 34814 56171
rect 35458 56161 35486 59200
rect 35938 56513 35966 59200
rect 36514 56901 36542 59200
rect 36994 57614 37022 59200
rect 36994 57586 37118 57614
rect 36502 56895 36554 56901
rect 36502 56837 36554 56843
rect 36694 56747 36746 56753
rect 36694 56689 36746 56695
rect 36022 56525 36074 56531
rect 35938 56485 36022 56513
rect 36022 56467 36074 56473
rect 36022 56303 36074 56309
rect 36022 56245 36074 56251
rect 35830 56229 35882 56235
rect 35830 56171 35882 56177
rect 35446 56155 35498 56161
rect 35446 56097 35498 56103
rect 34988 55972 35284 55992
rect 35044 55970 35068 55972
rect 35124 55970 35148 55972
rect 35204 55970 35228 55972
rect 35066 55918 35068 55970
rect 35130 55918 35142 55970
rect 35204 55918 35206 55970
rect 35044 55916 35068 55918
rect 35124 55916 35148 55918
rect 35204 55916 35228 55918
rect 34988 55896 35284 55916
rect 34988 54640 35284 54660
rect 35044 54638 35068 54640
rect 35124 54638 35148 54640
rect 35204 54638 35228 54640
rect 35066 54586 35068 54638
rect 35130 54586 35142 54638
rect 35204 54586 35206 54638
rect 35044 54584 35068 54586
rect 35124 54584 35148 54586
rect 35204 54584 35228 54586
rect 34988 54564 35284 54584
rect 34988 53308 35284 53328
rect 35044 53306 35068 53308
rect 35124 53306 35148 53308
rect 35204 53306 35228 53308
rect 35066 53254 35068 53306
rect 35130 53254 35142 53306
rect 35204 53254 35206 53306
rect 35044 53252 35068 53254
rect 35124 53252 35148 53254
rect 35204 53252 35228 53254
rect 34988 53232 35284 53252
rect 34988 51976 35284 51996
rect 35044 51974 35068 51976
rect 35124 51974 35148 51976
rect 35204 51974 35228 51976
rect 35066 51922 35068 51974
rect 35130 51922 35142 51974
rect 35204 51922 35206 51974
rect 35044 51920 35068 51922
rect 35124 51920 35148 51922
rect 35204 51920 35228 51922
rect 34988 51900 35284 51920
rect 34988 50644 35284 50664
rect 35044 50642 35068 50644
rect 35124 50642 35148 50644
rect 35204 50642 35228 50644
rect 35066 50590 35068 50642
rect 35130 50590 35142 50642
rect 35204 50590 35206 50642
rect 35044 50588 35068 50590
rect 35124 50588 35148 50590
rect 35204 50588 35228 50590
rect 34988 50568 35284 50588
rect 34988 49312 35284 49332
rect 35044 49310 35068 49312
rect 35124 49310 35148 49312
rect 35204 49310 35228 49312
rect 35066 49258 35068 49310
rect 35130 49258 35142 49310
rect 35204 49258 35206 49310
rect 35044 49256 35068 49258
rect 35124 49256 35148 49258
rect 35204 49256 35228 49258
rect 34988 49236 35284 49256
rect 34988 47980 35284 48000
rect 35044 47978 35068 47980
rect 35124 47978 35148 47980
rect 35204 47978 35228 47980
rect 35066 47926 35068 47978
rect 35130 47926 35142 47978
rect 35204 47926 35206 47978
rect 35044 47924 35068 47926
rect 35124 47924 35148 47926
rect 35204 47924 35228 47926
rect 34988 47904 35284 47924
rect 34988 46648 35284 46668
rect 35044 46646 35068 46648
rect 35124 46646 35148 46648
rect 35204 46646 35228 46648
rect 35066 46594 35068 46646
rect 35130 46594 35142 46646
rect 35204 46594 35206 46646
rect 35044 46592 35068 46594
rect 35124 46592 35148 46594
rect 35204 46592 35228 46594
rect 34988 46572 35284 46592
rect 34988 45316 35284 45336
rect 35044 45314 35068 45316
rect 35124 45314 35148 45316
rect 35204 45314 35228 45316
rect 35066 45262 35068 45314
rect 35130 45262 35142 45314
rect 35204 45262 35206 45314
rect 35044 45260 35068 45262
rect 35124 45260 35148 45262
rect 35204 45260 35228 45262
rect 34988 45240 35284 45260
rect 34988 43984 35284 44004
rect 35044 43982 35068 43984
rect 35124 43982 35148 43984
rect 35204 43982 35228 43984
rect 35066 43930 35068 43982
rect 35130 43930 35142 43982
rect 35204 43930 35206 43982
rect 35044 43928 35068 43930
rect 35124 43928 35148 43930
rect 35204 43928 35228 43930
rect 34988 43908 35284 43928
rect 34988 42652 35284 42672
rect 35044 42650 35068 42652
rect 35124 42650 35148 42652
rect 35204 42650 35228 42652
rect 35066 42598 35068 42650
rect 35130 42598 35142 42650
rect 35204 42598 35206 42650
rect 35044 42596 35068 42598
rect 35124 42596 35148 42598
rect 35204 42596 35228 42598
rect 34988 42576 35284 42596
rect 34988 41320 35284 41340
rect 35044 41318 35068 41320
rect 35124 41318 35148 41320
rect 35204 41318 35228 41320
rect 35066 41266 35068 41318
rect 35130 41266 35142 41318
rect 35204 41266 35206 41318
rect 35044 41264 35068 41266
rect 35124 41264 35148 41266
rect 35204 41264 35228 41266
rect 34988 41244 35284 41264
rect 34988 39988 35284 40008
rect 35044 39986 35068 39988
rect 35124 39986 35148 39988
rect 35204 39986 35228 39988
rect 35066 39934 35068 39986
rect 35130 39934 35142 39986
rect 35204 39934 35206 39986
rect 35044 39932 35068 39934
rect 35124 39932 35148 39934
rect 35204 39932 35228 39934
rect 34988 39912 35284 39932
rect 34988 38656 35284 38676
rect 35044 38654 35068 38656
rect 35124 38654 35148 38656
rect 35204 38654 35228 38656
rect 35066 38602 35068 38654
rect 35130 38602 35142 38654
rect 35204 38602 35206 38654
rect 35044 38600 35068 38602
rect 35124 38600 35148 38602
rect 35204 38600 35228 38602
rect 34988 38580 35284 38600
rect 34988 37324 35284 37344
rect 35044 37322 35068 37324
rect 35124 37322 35148 37324
rect 35204 37322 35228 37324
rect 35066 37270 35068 37322
rect 35130 37270 35142 37322
rect 35204 37270 35206 37322
rect 35044 37268 35068 37270
rect 35124 37268 35148 37270
rect 35204 37268 35228 37270
rect 34988 37248 35284 37268
rect 34988 35992 35284 36012
rect 35044 35990 35068 35992
rect 35124 35990 35148 35992
rect 35204 35990 35228 35992
rect 35066 35938 35068 35990
rect 35130 35938 35142 35990
rect 35204 35938 35206 35990
rect 35044 35936 35068 35938
rect 35124 35936 35148 35938
rect 35204 35936 35228 35938
rect 34988 35916 35284 35936
rect 34988 34660 35284 34680
rect 35044 34658 35068 34660
rect 35124 34658 35148 34660
rect 35204 34658 35228 34660
rect 35066 34606 35068 34658
rect 35130 34606 35142 34658
rect 35204 34606 35206 34658
rect 35044 34604 35068 34606
rect 35124 34604 35148 34606
rect 35204 34604 35228 34606
rect 34988 34584 35284 34604
rect 34774 33585 34826 33591
rect 34774 33527 34826 33533
rect 35350 33511 35402 33517
rect 35350 33453 35402 33459
rect 34678 33437 34730 33443
rect 34678 33379 34730 33385
rect 34690 8579 34718 33379
rect 34988 33328 35284 33348
rect 35044 33326 35068 33328
rect 35124 33326 35148 33328
rect 35204 33326 35228 33328
rect 35066 33274 35068 33326
rect 35130 33274 35142 33326
rect 35204 33274 35206 33326
rect 35044 33272 35068 33274
rect 35124 33272 35148 33274
rect 35204 33272 35228 33274
rect 34988 33252 35284 33272
rect 34988 31996 35284 32016
rect 35044 31994 35068 31996
rect 35124 31994 35148 31996
rect 35204 31994 35228 31996
rect 35066 31942 35068 31994
rect 35130 31942 35142 31994
rect 35204 31942 35206 31994
rect 35044 31940 35068 31942
rect 35124 31940 35148 31942
rect 35204 31940 35228 31942
rect 34988 31920 35284 31940
rect 34774 30773 34826 30779
rect 34774 30715 34826 30721
rect 34678 8573 34730 8579
rect 34678 8515 34730 8521
rect 34582 7759 34634 7765
rect 34582 7701 34634 7707
rect 34486 7611 34538 7617
rect 34486 7553 34538 7559
rect 34390 7463 34442 7469
rect 34390 7405 34442 7411
rect 34294 6427 34346 6433
rect 34294 6369 34346 6375
rect 34102 5021 34154 5027
rect 34102 4963 34154 4969
rect 34114 3177 34142 4963
rect 34198 4281 34250 4287
rect 34198 4223 34250 4229
rect 34102 3171 34154 3177
rect 34102 3113 34154 3119
rect 34210 2160 34238 4223
rect 34294 3689 34346 3695
rect 34294 3631 34346 3637
rect 34114 2132 34238 2160
rect 34114 800 34142 2132
rect 34306 800 34334 3631
rect 34402 800 34430 7405
rect 34498 7025 34526 7553
rect 34678 7463 34730 7469
rect 34678 7405 34730 7411
rect 34486 7019 34538 7025
rect 34486 6961 34538 6967
rect 34582 4947 34634 4953
rect 34582 4889 34634 4895
rect 34594 4528 34622 4889
rect 34498 4500 34622 4528
rect 34498 800 34526 4500
rect 34582 4355 34634 4361
rect 34582 4297 34634 4303
rect 34594 800 34622 4297
rect 34690 3640 34718 7405
rect 34786 7099 34814 30715
rect 34988 30664 35284 30684
rect 35044 30662 35068 30664
rect 35124 30662 35148 30664
rect 35204 30662 35228 30664
rect 35066 30610 35068 30662
rect 35130 30610 35142 30662
rect 35204 30610 35206 30662
rect 35044 30608 35068 30610
rect 35124 30608 35148 30610
rect 35204 30608 35228 30610
rect 34988 30588 35284 30608
rect 34988 29332 35284 29352
rect 35044 29330 35068 29332
rect 35124 29330 35148 29332
rect 35204 29330 35228 29332
rect 35066 29278 35068 29330
rect 35130 29278 35142 29330
rect 35204 29278 35206 29330
rect 35044 29276 35068 29278
rect 35124 29276 35148 29278
rect 35204 29276 35228 29278
rect 34988 29256 35284 29276
rect 34988 28000 35284 28020
rect 35044 27998 35068 28000
rect 35124 27998 35148 28000
rect 35204 27998 35228 28000
rect 35066 27946 35068 27998
rect 35130 27946 35142 27998
rect 35204 27946 35206 27998
rect 35044 27944 35068 27946
rect 35124 27944 35148 27946
rect 35204 27944 35228 27946
rect 34988 27924 35284 27944
rect 34988 26668 35284 26688
rect 35044 26666 35068 26668
rect 35124 26666 35148 26668
rect 35204 26666 35228 26668
rect 35066 26614 35068 26666
rect 35130 26614 35142 26666
rect 35204 26614 35206 26666
rect 35044 26612 35068 26614
rect 35124 26612 35148 26614
rect 35204 26612 35228 26614
rect 34988 26592 35284 26612
rect 34988 25336 35284 25356
rect 35044 25334 35068 25336
rect 35124 25334 35148 25336
rect 35204 25334 35228 25336
rect 35066 25282 35068 25334
rect 35130 25282 35142 25334
rect 35204 25282 35206 25334
rect 35044 25280 35068 25282
rect 35124 25280 35148 25282
rect 35204 25280 35228 25282
rect 34988 25260 35284 25280
rect 34988 24004 35284 24024
rect 35044 24002 35068 24004
rect 35124 24002 35148 24004
rect 35204 24002 35228 24004
rect 35066 23950 35068 24002
rect 35130 23950 35142 24002
rect 35204 23950 35206 24002
rect 35044 23948 35068 23950
rect 35124 23948 35148 23950
rect 35204 23948 35228 23950
rect 34988 23928 35284 23948
rect 34988 22672 35284 22692
rect 35044 22670 35068 22672
rect 35124 22670 35148 22672
rect 35204 22670 35228 22672
rect 35066 22618 35068 22670
rect 35130 22618 35142 22670
rect 35204 22618 35206 22670
rect 35044 22616 35068 22618
rect 35124 22616 35148 22618
rect 35204 22616 35228 22618
rect 34988 22596 35284 22616
rect 34988 21340 35284 21360
rect 35044 21338 35068 21340
rect 35124 21338 35148 21340
rect 35204 21338 35228 21340
rect 35066 21286 35068 21338
rect 35130 21286 35142 21338
rect 35204 21286 35206 21338
rect 35044 21284 35068 21286
rect 35124 21284 35148 21286
rect 35204 21284 35228 21286
rect 34988 21264 35284 21284
rect 34988 20008 35284 20028
rect 35044 20006 35068 20008
rect 35124 20006 35148 20008
rect 35204 20006 35228 20008
rect 35066 19954 35068 20006
rect 35130 19954 35142 20006
rect 35204 19954 35206 20006
rect 35044 19952 35068 19954
rect 35124 19952 35148 19954
rect 35204 19952 35228 19954
rect 34988 19932 35284 19952
rect 34988 18676 35284 18696
rect 35044 18674 35068 18676
rect 35124 18674 35148 18676
rect 35204 18674 35228 18676
rect 35066 18622 35068 18674
rect 35130 18622 35142 18674
rect 35204 18622 35206 18674
rect 35044 18620 35068 18622
rect 35124 18620 35148 18622
rect 35204 18620 35228 18622
rect 34988 18600 35284 18620
rect 34988 17344 35284 17364
rect 35044 17342 35068 17344
rect 35124 17342 35148 17344
rect 35204 17342 35228 17344
rect 35066 17290 35068 17342
rect 35130 17290 35142 17342
rect 35204 17290 35206 17342
rect 35044 17288 35068 17290
rect 35124 17288 35148 17290
rect 35204 17288 35228 17290
rect 34988 17268 35284 17288
rect 34988 16012 35284 16032
rect 35044 16010 35068 16012
rect 35124 16010 35148 16012
rect 35204 16010 35228 16012
rect 35066 15958 35068 16010
rect 35130 15958 35142 16010
rect 35204 15958 35206 16010
rect 35044 15956 35068 15958
rect 35124 15956 35148 15958
rect 35204 15956 35228 15958
rect 34988 15936 35284 15956
rect 34870 14937 34922 14943
rect 34870 14879 34922 14885
rect 34774 7093 34826 7099
rect 34774 7035 34826 7041
rect 34882 6433 34910 14879
rect 34988 14680 35284 14700
rect 35044 14678 35068 14680
rect 35124 14678 35148 14680
rect 35204 14678 35228 14680
rect 35066 14626 35068 14678
rect 35130 14626 35142 14678
rect 35204 14626 35206 14678
rect 35044 14624 35068 14626
rect 35124 14624 35148 14626
rect 35204 14624 35228 14626
rect 34988 14604 35284 14624
rect 34988 13348 35284 13368
rect 35044 13346 35068 13348
rect 35124 13346 35148 13348
rect 35204 13346 35228 13348
rect 35066 13294 35068 13346
rect 35130 13294 35142 13346
rect 35204 13294 35206 13346
rect 35044 13292 35068 13294
rect 35124 13292 35148 13294
rect 35204 13292 35228 13294
rect 34988 13272 35284 13292
rect 34988 12016 35284 12036
rect 35044 12014 35068 12016
rect 35124 12014 35148 12016
rect 35204 12014 35228 12016
rect 35066 11962 35068 12014
rect 35130 11962 35142 12014
rect 35204 11962 35206 12014
rect 35044 11960 35068 11962
rect 35124 11960 35148 11962
rect 35204 11960 35228 11962
rect 34988 11940 35284 11960
rect 34988 10684 35284 10704
rect 35044 10682 35068 10684
rect 35124 10682 35148 10684
rect 35204 10682 35228 10684
rect 35066 10630 35068 10682
rect 35130 10630 35142 10682
rect 35204 10630 35206 10682
rect 35044 10628 35068 10630
rect 35124 10628 35148 10630
rect 35204 10628 35228 10630
rect 34988 10608 35284 10628
rect 34988 9352 35284 9372
rect 35044 9350 35068 9352
rect 35124 9350 35148 9352
rect 35204 9350 35228 9352
rect 35066 9298 35068 9350
rect 35130 9298 35142 9350
rect 35204 9298 35206 9350
rect 35044 9296 35068 9298
rect 35124 9296 35148 9298
rect 35204 9296 35228 9298
rect 34988 9276 35284 9296
rect 34988 8020 35284 8040
rect 35044 8018 35068 8020
rect 35124 8018 35148 8020
rect 35204 8018 35228 8020
rect 35066 7966 35068 8018
rect 35130 7966 35142 8018
rect 35204 7966 35206 8018
rect 35044 7964 35068 7966
rect 35124 7964 35148 7966
rect 35204 7964 35228 7966
rect 34988 7944 35284 7964
rect 35362 7765 35390 33453
rect 35842 11835 35870 56171
rect 36034 55643 36062 56245
rect 36598 56229 36650 56235
rect 36598 56171 36650 56177
rect 36022 55637 36074 55643
rect 36022 55579 36074 55585
rect 36406 46757 36458 46763
rect 36406 46699 36458 46705
rect 36214 19155 36266 19161
rect 36214 19097 36266 19103
rect 36118 18785 36170 18791
rect 36118 18727 36170 18733
rect 35830 11829 35882 11835
rect 35830 11771 35882 11777
rect 36130 7765 36158 18727
rect 35350 7759 35402 7765
rect 35350 7701 35402 7707
rect 36118 7759 36170 7765
rect 36118 7701 36170 7707
rect 36022 7463 36074 7469
rect 36022 7405 36074 7411
rect 35542 6945 35594 6951
rect 35542 6887 35594 6893
rect 34988 6688 35284 6708
rect 35044 6686 35068 6688
rect 35124 6686 35148 6688
rect 35204 6686 35228 6688
rect 35066 6634 35068 6686
rect 35130 6634 35142 6686
rect 35204 6634 35206 6686
rect 35044 6632 35068 6634
rect 35124 6632 35148 6634
rect 35204 6632 35228 6634
rect 34988 6612 35284 6632
rect 34870 6427 34922 6433
rect 34870 6369 34922 6375
rect 35350 6131 35402 6137
rect 35350 6073 35402 6079
rect 34774 5687 34826 5693
rect 34774 5629 34826 5635
rect 34786 3751 34814 5629
rect 34988 5356 35284 5376
rect 35044 5354 35068 5356
rect 35124 5354 35148 5356
rect 35204 5354 35228 5356
rect 35066 5302 35068 5354
rect 35130 5302 35142 5354
rect 35204 5302 35206 5354
rect 35044 5300 35068 5302
rect 35124 5300 35148 5302
rect 35204 5300 35228 5302
rect 34988 5280 35284 5300
rect 34870 5021 34922 5027
rect 34870 4963 34922 4969
rect 34882 3843 34910 4963
rect 34988 4024 35284 4044
rect 35044 4022 35068 4024
rect 35124 4022 35148 4024
rect 35204 4022 35228 4024
rect 35066 3970 35068 4022
rect 35130 3970 35142 4022
rect 35204 3970 35206 4022
rect 35044 3968 35068 3970
rect 35124 3968 35148 3970
rect 35204 3968 35228 3970
rect 34988 3948 35284 3968
rect 34870 3837 34922 3843
rect 34870 3779 34922 3785
rect 34786 3723 35102 3751
rect 34966 3689 35018 3695
rect 34882 3649 34966 3677
rect 34690 3612 34814 3640
rect 34678 3171 34730 3177
rect 34678 3113 34730 3119
rect 34690 1475 34718 3113
rect 34678 1469 34730 1475
rect 34678 1411 34730 1417
rect 34786 800 34814 3612
rect 34882 1864 34910 3649
rect 34966 3631 35018 3637
rect 35074 3251 35102 3723
rect 35062 3245 35114 3251
rect 35062 3187 35114 3193
rect 35362 3177 35390 6073
rect 35350 3171 35402 3177
rect 35350 3113 35402 3119
rect 35446 3097 35498 3103
rect 35446 3039 35498 3045
rect 35350 3023 35402 3029
rect 35350 2965 35402 2971
rect 34988 2692 35284 2712
rect 35044 2690 35068 2692
rect 35124 2690 35148 2692
rect 35204 2690 35228 2692
rect 35066 2638 35068 2690
rect 35130 2638 35142 2690
rect 35204 2638 35206 2690
rect 35044 2636 35068 2638
rect 35124 2636 35148 2638
rect 35204 2636 35228 2638
rect 34988 2616 35284 2636
rect 35158 2579 35210 2585
rect 35158 2521 35210 2527
rect 34882 1836 35006 1864
rect 34870 1765 34922 1771
rect 34870 1707 34922 1713
rect 34882 800 34910 1707
rect 34978 800 35006 1836
rect 35170 800 35198 2521
rect 35362 2456 35390 2965
rect 35266 2428 35390 2456
rect 35266 800 35294 2428
rect 35458 1568 35486 3039
rect 35554 2585 35582 6887
rect 35638 3837 35690 3843
rect 35638 3779 35690 3785
rect 35542 2579 35594 2585
rect 35542 2521 35594 2527
rect 35650 1771 35678 3779
rect 35734 3689 35786 3695
rect 36034 3640 36062 7405
rect 36226 7099 36254 19097
rect 36214 7093 36266 7099
rect 36214 7035 36266 7041
rect 36418 6803 36446 46699
rect 36502 21745 36554 21751
rect 36502 21687 36554 21693
rect 36514 7913 36542 21687
rect 36610 13167 36638 56171
rect 36706 14351 36734 56689
rect 37090 56161 37118 57586
rect 37570 56531 37598 59200
rect 38050 56975 38078 59200
rect 38038 56969 38090 56975
rect 38038 56911 38090 56917
rect 38626 56531 38654 59200
rect 37558 56525 37610 56531
rect 37558 56467 37610 56473
rect 38614 56525 38666 56531
rect 38614 56467 38666 56473
rect 37078 56155 37130 56161
rect 37078 56097 37130 56103
rect 39106 55717 39134 59200
rect 39682 56901 39710 59200
rect 39670 56895 39722 56901
rect 39670 56837 39722 56843
rect 39766 56747 39818 56753
rect 39766 56689 39818 56695
rect 39094 55711 39146 55717
rect 39094 55653 39146 55659
rect 38902 55563 38954 55569
rect 38902 55505 38954 55511
rect 38914 55421 38942 55505
rect 38902 55415 38954 55421
rect 38902 55357 38954 55363
rect 36790 54971 36842 54977
rect 36790 54913 36842 54919
rect 36694 14345 36746 14351
rect 36694 14287 36746 14293
rect 36598 13161 36650 13167
rect 36598 13103 36650 13109
rect 36802 9615 36830 54913
rect 37750 48089 37802 48095
rect 37750 48031 37802 48037
rect 37174 36323 37226 36329
rect 37174 36265 37226 36271
rect 37186 36107 37214 36265
rect 37174 36101 37226 36107
rect 37174 36043 37226 36049
rect 36790 9609 36842 9615
rect 36790 9551 36842 9557
rect 37270 9461 37322 9467
rect 37270 9403 37322 9409
rect 36502 7907 36554 7913
rect 36502 7849 36554 7855
rect 36598 7463 36650 7469
rect 36598 7405 36650 7411
rect 36502 6945 36554 6951
rect 36502 6887 36554 6893
rect 36406 6797 36458 6803
rect 36406 6739 36458 6745
rect 36310 6353 36362 6359
rect 36310 6295 36362 6301
rect 36118 5687 36170 5693
rect 36118 5629 36170 5635
rect 36214 5687 36266 5693
rect 36214 5629 36266 5635
rect 35734 3631 35786 3637
rect 35638 1765 35690 1771
rect 35638 1707 35690 1713
rect 35362 1540 35486 1568
rect 35638 1617 35690 1623
rect 35638 1559 35690 1565
rect 35362 800 35390 1540
rect 35446 1469 35498 1475
rect 35446 1411 35498 1417
rect 35458 800 35486 1411
rect 35650 800 35678 1559
rect 35746 800 35774 3631
rect 35842 3612 36062 3640
rect 35842 800 35870 3612
rect 35926 3541 35978 3547
rect 35926 3483 35978 3489
rect 35938 1623 35966 3483
rect 36022 3467 36074 3473
rect 36022 3409 36074 3415
rect 35926 1617 35978 1623
rect 35926 1559 35978 1565
rect 36034 800 36062 3409
rect 36130 3029 36158 5629
rect 36226 3473 36254 5629
rect 36214 3467 36266 3473
rect 36214 3409 36266 3415
rect 36214 3171 36266 3177
rect 36214 3113 36266 3119
rect 36118 3023 36170 3029
rect 36118 2965 36170 2971
rect 36226 1568 36254 3113
rect 36130 1540 36254 1568
rect 36322 1549 36350 6295
rect 36406 5021 36458 5027
rect 36406 4963 36458 4969
rect 36418 3843 36446 4963
rect 36406 3837 36458 3843
rect 36406 3779 36458 3785
rect 36514 3751 36542 6887
rect 36418 3723 36542 3751
rect 36310 1543 36362 1549
rect 36130 800 36158 1540
rect 36310 1485 36362 1491
rect 36418 1420 36446 3723
rect 36502 3689 36554 3695
rect 36502 3631 36554 3637
rect 36226 1392 36446 1420
rect 36226 800 36254 1392
rect 36310 1173 36362 1179
rect 36310 1115 36362 1121
rect 36322 800 36350 1115
rect 36514 800 36542 3631
rect 36610 800 36638 7405
rect 37078 6945 37130 6951
rect 36994 6905 37078 6933
rect 36694 5021 36746 5027
rect 36694 4963 36746 4969
rect 36706 3547 36734 4963
rect 36790 4355 36842 4361
rect 36790 4297 36842 4303
rect 36694 3541 36746 3547
rect 36694 3483 36746 3489
rect 36694 3245 36746 3251
rect 36694 3187 36746 3193
rect 36706 800 36734 3187
rect 36802 800 36830 4297
rect 36994 800 37022 6905
rect 37078 6887 37130 6893
rect 37282 6433 37310 9403
rect 37654 7167 37706 7173
rect 37654 7109 37706 7115
rect 37366 7019 37418 7025
rect 37366 6961 37418 6967
rect 37270 6427 37322 6433
rect 37270 6369 37322 6375
rect 37174 4281 37226 4287
rect 37174 4223 37226 4229
rect 37078 3467 37130 3473
rect 37078 3409 37130 3415
rect 37090 800 37118 3409
rect 37186 800 37214 4223
rect 37378 800 37406 6961
rect 37462 5761 37514 5767
rect 37462 5703 37514 5709
rect 37474 800 37502 5703
rect 37558 5687 37610 5693
rect 37558 5629 37610 5635
rect 37570 3251 37598 5629
rect 37558 3245 37610 3251
rect 37558 3187 37610 3193
rect 37558 3023 37610 3029
rect 37558 2965 37610 2971
rect 37570 800 37598 2965
rect 37666 800 37694 7109
rect 37762 7099 37790 48031
rect 38710 38765 38762 38771
rect 38710 38707 38762 38713
rect 38230 33437 38282 33443
rect 38230 33379 38282 33385
rect 38038 7463 38090 7469
rect 38038 7405 38090 7411
rect 37750 7093 37802 7099
rect 37750 7035 37802 7041
rect 37846 3837 37898 3843
rect 37846 3779 37898 3785
rect 37750 3763 37802 3769
rect 37750 3705 37802 3711
rect 37762 2955 37790 3705
rect 37750 2949 37802 2955
rect 37750 2891 37802 2897
rect 37858 800 37886 3779
rect 37942 3689 37994 3695
rect 37942 3631 37994 3637
rect 37954 800 37982 3631
rect 38050 800 38078 7405
rect 38242 6877 38270 33379
rect 38518 12125 38570 12131
rect 38518 12067 38570 12073
rect 38530 7099 38558 12067
rect 38722 7765 38750 38707
rect 38914 14129 38942 55357
rect 39478 48903 39530 48909
rect 39478 48845 39530 48851
rect 38902 14123 38954 14129
rect 38902 14065 38954 14071
rect 38806 10275 38858 10281
rect 38806 10217 38858 10223
rect 38818 7839 38846 10217
rect 38806 7833 38858 7839
rect 38806 7775 38858 7781
rect 39490 7765 39518 48845
rect 39778 15535 39806 56689
rect 40162 56531 40190 59200
rect 40438 56747 40490 56753
rect 40438 56689 40490 56695
rect 40150 56525 40202 56531
rect 40150 56467 40202 56473
rect 40246 56229 40298 56235
rect 40246 56171 40298 56177
rect 40258 40769 40286 56171
rect 40246 40763 40298 40769
rect 40246 40705 40298 40711
rect 40450 26117 40478 56689
rect 40738 55717 40766 59200
rect 41218 56975 41246 59200
rect 41206 56969 41258 56975
rect 41206 56911 41258 56917
rect 40822 56747 40874 56753
rect 40822 56689 40874 56695
rect 40834 56161 40862 56689
rect 41794 56531 41822 59200
rect 42274 56531 42302 59200
rect 42850 56901 42878 59200
rect 42838 56895 42890 56901
rect 42838 56837 42890 56843
rect 42934 56747 42986 56753
rect 42934 56689 42986 56695
rect 41782 56525 41834 56531
rect 41782 56467 41834 56473
rect 42262 56525 42314 56531
rect 42262 56467 42314 56473
rect 42070 56229 42122 56235
rect 42070 56171 42122 56177
rect 42358 56229 42410 56235
rect 42358 56171 42410 56177
rect 40822 56155 40874 56161
rect 40822 56097 40874 56103
rect 40726 55711 40778 55717
rect 40726 55653 40778 55659
rect 40918 55563 40970 55569
rect 40918 55505 40970 55511
rect 40930 54755 40958 55505
rect 40918 54749 40970 54755
rect 40918 54691 40970 54697
rect 41110 44093 41162 44099
rect 41110 44035 41162 44041
rect 40438 26111 40490 26117
rect 40438 26053 40490 26059
rect 39958 18785 40010 18791
rect 39958 18727 40010 18733
rect 39766 15529 39818 15535
rect 39766 15471 39818 15477
rect 38710 7759 38762 7765
rect 38710 7701 38762 7707
rect 39478 7759 39530 7765
rect 39478 7701 39530 7707
rect 38806 7685 38858 7691
rect 38806 7627 38858 7633
rect 38518 7093 38570 7099
rect 38518 7035 38570 7041
rect 38518 6945 38570 6951
rect 38434 6905 38518 6933
rect 38134 6871 38186 6877
rect 38134 6813 38186 6819
rect 38230 6871 38282 6877
rect 38230 6813 38282 6819
rect 38146 6285 38174 6813
rect 38134 6279 38186 6285
rect 38134 6221 38186 6227
rect 38134 5243 38186 5249
rect 38134 5185 38186 5191
rect 38146 4583 38174 5185
rect 38134 4577 38186 4583
rect 38134 4519 38186 4525
rect 38326 3097 38378 3103
rect 38326 3039 38378 3045
rect 38134 2949 38186 2955
rect 38134 2891 38186 2897
rect 38146 800 38174 2891
rect 38338 800 38366 3039
rect 38434 800 38462 6905
rect 38518 6887 38570 6893
rect 38614 5021 38666 5027
rect 38614 4963 38666 4969
rect 38518 3911 38570 3917
rect 38518 3853 38570 3859
rect 38530 800 38558 3853
rect 38626 3473 38654 4963
rect 38710 3689 38762 3695
rect 38710 3631 38762 3637
rect 38614 3467 38666 3473
rect 38614 3409 38666 3415
rect 38722 800 38750 3631
rect 38818 800 38846 7627
rect 39970 7617 39998 18727
rect 40342 18267 40394 18273
rect 40342 18209 40394 18215
rect 40354 7765 40382 18209
rect 40342 7759 40394 7765
rect 40342 7701 40394 7707
rect 40246 7685 40298 7691
rect 40246 7627 40298 7633
rect 39958 7611 40010 7617
rect 39958 7553 40010 7559
rect 39478 7537 39530 7543
rect 39478 7479 39530 7485
rect 38902 6353 38954 6359
rect 38902 6295 38954 6301
rect 38914 800 38942 6295
rect 39190 6131 39242 6137
rect 39190 6073 39242 6079
rect 39094 5687 39146 5693
rect 39094 5629 39146 5635
rect 38998 4355 39050 4361
rect 38998 4297 39050 4303
rect 39010 800 39038 4297
rect 39106 2955 39134 5629
rect 39094 2949 39146 2955
rect 39094 2891 39146 2897
rect 39202 800 39230 6073
rect 39286 5687 39338 5693
rect 39286 5629 39338 5635
rect 39298 800 39326 5629
rect 39382 5021 39434 5027
rect 39382 4963 39434 4969
rect 39394 3843 39422 4963
rect 39382 3837 39434 3843
rect 39382 3779 39434 3785
rect 39382 3541 39434 3547
rect 39382 3483 39434 3489
rect 39394 800 39422 3483
rect 39490 800 39518 7479
rect 39862 6871 39914 6877
rect 39862 6813 39914 6819
rect 39766 4355 39818 4361
rect 39766 4297 39818 4303
rect 39670 3171 39722 3177
rect 39670 3113 39722 3119
rect 39682 800 39710 3113
rect 39778 800 39806 4297
rect 39874 800 39902 6813
rect 40150 5021 40202 5027
rect 40150 4963 40202 4969
rect 40054 4133 40106 4139
rect 40054 4075 40106 4081
rect 40066 800 40094 4075
rect 40162 3917 40190 4963
rect 40150 3911 40202 3917
rect 40150 3853 40202 3859
rect 40150 3467 40202 3473
rect 40150 3409 40202 3415
rect 40162 800 40190 3409
rect 40258 800 40286 7627
rect 41122 7173 41150 44035
rect 42082 33739 42110 56171
rect 42262 44093 42314 44099
rect 42262 44035 42314 44041
rect 42070 33733 42122 33739
rect 42070 33675 42122 33681
rect 41302 28923 41354 28929
rect 41302 28865 41354 28871
rect 41110 7167 41162 7173
rect 41110 7109 41162 7115
rect 41314 6433 41342 28865
rect 41494 14567 41546 14573
rect 41494 14509 41546 14515
rect 41506 7913 41534 14509
rect 42274 7913 42302 44035
rect 42370 15461 42398 56171
rect 42742 20117 42794 20123
rect 42742 20059 42794 20065
rect 42358 15455 42410 15461
rect 42358 15397 42410 15403
rect 41494 7907 41546 7913
rect 41494 7849 41546 7855
rect 42262 7907 42314 7913
rect 42262 7849 42314 7855
rect 41398 7759 41450 7765
rect 41398 7701 41450 7707
rect 41302 6427 41354 6433
rect 41302 6369 41354 6375
rect 40342 6353 40394 6359
rect 40342 6295 40394 6301
rect 40354 800 40382 6295
rect 40630 6205 40682 6211
rect 40630 6147 40682 6153
rect 40534 3023 40586 3029
rect 40534 2965 40586 2971
rect 40546 800 40574 2965
rect 40642 800 40670 6147
rect 40726 5687 40778 5693
rect 40726 5629 40778 5635
rect 40738 800 40766 5629
rect 40918 5021 40970 5027
rect 40918 4963 40970 4969
rect 40930 3177 40958 4963
rect 41302 3911 41354 3917
rect 41302 3853 41354 3859
rect 41014 3689 41066 3695
rect 41014 3631 41066 3637
rect 40918 3171 40970 3177
rect 40918 3113 40970 3119
rect 41026 1864 41054 3631
rect 41110 3171 41162 3177
rect 41110 3113 41162 3119
rect 40930 1836 41054 1864
rect 40930 800 40958 1836
rect 41014 1765 41066 1771
rect 41014 1707 41066 1713
rect 41026 800 41054 1707
rect 41122 800 41150 3113
rect 41206 3097 41258 3103
rect 41206 3039 41258 3045
rect 41218 800 41246 3039
rect 41314 1771 41342 3853
rect 41302 1765 41354 1771
rect 41302 1707 41354 1713
rect 41410 800 41438 7701
rect 41506 7617 41534 7849
rect 41494 7611 41546 7617
rect 41494 7553 41546 7559
rect 42454 7463 42506 7469
rect 42454 7405 42506 7411
rect 41494 7167 41546 7173
rect 41494 7109 41546 7115
rect 41506 3917 41534 7109
rect 42262 6945 42314 6951
rect 42262 6887 42314 6893
rect 41590 6871 41642 6877
rect 41590 6813 41642 6819
rect 41602 3936 41630 6813
rect 42274 6581 42302 6887
rect 42262 6575 42314 6581
rect 42262 6517 42314 6523
rect 41878 6353 41930 6359
rect 41878 6295 41930 6301
rect 41782 5687 41834 5693
rect 41782 5629 41834 5635
rect 41686 5021 41738 5027
rect 41686 4963 41738 4969
rect 41698 4139 41726 4963
rect 41686 4133 41738 4139
rect 41686 4075 41738 4081
rect 41494 3911 41546 3917
rect 41602 3908 41726 3936
rect 41494 3853 41546 3859
rect 41590 3615 41642 3621
rect 41590 3557 41642 3563
rect 41494 3245 41546 3251
rect 41494 3187 41546 3193
rect 41506 800 41534 3187
rect 41602 800 41630 3557
rect 41698 800 41726 3908
rect 41794 3251 41822 5629
rect 41782 3245 41834 3251
rect 41782 3187 41834 3193
rect 41780 3062 41836 3071
rect 41780 2997 41836 3006
rect 41794 2955 41822 2997
rect 41782 2949 41834 2955
rect 41782 2891 41834 2897
rect 41890 800 41918 6295
rect 42166 6205 42218 6211
rect 42166 6147 42218 6153
rect 42070 5021 42122 5027
rect 42070 4963 42122 4969
rect 41974 4355 42026 4361
rect 41974 4297 42026 4303
rect 41986 800 42014 4297
rect 42082 3177 42110 4963
rect 42070 3171 42122 3177
rect 42070 3113 42122 3119
rect 42178 3085 42206 6147
rect 42262 5687 42314 5693
rect 42262 5629 42314 5635
rect 42082 3057 42206 3085
rect 42082 800 42110 3057
rect 42274 800 42302 5629
rect 42358 4355 42410 4361
rect 42358 4297 42410 4303
rect 42370 800 42398 4297
rect 42466 800 42494 7405
rect 42754 5841 42782 20059
rect 42838 19229 42890 19235
rect 42838 19171 42890 19177
rect 42850 6433 42878 19171
rect 42946 17237 42974 56689
rect 43330 56531 43358 59200
rect 43906 56531 43934 59200
rect 44386 56975 44414 59200
rect 44374 56969 44426 56975
rect 44374 56911 44426 56917
rect 44962 56531 44990 59200
rect 43318 56525 43370 56531
rect 43318 56467 43370 56473
rect 43894 56525 43946 56531
rect 43894 56467 43946 56473
rect 44950 56525 45002 56531
rect 44950 56467 45002 56473
rect 43318 56377 43370 56383
rect 43318 56319 43370 56325
rect 43030 21449 43082 21455
rect 43030 21391 43082 21397
rect 42934 17231 42986 17237
rect 42934 17173 42986 17179
rect 43042 7099 43070 21391
rect 43030 7093 43082 7099
rect 43030 7035 43082 7041
rect 43030 6945 43082 6951
rect 42946 6905 43030 6933
rect 42838 6427 42890 6433
rect 42838 6369 42890 6375
rect 42742 5835 42794 5841
rect 42742 5777 42794 5783
rect 42742 3689 42794 3695
rect 42742 3631 42794 3637
rect 42550 3467 42602 3473
rect 42550 3409 42602 3415
rect 42562 800 42590 3409
rect 42754 800 42782 3631
rect 42946 3492 42974 6905
rect 43030 6887 43082 6893
rect 43222 5687 43274 5693
rect 43222 5629 43274 5635
rect 42850 3464 42974 3492
rect 42850 800 42878 3464
rect 43234 2900 43262 5629
rect 43330 3251 43358 56319
rect 43414 56229 43466 56235
rect 43414 56171 43466 56177
rect 43426 31001 43454 56171
rect 45442 55717 45470 59200
rect 45922 56901 45950 59200
rect 45910 56895 45962 56901
rect 45910 56837 45962 56843
rect 46102 56747 46154 56753
rect 46102 56689 46154 56695
rect 45430 55711 45482 55717
rect 45430 55653 45482 55659
rect 45238 55563 45290 55569
rect 45238 55505 45290 55511
rect 45250 55421 45278 55505
rect 45238 55415 45290 55421
rect 45238 55357 45290 55363
rect 44182 49421 44234 49427
rect 44182 49363 44234 49369
rect 44194 49205 44222 49363
rect 44182 49199 44234 49205
rect 44182 49141 44234 49147
rect 43894 36175 43946 36181
rect 43894 36117 43946 36123
rect 43414 30995 43466 31001
rect 43414 30937 43466 30943
rect 43798 20117 43850 20123
rect 43798 20059 43850 20065
rect 43606 7167 43658 7173
rect 43606 7109 43658 7115
rect 43510 5021 43562 5027
rect 43510 4963 43562 4969
rect 43414 4355 43466 4361
rect 43414 4297 43466 4303
rect 43426 3344 43454 4297
rect 43522 3473 43550 4963
rect 43510 3467 43562 3473
rect 43510 3409 43562 3415
rect 43426 3316 43550 3344
rect 43318 3245 43370 3251
rect 43318 3187 43370 3193
rect 43318 3023 43370 3029
rect 43318 2965 43370 2971
rect 42946 2872 43262 2900
rect 42946 800 42974 2872
rect 43330 1420 43358 2965
rect 43522 2160 43550 3316
rect 43234 1392 43358 1420
rect 43426 2132 43550 2160
rect 43030 951 43082 957
rect 43030 893 43082 899
rect 43042 800 43070 893
rect 43234 800 43262 1392
rect 43318 1321 43370 1327
rect 43318 1263 43370 1269
rect 43330 800 43358 1263
rect 43426 800 43454 2132
rect 43618 800 43646 7109
rect 43810 7099 43838 20059
rect 43906 17294 43934 36117
rect 44950 33585 45002 33591
rect 44950 33527 45002 33533
rect 44962 33147 44990 33527
rect 44950 33141 45002 33147
rect 44950 33083 45002 33089
rect 45142 30329 45194 30335
rect 45142 30271 45194 30277
rect 45046 29441 45098 29447
rect 45046 29383 45098 29389
rect 44086 23595 44138 23601
rect 44086 23537 44138 23543
rect 43906 17266 44030 17294
rect 43894 7463 43946 7469
rect 43894 7405 43946 7411
rect 43798 7093 43850 7099
rect 43798 7035 43850 7041
rect 43702 5687 43754 5693
rect 43702 5629 43754 5635
rect 43714 800 43742 5629
rect 43798 4207 43850 4213
rect 43798 4149 43850 4155
rect 43810 3917 43838 4149
rect 43798 3911 43850 3917
rect 43798 3853 43850 3859
rect 43798 3615 43850 3621
rect 43798 3557 43850 3563
rect 43810 800 43838 3557
rect 43906 800 43934 7405
rect 44002 6877 44030 17266
rect 44098 12974 44126 23537
rect 44950 22781 45002 22787
rect 44950 22723 45002 22729
rect 44758 21227 44810 21233
rect 44758 21169 44810 21175
rect 44098 12946 44222 12974
rect 44194 11687 44222 12946
rect 44086 11681 44138 11687
rect 44086 11623 44138 11629
rect 44182 11681 44234 11687
rect 44182 11623 44234 11629
rect 43990 6871 44042 6877
rect 43990 6813 44042 6819
rect 44098 6433 44126 11623
rect 44278 11607 44330 11613
rect 44278 11549 44330 11555
rect 44290 7691 44318 11549
rect 44374 8129 44426 8135
rect 44374 8071 44426 8077
rect 44278 7685 44330 7691
rect 44278 7627 44330 7633
rect 44278 7093 44330 7099
rect 44278 7035 44330 7041
rect 44086 6427 44138 6433
rect 44086 6369 44138 6375
rect 44182 6131 44234 6137
rect 44182 6073 44234 6079
rect 43990 3911 44042 3917
rect 43990 3853 44042 3859
rect 44002 1327 44030 3853
rect 44086 3837 44138 3843
rect 44086 3779 44138 3785
rect 43990 1321 44042 1327
rect 43990 1263 44042 1269
rect 44098 800 44126 3779
rect 44194 3251 44222 6073
rect 44182 3245 44234 3251
rect 44182 3187 44234 3193
rect 44182 3097 44234 3103
rect 44182 3039 44234 3045
rect 44194 800 44222 3039
rect 44290 800 44318 7035
rect 44386 7025 44414 8071
rect 44770 7765 44798 21169
rect 44854 20931 44906 20937
rect 44854 20873 44906 20879
rect 44866 20419 44894 20873
rect 44854 20413 44906 20419
rect 44854 20355 44906 20361
rect 44758 7759 44810 7765
rect 44758 7701 44810 7707
rect 44662 7463 44714 7469
rect 44662 7405 44714 7411
rect 44374 7019 44426 7025
rect 44374 6961 44426 6967
rect 44470 4281 44522 4287
rect 44470 4223 44522 4229
rect 44374 3171 44426 3177
rect 44374 3113 44426 3119
rect 44386 3071 44414 3113
rect 44372 3062 44428 3071
rect 44372 2997 44428 3006
rect 44374 2949 44426 2955
rect 44374 2891 44426 2897
rect 44386 957 44414 2891
rect 44374 951 44426 957
rect 44374 893 44426 899
rect 44482 800 44510 4223
rect 44566 3615 44618 3621
rect 44566 3557 44618 3563
rect 44578 800 44606 3557
rect 44674 800 44702 7405
rect 44962 6433 44990 22723
rect 45058 7913 45086 29383
rect 45046 7907 45098 7913
rect 45046 7849 45098 7855
rect 45046 7463 45098 7469
rect 45046 7405 45098 7411
rect 44950 6427 45002 6433
rect 44950 6369 45002 6375
rect 44758 5021 44810 5027
rect 44758 4963 44810 4969
rect 44770 3917 44798 4963
rect 44950 4355 45002 4361
rect 44950 4297 45002 4303
rect 44758 3911 44810 3917
rect 44758 3853 44810 3859
rect 44758 3541 44810 3547
rect 44758 3483 44810 3489
rect 44770 800 44798 3483
rect 44962 800 44990 4297
rect 45058 800 45086 7405
rect 45154 7099 45182 30271
rect 45250 16793 45278 55357
rect 45334 42095 45386 42101
rect 45334 42037 45386 42043
rect 45238 16787 45290 16793
rect 45238 16729 45290 16735
rect 45346 7617 45374 42037
rect 45430 36545 45482 36551
rect 45430 36487 45482 36493
rect 45442 7691 45470 36487
rect 45910 19599 45962 19605
rect 45910 19541 45962 19547
rect 45922 19161 45950 19541
rect 45910 19155 45962 19161
rect 45910 19097 45962 19103
rect 46114 18421 46142 56689
rect 46498 56531 46526 59200
rect 46486 56525 46538 56531
rect 46486 56467 46538 56473
rect 46870 56303 46922 56309
rect 46870 56245 46922 56251
rect 46678 56229 46730 56235
rect 46882 56217 46910 56245
rect 46730 56189 46910 56217
rect 46678 56171 46730 56177
rect 46486 55563 46538 55569
rect 46486 55505 46538 55511
rect 46498 55421 46526 55505
rect 46486 55415 46538 55421
rect 46486 55357 46538 55363
rect 46102 18415 46154 18421
rect 46102 18357 46154 18363
rect 46294 8943 46346 8949
rect 46294 8885 46346 8891
rect 46306 7765 46334 8885
rect 46294 7759 46346 7765
rect 46294 7701 46346 7707
rect 45430 7685 45482 7691
rect 45430 7627 45482 7633
rect 45334 7611 45386 7617
rect 45334 7553 45386 7559
rect 45814 7463 45866 7469
rect 45814 7405 45866 7411
rect 45142 7093 45194 7099
rect 45142 7035 45194 7041
rect 45718 6871 45770 6877
rect 45718 6813 45770 6819
rect 45526 6353 45578 6359
rect 45526 6295 45578 6301
rect 45142 5687 45194 5693
rect 45142 5629 45194 5635
rect 45154 4287 45182 5629
rect 45430 5021 45482 5027
rect 45430 4963 45482 4969
rect 45142 4281 45194 4287
rect 45142 4223 45194 4229
rect 45334 4133 45386 4139
rect 45334 4075 45386 4081
rect 45238 3763 45290 3769
rect 45238 3705 45290 3711
rect 45142 1099 45194 1105
rect 45142 1041 45194 1047
rect 45154 800 45182 1041
rect 45250 800 45278 3705
rect 45346 1105 45374 4075
rect 45442 3843 45470 4963
rect 45430 3837 45482 3843
rect 45430 3779 45482 3785
rect 45430 1469 45482 1475
rect 45430 1411 45482 1417
rect 45334 1099 45386 1105
rect 45334 1041 45386 1047
rect 45442 800 45470 1411
rect 45538 800 45566 6295
rect 45622 3023 45674 3029
rect 45622 2965 45674 2971
rect 45634 800 45662 2965
rect 45730 1475 45758 6813
rect 45718 1469 45770 1475
rect 45718 1411 45770 1417
rect 45826 800 45854 7405
rect 46498 6581 46526 55357
rect 46582 54749 46634 54755
rect 46582 54691 46634 54697
rect 46594 12974 46622 54691
rect 46690 17294 46718 56171
rect 46978 55717 47006 59200
rect 47554 56975 47582 59200
rect 47542 56969 47594 56975
rect 47542 56911 47594 56917
rect 47926 56821 47978 56827
rect 47926 56763 47978 56769
rect 47938 56235 47966 56763
rect 48034 56531 48062 59200
rect 48022 56525 48074 56531
rect 48022 56467 48074 56473
rect 47926 56229 47978 56235
rect 47926 56171 47978 56177
rect 48214 56229 48266 56235
rect 48214 56171 48266 56177
rect 46966 55711 47018 55717
rect 46966 55653 47018 55659
rect 47542 49495 47594 49501
rect 47542 49437 47594 49443
rect 47254 40097 47306 40103
rect 47254 40039 47306 40045
rect 47266 39881 47294 40039
rect 47254 39875 47306 39881
rect 47254 39817 47306 39823
rect 47350 37433 47402 37439
rect 47350 37375 47402 37381
rect 46690 17266 47102 17294
rect 47074 12974 47102 17266
rect 46594 12946 46718 12974
rect 47074 12946 47198 12974
rect 46582 7463 46634 7469
rect 46582 7405 46634 7411
rect 46486 6575 46538 6581
rect 46486 6517 46538 6523
rect 46102 5687 46154 5693
rect 46102 5629 46154 5635
rect 46114 4232 46142 5629
rect 46594 5120 46622 7405
rect 46690 6285 46718 12946
rect 47062 6945 47114 6951
rect 47062 6887 47114 6893
rect 46870 6871 46922 6877
rect 46870 6813 46922 6819
rect 46678 6279 46730 6285
rect 46678 6221 46730 6227
rect 46678 5687 46730 5693
rect 46678 5629 46730 5635
rect 46498 5092 46622 5120
rect 46198 5021 46250 5027
rect 46198 4963 46250 4969
rect 46294 5021 46346 5027
rect 46294 4963 46346 4969
rect 45922 4204 46142 4232
rect 45922 800 45950 4204
rect 46102 3837 46154 3843
rect 46102 3779 46154 3785
rect 46006 3615 46058 3621
rect 46006 3557 46058 3563
rect 46018 800 46046 3557
rect 46114 800 46142 3779
rect 46210 3547 46238 4963
rect 46306 4139 46334 4963
rect 46294 4133 46346 4139
rect 46294 4075 46346 4081
rect 46294 3911 46346 3917
rect 46294 3853 46346 3859
rect 46198 3541 46250 3547
rect 46198 3483 46250 3489
rect 46306 800 46334 3853
rect 46390 2949 46442 2955
rect 46390 2891 46442 2897
rect 46402 800 46430 2891
rect 46498 800 46526 5092
rect 46690 2894 46718 5629
rect 46774 4355 46826 4361
rect 46774 4297 46826 4303
rect 46594 2866 46718 2894
rect 46594 800 46622 2866
rect 46786 800 46814 4297
rect 46882 800 46910 6813
rect 46966 6353 47018 6359
rect 46966 6295 47018 6301
rect 46978 800 47006 6295
rect 47074 3843 47102 6887
rect 47170 4213 47198 12946
rect 47254 7463 47306 7469
rect 47254 7405 47306 7411
rect 47158 4207 47210 4213
rect 47158 4149 47210 4155
rect 47062 3837 47114 3843
rect 47062 3779 47114 3785
rect 47158 3689 47210 3695
rect 47158 3631 47210 3637
rect 47170 800 47198 3631
rect 47266 800 47294 7405
rect 47362 7099 47390 37375
rect 47554 7913 47582 49437
rect 48226 47059 48254 56171
rect 48610 56161 48638 59200
rect 49090 56901 49118 59200
rect 49078 56895 49130 56901
rect 49078 56837 49130 56843
rect 48694 56747 48746 56753
rect 48694 56689 48746 56695
rect 48598 56155 48650 56161
rect 48598 56097 48650 56103
rect 48214 47053 48266 47059
rect 48214 46995 48266 47001
rect 48598 35583 48650 35589
rect 48598 35525 48650 35531
rect 48214 9461 48266 9467
rect 48214 9403 48266 9409
rect 48226 9171 48254 9403
rect 48214 9165 48266 9171
rect 48214 9107 48266 9113
rect 48610 8579 48638 35525
rect 48706 19457 48734 56689
rect 49666 56531 49694 59200
rect 49942 56969 49994 56975
rect 49942 56911 49994 56917
rect 49654 56525 49706 56531
rect 49654 56467 49706 56473
rect 49174 56377 49226 56383
rect 49174 56319 49226 56325
rect 48886 56229 48938 56235
rect 48886 56171 48938 56177
rect 48790 45425 48842 45431
rect 48790 45367 48842 45373
rect 48802 45209 48830 45367
rect 48790 45203 48842 45209
rect 48790 45145 48842 45151
rect 48790 34103 48842 34109
rect 48790 34045 48842 34051
rect 48694 19451 48746 19457
rect 48694 19393 48746 19399
rect 48598 8573 48650 8579
rect 48598 8515 48650 8521
rect 48022 8277 48074 8283
rect 48022 8219 48074 8225
rect 47542 7907 47594 7913
rect 47542 7849 47594 7855
rect 47350 7093 47402 7099
rect 47350 7035 47402 7041
rect 47734 6353 47786 6359
rect 47734 6295 47786 6301
rect 47542 5687 47594 5693
rect 47542 5629 47594 5635
rect 47554 4380 47582 5629
rect 47638 5021 47690 5027
rect 47638 4963 47690 4969
rect 47362 4352 47582 4380
rect 47362 800 47390 4352
rect 47446 4281 47498 4287
rect 47446 4223 47498 4229
rect 47458 800 47486 4223
rect 47650 3917 47678 4963
rect 47638 3911 47690 3917
rect 47638 3853 47690 3859
rect 47638 3615 47690 3621
rect 47638 3557 47690 3563
rect 47650 800 47678 3557
rect 47746 800 47774 6295
rect 47830 4355 47882 4361
rect 47830 4297 47882 4303
rect 47842 800 47870 4297
rect 48034 800 48062 8219
rect 48694 8203 48746 8209
rect 48694 8145 48746 8151
rect 48310 7463 48362 7469
rect 48310 7405 48362 7411
rect 48118 4133 48170 4139
rect 48118 4075 48170 4081
rect 48130 800 48158 4075
rect 48214 3689 48266 3695
rect 48214 3631 48266 3637
rect 48226 800 48254 3631
rect 48322 800 48350 7405
rect 48406 6945 48458 6951
rect 48406 6887 48458 6893
rect 48418 3621 48446 6887
rect 48598 4281 48650 4287
rect 48598 4223 48650 4229
rect 48502 3911 48554 3917
rect 48502 3853 48554 3859
rect 48406 3615 48458 3621
rect 48406 3557 48458 3563
rect 48514 800 48542 3853
rect 48610 800 48638 4223
rect 48706 800 48734 8145
rect 48802 7173 48830 34045
rect 48898 18569 48926 56171
rect 49186 47503 49214 56319
rect 49654 56303 49706 56309
rect 49654 56245 49706 56251
rect 49174 47497 49226 47503
rect 49174 47439 49226 47445
rect 49558 43797 49610 43803
rect 49558 43739 49610 43745
rect 49462 39579 49514 39585
rect 49462 39521 49514 39527
rect 48886 18563 48938 18569
rect 48886 18505 48938 18511
rect 49366 16195 49418 16201
rect 49366 16137 49418 16143
rect 48982 15899 49034 15905
rect 48982 15841 49034 15847
rect 48886 8277 48938 8283
rect 48994 8265 49022 15841
rect 48938 8237 49022 8265
rect 48886 8219 48938 8225
rect 49378 7765 49406 16137
rect 49474 8376 49502 39521
rect 49570 8524 49598 43739
rect 49666 33221 49694 56245
rect 49846 56229 49898 56235
rect 49846 56171 49898 56177
rect 49750 54231 49802 54237
rect 49750 54173 49802 54179
rect 49654 33215 49706 33221
rect 49654 33157 49706 33163
rect 49654 27591 49706 27597
rect 49654 27533 49706 27539
rect 49666 8672 49694 27533
rect 49762 8875 49790 54173
rect 49858 36773 49886 56171
rect 49846 36767 49898 36773
rect 49846 36709 49898 36715
rect 49954 35737 49982 56911
rect 50146 56531 50174 59200
rect 50722 56901 50750 59200
rect 50710 56895 50762 56901
rect 50710 56837 50762 56843
rect 50806 56747 50858 56753
rect 50806 56689 50858 56695
rect 50348 56638 50644 56658
rect 50404 56636 50428 56638
rect 50484 56636 50508 56638
rect 50564 56636 50588 56638
rect 50426 56584 50428 56636
rect 50490 56584 50502 56636
rect 50564 56584 50566 56636
rect 50404 56582 50428 56584
rect 50484 56582 50508 56584
rect 50564 56582 50588 56584
rect 50348 56562 50644 56582
rect 50134 56525 50186 56531
rect 50134 56467 50186 56473
rect 50710 55415 50762 55421
rect 50710 55357 50762 55363
rect 50348 55306 50644 55326
rect 50404 55304 50428 55306
rect 50484 55304 50508 55306
rect 50564 55304 50588 55306
rect 50426 55252 50428 55304
rect 50490 55252 50502 55304
rect 50564 55252 50566 55304
rect 50404 55250 50428 55252
rect 50484 55250 50508 55252
rect 50564 55250 50588 55252
rect 50348 55230 50644 55250
rect 50348 53974 50644 53994
rect 50404 53972 50428 53974
rect 50484 53972 50508 53974
rect 50564 53972 50588 53974
rect 50426 53920 50428 53972
rect 50490 53920 50502 53972
rect 50564 53920 50566 53972
rect 50404 53918 50428 53920
rect 50484 53918 50508 53920
rect 50564 53918 50588 53920
rect 50348 53898 50644 53918
rect 50348 52642 50644 52662
rect 50404 52640 50428 52642
rect 50484 52640 50508 52642
rect 50564 52640 50588 52642
rect 50426 52588 50428 52640
rect 50490 52588 50502 52640
rect 50564 52588 50566 52640
rect 50404 52586 50428 52588
rect 50484 52586 50508 52588
rect 50564 52586 50588 52588
rect 50348 52566 50644 52586
rect 50348 51310 50644 51330
rect 50404 51308 50428 51310
rect 50484 51308 50508 51310
rect 50564 51308 50588 51310
rect 50426 51256 50428 51308
rect 50490 51256 50502 51308
rect 50564 51256 50566 51308
rect 50404 51254 50428 51256
rect 50484 51254 50508 51256
rect 50564 51254 50588 51256
rect 50348 51234 50644 51254
rect 50230 50753 50282 50759
rect 50230 50695 50282 50701
rect 49942 35731 49994 35737
rect 49942 35673 49994 35679
rect 49942 34251 49994 34257
rect 49942 34193 49994 34199
rect 49846 30773 49898 30779
rect 49846 30715 49898 30721
rect 49750 8869 49802 8875
rect 49750 8811 49802 8817
rect 49666 8644 49790 8672
rect 49570 8496 49694 8524
rect 49474 8348 49598 8376
rect 49462 8277 49514 8283
rect 49462 8219 49514 8225
rect 49366 7759 49418 7765
rect 49366 7701 49418 7707
rect 48790 7167 48842 7173
rect 48790 7109 48842 7115
rect 48790 6353 48842 6359
rect 48790 6295 48842 6301
rect 48802 800 48830 6295
rect 49078 5687 49130 5693
rect 49078 5629 49130 5635
rect 48982 4207 49034 4213
rect 48982 4149 49034 4155
rect 48994 800 49022 4149
rect 49090 4139 49118 5629
rect 49366 5021 49418 5027
rect 49366 4963 49418 4969
rect 49078 4133 49130 4139
rect 49078 4075 49130 4081
rect 49174 4133 49226 4139
rect 49174 4075 49226 4081
rect 49078 3837 49130 3843
rect 49078 3779 49130 3785
rect 49090 800 49118 3779
rect 49186 800 49214 4075
rect 49378 800 49406 4963
rect 49474 800 49502 8219
rect 49570 7913 49598 8348
rect 49558 7907 49610 7913
rect 49558 7849 49610 7855
rect 49666 6581 49694 8496
rect 49762 7691 49790 8644
rect 49858 8357 49886 30715
rect 49846 8351 49898 8357
rect 49846 8293 49898 8299
rect 49750 7685 49802 7691
rect 49750 7627 49802 7633
rect 49954 7173 49982 34193
rect 50242 17294 50270 50695
rect 50348 49978 50644 49998
rect 50404 49976 50428 49978
rect 50484 49976 50508 49978
rect 50564 49976 50588 49978
rect 50426 49924 50428 49976
rect 50490 49924 50502 49976
rect 50564 49924 50566 49976
rect 50404 49922 50428 49924
rect 50484 49922 50508 49924
rect 50564 49922 50588 49924
rect 50348 49902 50644 49922
rect 50348 48646 50644 48666
rect 50404 48644 50428 48646
rect 50484 48644 50508 48646
rect 50564 48644 50588 48646
rect 50426 48592 50428 48644
rect 50490 48592 50502 48644
rect 50564 48592 50566 48644
rect 50404 48590 50428 48592
rect 50484 48590 50508 48592
rect 50564 48590 50588 48592
rect 50348 48570 50644 48590
rect 50348 47314 50644 47334
rect 50404 47312 50428 47314
rect 50484 47312 50508 47314
rect 50564 47312 50588 47314
rect 50426 47260 50428 47312
rect 50490 47260 50502 47312
rect 50564 47260 50566 47312
rect 50404 47258 50428 47260
rect 50484 47258 50508 47260
rect 50564 47258 50588 47260
rect 50348 47238 50644 47258
rect 50348 45982 50644 46002
rect 50404 45980 50428 45982
rect 50484 45980 50508 45982
rect 50564 45980 50588 45982
rect 50426 45928 50428 45980
rect 50490 45928 50502 45980
rect 50564 45928 50566 45980
rect 50404 45926 50428 45928
rect 50484 45926 50508 45928
rect 50564 45926 50588 45928
rect 50348 45906 50644 45926
rect 50348 44650 50644 44670
rect 50404 44648 50428 44650
rect 50484 44648 50508 44650
rect 50564 44648 50588 44650
rect 50426 44596 50428 44648
rect 50490 44596 50502 44648
rect 50564 44596 50566 44648
rect 50404 44594 50428 44596
rect 50484 44594 50508 44596
rect 50564 44594 50588 44596
rect 50348 44574 50644 44594
rect 50348 43318 50644 43338
rect 50404 43316 50428 43318
rect 50484 43316 50508 43318
rect 50564 43316 50588 43318
rect 50426 43264 50428 43316
rect 50490 43264 50502 43316
rect 50564 43264 50566 43316
rect 50404 43262 50428 43264
rect 50484 43262 50508 43264
rect 50564 43262 50588 43264
rect 50348 43242 50644 43262
rect 50348 41986 50644 42006
rect 50404 41984 50428 41986
rect 50484 41984 50508 41986
rect 50564 41984 50588 41986
rect 50426 41932 50428 41984
rect 50490 41932 50502 41984
rect 50564 41932 50566 41984
rect 50404 41930 50428 41932
rect 50484 41930 50508 41932
rect 50564 41930 50588 41932
rect 50348 41910 50644 41930
rect 50348 40654 50644 40674
rect 50404 40652 50428 40654
rect 50484 40652 50508 40654
rect 50564 40652 50588 40654
rect 50426 40600 50428 40652
rect 50490 40600 50502 40652
rect 50564 40600 50566 40652
rect 50404 40598 50428 40600
rect 50484 40598 50508 40600
rect 50564 40598 50588 40600
rect 50348 40578 50644 40598
rect 50348 39322 50644 39342
rect 50404 39320 50428 39322
rect 50484 39320 50508 39322
rect 50564 39320 50588 39322
rect 50426 39268 50428 39320
rect 50490 39268 50502 39320
rect 50564 39268 50566 39320
rect 50404 39266 50428 39268
rect 50484 39266 50508 39268
rect 50564 39266 50588 39268
rect 50348 39246 50644 39266
rect 50348 37990 50644 38010
rect 50404 37988 50428 37990
rect 50484 37988 50508 37990
rect 50564 37988 50588 37990
rect 50426 37936 50428 37988
rect 50490 37936 50502 37988
rect 50564 37936 50566 37988
rect 50404 37934 50428 37936
rect 50484 37934 50508 37936
rect 50564 37934 50588 37936
rect 50348 37914 50644 37934
rect 50348 36658 50644 36678
rect 50404 36656 50428 36658
rect 50484 36656 50508 36658
rect 50564 36656 50588 36658
rect 50426 36604 50428 36656
rect 50490 36604 50502 36656
rect 50564 36604 50566 36656
rect 50404 36602 50428 36604
rect 50484 36602 50508 36604
rect 50564 36602 50588 36604
rect 50348 36582 50644 36602
rect 50348 35326 50644 35346
rect 50404 35324 50428 35326
rect 50484 35324 50508 35326
rect 50564 35324 50588 35326
rect 50426 35272 50428 35324
rect 50490 35272 50502 35324
rect 50564 35272 50566 35324
rect 50404 35270 50428 35272
rect 50484 35270 50508 35272
rect 50564 35270 50588 35272
rect 50348 35250 50644 35270
rect 50348 33994 50644 34014
rect 50404 33992 50428 33994
rect 50484 33992 50508 33994
rect 50564 33992 50588 33994
rect 50426 33940 50428 33992
rect 50490 33940 50502 33992
rect 50564 33940 50566 33992
rect 50404 33938 50428 33940
rect 50484 33938 50508 33940
rect 50564 33938 50588 33940
rect 50348 33918 50644 33938
rect 50348 32662 50644 32682
rect 50404 32660 50428 32662
rect 50484 32660 50508 32662
rect 50564 32660 50588 32662
rect 50426 32608 50428 32660
rect 50490 32608 50502 32660
rect 50564 32608 50566 32660
rect 50404 32606 50428 32608
rect 50484 32606 50508 32608
rect 50564 32606 50588 32608
rect 50348 32586 50644 32606
rect 50348 31330 50644 31350
rect 50404 31328 50428 31330
rect 50484 31328 50508 31330
rect 50564 31328 50588 31330
rect 50426 31276 50428 31328
rect 50490 31276 50502 31328
rect 50564 31276 50566 31328
rect 50404 31274 50428 31276
rect 50484 31274 50508 31276
rect 50564 31274 50588 31276
rect 50348 31254 50644 31274
rect 50348 29998 50644 30018
rect 50404 29996 50428 29998
rect 50484 29996 50508 29998
rect 50564 29996 50588 29998
rect 50426 29944 50428 29996
rect 50490 29944 50502 29996
rect 50564 29944 50566 29996
rect 50404 29942 50428 29944
rect 50484 29942 50508 29944
rect 50564 29942 50588 29944
rect 50348 29922 50644 29942
rect 50348 28666 50644 28686
rect 50404 28664 50428 28666
rect 50484 28664 50508 28666
rect 50564 28664 50588 28666
rect 50426 28612 50428 28664
rect 50490 28612 50502 28664
rect 50564 28612 50566 28664
rect 50404 28610 50428 28612
rect 50484 28610 50508 28612
rect 50564 28610 50588 28612
rect 50348 28590 50644 28610
rect 50348 27334 50644 27354
rect 50404 27332 50428 27334
rect 50484 27332 50508 27334
rect 50564 27332 50588 27334
rect 50426 27280 50428 27332
rect 50490 27280 50502 27332
rect 50564 27280 50566 27332
rect 50404 27278 50428 27280
rect 50484 27278 50508 27280
rect 50564 27278 50588 27280
rect 50348 27258 50644 27278
rect 50348 26002 50644 26022
rect 50404 26000 50428 26002
rect 50484 26000 50508 26002
rect 50564 26000 50588 26002
rect 50426 25948 50428 26000
rect 50490 25948 50502 26000
rect 50564 25948 50566 26000
rect 50404 25946 50428 25948
rect 50484 25946 50508 25948
rect 50564 25946 50588 25948
rect 50348 25926 50644 25946
rect 50348 24670 50644 24690
rect 50404 24668 50428 24670
rect 50484 24668 50508 24670
rect 50564 24668 50588 24670
rect 50426 24616 50428 24668
rect 50490 24616 50502 24668
rect 50564 24616 50566 24668
rect 50404 24614 50428 24616
rect 50484 24614 50508 24616
rect 50564 24614 50588 24616
rect 50348 24594 50644 24614
rect 50348 23338 50644 23358
rect 50404 23336 50428 23338
rect 50484 23336 50508 23338
rect 50564 23336 50588 23338
rect 50426 23284 50428 23336
rect 50490 23284 50502 23336
rect 50564 23284 50566 23336
rect 50404 23282 50428 23284
rect 50484 23282 50508 23284
rect 50564 23282 50588 23284
rect 50348 23262 50644 23282
rect 50348 22006 50644 22026
rect 50404 22004 50428 22006
rect 50484 22004 50508 22006
rect 50564 22004 50588 22006
rect 50426 21952 50428 22004
rect 50490 21952 50502 22004
rect 50564 21952 50566 22004
rect 50404 21950 50428 21952
rect 50484 21950 50508 21952
rect 50564 21950 50588 21952
rect 50348 21930 50644 21950
rect 50348 20674 50644 20694
rect 50404 20672 50428 20674
rect 50484 20672 50508 20674
rect 50564 20672 50588 20674
rect 50426 20620 50428 20672
rect 50490 20620 50502 20672
rect 50564 20620 50566 20672
rect 50404 20618 50428 20620
rect 50484 20618 50508 20620
rect 50564 20618 50588 20620
rect 50348 20598 50644 20618
rect 50348 19342 50644 19362
rect 50404 19340 50428 19342
rect 50484 19340 50508 19342
rect 50564 19340 50588 19342
rect 50426 19288 50428 19340
rect 50490 19288 50502 19340
rect 50564 19288 50566 19340
rect 50404 19286 50428 19288
rect 50484 19286 50508 19288
rect 50564 19286 50588 19288
rect 50348 19266 50644 19286
rect 50348 18010 50644 18030
rect 50404 18008 50428 18010
rect 50484 18008 50508 18010
rect 50564 18008 50588 18010
rect 50426 17956 50428 18008
rect 50490 17956 50502 18008
rect 50564 17956 50566 18008
rect 50404 17954 50428 17956
rect 50484 17954 50508 17956
rect 50564 17954 50588 17956
rect 50348 17934 50644 17954
rect 50146 17266 50270 17294
rect 50038 16121 50090 16127
rect 50038 16063 50090 16069
rect 50050 7765 50078 16063
rect 50146 8579 50174 17266
rect 50348 16678 50644 16698
rect 50404 16676 50428 16678
rect 50484 16676 50508 16678
rect 50564 16676 50588 16678
rect 50426 16624 50428 16676
rect 50490 16624 50502 16676
rect 50564 16624 50566 16676
rect 50404 16622 50428 16624
rect 50484 16622 50508 16624
rect 50564 16622 50588 16624
rect 50348 16602 50644 16622
rect 50348 15346 50644 15366
rect 50404 15344 50428 15346
rect 50484 15344 50508 15346
rect 50564 15344 50588 15346
rect 50426 15292 50428 15344
rect 50490 15292 50502 15344
rect 50564 15292 50566 15344
rect 50404 15290 50428 15292
rect 50484 15290 50508 15292
rect 50564 15290 50588 15292
rect 50348 15270 50644 15290
rect 50348 14014 50644 14034
rect 50404 14012 50428 14014
rect 50484 14012 50508 14014
rect 50564 14012 50588 14014
rect 50426 13960 50428 14012
rect 50490 13960 50502 14012
rect 50564 13960 50566 14012
rect 50404 13958 50428 13960
rect 50484 13958 50508 13960
rect 50564 13958 50588 13960
rect 50348 13938 50644 13958
rect 50348 12682 50644 12702
rect 50404 12680 50428 12682
rect 50484 12680 50508 12682
rect 50564 12680 50588 12682
rect 50426 12628 50428 12680
rect 50490 12628 50502 12680
rect 50564 12628 50566 12680
rect 50404 12626 50428 12628
rect 50484 12626 50508 12628
rect 50564 12626 50588 12628
rect 50348 12606 50644 12626
rect 50348 11350 50644 11370
rect 50404 11348 50428 11350
rect 50484 11348 50508 11350
rect 50564 11348 50588 11350
rect 50426 11296 50428 11348
rect 50490 11296 50502 11348
rect 50564 11296 50566 11348
rect 50404 11294 50428 11296
rect 50484 11294 50508 11296
rect 50564 11294 50588 11296
rect 50348 11274 50644 11294
rect 50348 10018 50644 10038
rect 50404 10016 50428 10018
rect 50484 10016 50508 10018
rect 50564 10016 50588 10018
rect 50426 9964 50428 10016
rect 50490 9964 50502 10016
rect 50564 9964 50566 10016
rect 50404 9962 50428 9964
rect 50484 9962 50508 9964
rect 50564 9962 50588 9964
rect 50348 9942 50644 9962
rect 50722 9541 50750 55357
rect 50818 19531 50846 56689
rect 51202 56161 51230 59200
rect 51190 56155 51242 56161
rect 51190 56097 51242 56103
rect 51778 55717 51806 59200
rect 52150 56969 52202 56975
rect 52150 56911 52202 56917
rect 52162 56383 52190 56911
rect 52258 56901 52286 59200
rect 52834 57614 52862 59200
rect 52834 57586 52958 57614
rect 52246 56895 52298 56901
rect 52246 56837 52298 56843
rect 52822 56747 52874 56753
rect 52822 56689 52874 56695
rect 52150 56377 52202 56383
rect 52150 56319 52202 56325
rect 51766 55711 51818 55717
rect 51766 55653 51818 55659
rect 51574 55415 51626 55421
rect 51574 55357 51626 55363
rect 51094 54823 51146 54829
rect 51094 54765 51146 54771
rect 50806 19525 50858 19531
rect 50806 19467 50858 19473
rect 50710 9535 50762 9541
rect 50710 9477 50762 9483
rect 50230 8869 50282 8875
rect 50230 8811 50282 8817
rect 50134 8573 50186 8579
rect 50134 8515 50186 8521
rect 50038 7759 50090 7765
rect 50038 7701 50090 7707
rect 50038 7463 50090 7469
rect 50038 7405 50090 7411
rect 49942 7167 49994 7173
rect 49942 7109 49994 7115
rect 49654 6575 49706 6581
rect 49654 6517 49706 6523
rect 49846 6427 49898 6433
rect 49846 6369 49898 6375
rect 49558 6353 49610 6359
rect 49558 6295 49610 6301
rect 49570 800 49598 6295
rect 49654 5687 49706 5693
rect 49654 5629 49706 5635
rect 49666 3917 49694 5629
rect 49654 3911 49706 3917
rect 49654 3853 49706 3859
rect 49654 3023 49706 3029
rect 49654 2965 49706 2971
rect 49666 800 49694 2965
rect 49858 800 49886 6369
rect 49942 4281 49994 4287
rect 49942 4223 49994 4229
rect 49954 800 49982 4223
rect 50050 3843 50078 7405
rect 50134 6871 50186 6877
rect 50134 6813 50186 6819
rect 50038 3837 50090 3843
rect 50038 3779 50090 3785
rect 50038 2875 50090 2881
rect 50038 2817 50090 2823
rect 50050 800 50078 2817
rect 50146 800 50174 6813
rect 50242 6803 50270 8811
rect 50348 8686 50644 8706
rect 50404 8684 50428 8686
rect 50484 8684 50508 8686
rect 50564 8684 50588 8686
rect 50426 8632 50428 8684
rect 50490 8632 50502 8684
rect 50564 8632 50566 8684
rect 50404 8630 50428 8632
rect 50484 8630 50508 8632
rect 50564 8630 50588 8632
rect 50348 8610 50644 8630
rect 50806 8129 50858 8135
rect 50806 8071 50858 8077
rect 50348 7354 50644 7374
rect 50404 7352 50428 7354
rect 50484 7352 50508 7354
rect 50564 7352 50588 7354
rect 50426 7300 50428 7352
rect 50490 7300 50502 7352
rect 50564 7300 50566 7352
rect 50404 7298 50428 7300
rect 50484 7298 50508 7300
rect 50564 7298 50588 7300
rect 50348 7278 50644 7298
rect 50422 6945 50474 6951
rect 50422 6887 50474 6893
rect 50230 6797 50282 6803
rect 50230 6739 50282 6745
rect 50434 6507 50462 6887
rect 50422 6501 50474 6507
rect 50422 6443 50474 6449
rect 50348 6022 50644 6042
rect 50404 6020 50428 6022
rect 50484 6020 50508 6022
rect 50564 6020 50588 6022
rect 50426 5968 50428 6020
rect 50490 5968 50502 6020
rect 50564 5968 50566 6020
rect 50404 5966 50428 5968
rect 50484 5966 50508 5968
rect 50564 5966 50588 5968
rect 50348 5946 50644 5966
rect 50710 5687 50762 5693
rect 50710 5629 50762 5635
rect 50422 5021 50474 5027
rect 50422 4963 50474 4969
rect 50434 4824 50462 4963
rect 50242 4796 50462 4824
rect 50242 2894 50270 4796
rect 50348 4690 50644 4710
rect 50404 4688 50428 4690
rect 50484 4688 50508 4690
rect 50564 4688 50588 4690
rect 50426 4636 50428 4688
rect 50490 4636 50502 4688
rect 50564 4636 50566 4688
rect 50404 4634 50428 4636
rect 50484 4634 50508 4636
rect 50564 4634 50588 4636
rect 50348 4614 50644 4634
rect 50722 4139 50750 5629
rect 50818 5619 50846 8071
rect 51106 6359 51134 54765
rect 51190 37507 51242 37513
rect 51190 37449 51242 37455
rect 51202 6951 51230 37449
rect 51586 36995 51614 55357
rect 52150 44093 52202 44099
rect 52150 44035 52202 44041
rect 51574 36989 51626 36995
rect 51574 36931 51626 36937
rect 51286 36249 51338 36255
rect 51286 36191 51338 36197
rect 51190 6945 51242 6951
rect 51190 6887 51242 6893
rect 51298 6581 51326 36191
rect 52054 19599 52106 19605
rect 52054 19541 52106 19547
rect 51670 7463 51722 7469
rect 51670 7405 51722 7411
rect 51574 6945 51626 6951
rect 51574 6887 51626 6893
rect 51286 6575 51338 6581
rect 51286 6517 51338 6523
rect 51094 6353 51146 6359
rect 51094 6295 51146 6301
rect 51478 6205 51530 6211
rect 51478 6147 51530 6153
rect 51094 6131 51146 6137
rect 51094 6073 51146 6079
rect 50806 5613 50858 5619
rect 50806 5555 50858 5561
rect 50902 5021 50954 5027
rect 50902 4963 50954 4969
rect 50710 4133 50762 4139
rect 50710 4075 50762 4081
rect 50710 3689 50762 3695
rect 50710 3631 50762 3637
rect 50806 3689 50858 3695
rect 50806 3631 50858 3637
rect 50348 3358 50644 3378
rect 50404 3356 50428 3358
rect 50484 3356 50508 3358
rect 50564 3356 50588 3358
rect 50426 3304 50428 3356
rect 50490 3304 50502 3356
rect 50564 3304 50566 3356
rect 50404 3302 50428 3304
rect 50484 3302 50508 3304
rect 50564 3302 50588 3304
rect 50348 3282 50644 3302
rect 50722 2894 50750 3631
rect 50242 2866 50366 2894
rect 50338 800 50366 2866
rect 50434 2866 50750 2894
rect 50434 800 50462 2866
rect 50518 1543 50570 1549
rect 50518 1485 50570 1491
rect 50530 800 50558 1485
rect 50710 1469 50762 1475
rect 50710 1411 50762 1417
rect 50722 800 50750 1411
rect 50818 800 50846 3631
rect 50914 1475 50942 4963
rect 50998 4281 51050 4287
rect 50998 4223 51050 4229
rect 50902 1469 50954 1475
rect 50902 1411 50954 1417
rect 50902 1321 50954 1327
rect 50902 1263 50954 1269
rect 50914 800 50942 1263
rect 51010 800 51038 4223
rect 51106 1549 51134 6073
rect 51382 3911 51434 3917
rect 51382 3853 51434 3859
rect 51286 3689 51338 3695
rect 51202 3649 51286 3677
rect 51094 1543 51146 1549
rect 51094 1485 51146 1491
rect 51202 800 51230 3649
rect 51286 3631 51338 3637
rect 51286 3541 51338 3547
rect 51286 3483 51338 3489
rect 51298 800 51326 3483
rect 51394 800 51422 3853
rect 51490 3344 51518 6147
rect 51586 3547 51614 6887
rect 51574 3541 51626 3547
rect 51574 3483 51626 3489
rect 51490 3316 51614 3344
rect 51478 3023 51530 3029
rect 51478 2965 51530 2971
rect 51490 800 51518 2965
rect 51586 1327 51614 3316
rect 51574 1321 51626 1327
rect 51574 1263 51626 1269
rect 51682 800 51710 7405
rect 52066 7099 52094 19541
rect 52162 8209 52190 44035
rect 52534 42761 52586 42767
rect 52534 42703 52586 42709
rect 52150 8203 52202 8209
rect 52150 8145 52202 8151
rect 52342 7463 52394 7469
rect 52342 7405 52394 7411
rect 52054 7093 52106 7099
rect 52054 7035 52106 7041
rect 52246 6871 52298 6877
rect 52246 6813 52298 6819
rect 52150 5687 52202 5693
rect 52150 5629 52202 5635
rect 51862 5021 51914 5027
rect 51862 4963 51914 4969
rect 51958 5021 52010 5027
rect 51958 4963 52010 4969
rect 51874 3917 51902 4963
rect 51862 3911 51914 3917
rect 51862 3853 51914 3859
rect 51970 3788 51998 4963
rect 51778 3760 51998 3788
rect 51778 800 51806 3760
rect 52054 3689 52106 3695
rect 51970 3649 52054 3677
rect 51970 976 51998 3649
rect 52054 3631 52106 3637
rect 52054 3541 52106 3547
rect 52054 3483 52106 3489
rect 51874 948 51998 976
rect 51874 800 51902 948
rect 52066 800 52094 3483
rect 52162 800 52190 5629
rect 52258 3547 52286 6813
rect 52246 3541 52298 3547
rect 52246 3483 52298 3489
rect 52246 2949 52298 2955
rect 52246 2891 52298 2897
rect 52258 800 52286 2891
rect 52354 800 52382 7405
rect 52546 7025 52574 42703
rect 52834 19901 52862 56689
rect 52930 56531 52958 57586
rect 53314 56531 53342 59200
rect 53890 56975 53918 59200
rect 53878 56969 53930 56975
rect 53878 56911 53930 56917
rect 54370 56531 54398 59200
rect 54838 56821 54890 56827
rect 54838 56763 54890 56769
rect 52918 56525 52970 56531
rect 52918 56467 52970 56473
rect 53302 56525 53354 56531
rect 53302 56467 53354 56473
rect 54358 56525 54410 56531
rect 54358 56467 54410 56473
rect 54358 56303 54410 56309
rect 54358 56245 54410 56251
rect 53014 56229 53066 56235
rect 53014 56171 53066 56177
rect 53398 56229 53450 56235
rect 53398 56171 53450 56177
rect 52918 39579 52970 39585
rect 52918 39521 52970 39527
rect 52822 19895 52874 19901
rect 52822 19837 52874 19843
rect 52930 8579 52958 39521
rect 53026 30927 53054 56171
rect 53014 30921 53066 30927
rect 53014 30863 53066 30869
rect 53410 20937 53438 56171
rect 54370 55051 54398 56245
rect 54454 56229 54506 56235
rect 54454 56171 54506 56177
rect 54358 55045 54410 55051
rect 54358 54987 54410 54993
rect 53398 20931 53450 20937
rect 53398 20873 53450 20879
rect 53398 14493 53450 14499
rect 53398 14435 53450 14441
rect 53410 9097 53438 14435
rect 53590 13531 53642 13537
rect 53590 13473 53642 13479
rect 53398 9091 53450 9097
rect 53398 9033 53450 9039
rect 52918 8573 52970 8579
rect 52918 8515 52970 8521
rect 53110 8277 53162 8283
rect 53110 8219 53162 8225
rect 53494 8277 53546 8283
rect 53494 8219 53546 8225
rect 52822 7611 52874 7617
rect 52822 7553 52874 7559
rect 52726 7463 52778 7469
rect 52726 7405 52778 7411
rect 52534 7019 52586 7025
rect 52534 6961 52586 6967
rect 52438 6279 52490 6285
rect 52438 6221 52490 6227
rect 52450 3103 52478 6221
rect 52534 5687 52586 5693
rect 52534 5629 52586 5635
rect 52438 3097 52490 3103
rect 52438 3039 52490 3045
rect 52546 800 52574 5629
rect 52630 4355 52682 4361
rect 52630 4297 52682 4303
rect 52642 800 52670 4297
rect 52738 800 52766 7405
rect 52834 2807 52862 7553
rect 53014 4281 53066 4287
rect 53014 4223 53066 4229
rect 52918 2949 52970 2955
rect 52918 2891 52970 2897
rect 52822 2801 52874 2807
rect 52822 2743 52874 2749
rect 52930 800 52958 2891
rect 53026 800 53054 4223
rect 53122 800 53150 8219
rect 53302 5021 53354 5027
rect 53302 4963 53354 4969
rect 53314 2900 53342 4963
rect 53398 3689 53450 3695
rect 53398 3631 53450 3637
rect 53218 2872 53342 2900
rect 53218 800 53246 2872
rect 53410 800 53438 3631
rect 53506 800 53534 8219
rect 53602 7765 53630 13473
rect 54466 10873 54494 56171
rect 54850 50537 54878 56763
rect 54946 56531 54974 59200
rect 55426 56901 55454 59200
rect 55414 56895 55466 56901
rect 55414 56837 55466 56843
rect 55414 56747 55466 56753
rect 55414 56689 55466 56695
rect 54934 56525 54986 56531
rect 54934 56467 54986 56473
rect 54838 50531 54890 50537
rect 54838 50473 54890 50479
rect 54646 46165 54698 46171
rect 54646 46107 54698 46113
rect 54454 10867 54506 10873
rect 54454 10809 54506 10815
rect 54658 9911 54686 46107
rect 55426 21529 55454 56689
rect 56002 56531 56030 59200
rect 55990 56525 56042 56531
rect 55990 56467 56042 56473
rect 55510 56229 55562 56235
rect 55510 56171 55562 56177
rect 55414 21523 55466 21529
rect 55414 21465 55466 21471
rect 55522 19679 55550 56171
rect 56482 55717 56510 59200
rect 57058 56901 57086 59200
rect 57046 56895 57098 56901
rect 57046 56837 57098 56843
rect 56758 56747 56810 56753
rect 56758 56689 56810 56695
rect 56770 56457 56798 56689
rect 56758 56451 56810 56457
rect 56758 56393 56810 56399
rect 57538 55717 57566 59200
rect 56470 55711 56522 55717
rect 56470 55653 56522 55659
rect 57526 55711 57578 55717
rect 57526 55653 57578 55659
rect 56662 55563 56714 55569
rect 56662 55505 56714 55511
rect 57526 55563 57578 55569
rect 57526 55505 57578 55511
rect 55606 55415 55658 55421
rect 55606 55357 55658 55363
rect 55618 55125 55646 55357
rect 55606 55119 55658 55125
rect 55606 55061 55658 55067
rect 55606 45425 55658 45431
rect 55606 45367 55658 45373
rect 55510 19673 55562 19679
rect 55510 19615 55562 19621
rect 54742 19599 54794 19605
rect 54742 19541 54794 19547
rect 54754 19235 54782 19541
rect 54742 19229 54794 19235
rect 54742 19171 54794 19177
rect 55618 9911 55646 45367
rect 56086 43649 56138 43655
rect 56086 43591 56138 43597
rect 56098 10577 56126 43591
rect 56674 13241 56702 55505
rect 57334 53417 57386 53423
rect 57334 53359 57386 53365
rect 56950 47867 57002 47873
rect 56950 47809 57002 47815
rect 56662 13235 56714 13241
rect 56662 13177 56714 13183
rect 56962 11243 56990 47809
rect 57346 12575 57374 53359
rect 57538 17294 57566 55505
rect 57910 54897 57962 54903
rect 57910 54839 57962 54845
rect 57622 54083 57674 54089
rect 57622 54025 57674 54031
rect 57442 17266 57566 17294
rect 57634 17294 57662 54025
rect 57718 53417 57770 53423
rect 57718 53359 57770 53365
rect 57730 20789 57758 53359
rect 57922 51055 57950 54839
rect 58114 54385 58142 59200
rect 58594 56309 58622 59200
rect 58582 56303 58634 56309
rect 58582 56245 58634 56251
rect 59170 55199 59198 59200
rect 59158 55193 59210 55199
rect 59158 55135 59210 55141
rect 58102 54379 58154 54385
rect 58102 54321 58154 54327
rect 59650 53867 59678 59200
rect 59638 53861 59690 53867
rect 59638 53803 59690 53809
rect 57910 51049 57962 51055
rect 57910 50991 57962 50997
rect 57718 20783 57770 20789
rect 57718 20725 57770 20731
rect 57634 17266 57758 17294
rect 57334 12569 57386 12575
rect 57334 12511 57386 12517
rect 57142 11755 57194 11761
rect 57142 11697 57194 11703
rect 56950 11237 57002 11243
rect 56950 11179 57002 11185
rect 56374 10941 56426 10947
rect 56374 10883 56426 10889
rect 56758 10941 56810 10947
rect 56758 10883 56810 10889
rect 56086 10571 56138 10577
rect 56086 10513 56138 10519
rect 55702 10127 55754 10133
rect 55702 10069 55754 10075
rect 56086 10127 56138 10133
rect 56086 10069 56138 10075
rect 54646 9905 54698 9911
rect 54646 9847 54698 9853
rect 55606 9905 55658 9911
rect 55606 9847 55658 9853
rect 54262 9609 54314 9615
rect 54262 9551 54314 9557
rect 55510 9609 55562 9615
rect 55510 9551 55562 9557
rect 53878 8795 53930 8801
rect 53878 8737 53930 8743
rect 53590 7759 53642 7765
rect 53590 7701 53642 7707
rect 53686 5687 53738 5693
rect 53686 5629 53738 5635
rect 53590 5613 53642 5619
rect 53590 5555 53642 5561
rect 53602 800 53630 5555
rect 53698 2955 53726 5629
rect 53782 3023 53834 3029
rect 53782 2965 53834 2971
rect 53686 2949 53738 2955
rect 53686 2891 53738 2897
rect 53794 1568 53822 2965
rect 53698 1540 53822 1568
rect 53698 800 53726 1540
rect 53890 800 53918 8737
rect 53974 6353 54026 6359
rect 53974 6295 54026 6301
rect 53986 800 54014 6295
rect 54070 4355 54122 4361
rect 54070 4297 54122 4303
rect 54082 800 54110 4297
rect 54274 800 54302 9551
rect 54934 9535 54986 9541
rect 54934 9477 54986 9483
rect 54550 8869 54602 8875
rect 54550 8811 54602 8817
rect 54358 3615 54410 3621
rect 54358 3557 54410 3563
rect 54370 1864 54398 3557
rect 54454 2801 54506 2807
rect 54454 2743 54506 2749
rect 54466 2511 54494 2743
rect 54454 2505 54506 2511
rect 54454 2447 54506 2453
rect 54370 1836 54494 1864
rect 54358 1765 54410 1771
rect 54358 1707 54410 1713
rect 54370 800 54398 1707
rect 54466 800 54494 1836
rect 54562 800 54590 8811
rect 54742 7019 54794 7025
rect 54742 6961 54794 6967
rect 54646 6353 54698 6359
rect 54646 6295 54698 6301
rect 54658 1771 54686 6295
rect 54646 1765 54698 1771
rect 54646 1707 54698 1713
rect 54754 800 54782 6961
rect 54838 2949 54890 2955
rect 54838 2891 54890 2897
rect 54850 800 54878 2891
rect 54946 800 54974 9477
rect 55414 7019 55466 7025
rect 55414 6961 55466 6967
rect 55030 6279 55082 6285
rect 55030 6221 55082 6227
rect 55042 800 55070 6221
rect 55318 3689 55370 3695
rect 55318 3631 55370 3637
rect 55330 3344 55358 3631
rect 55234 3316 55358 3344
rect 55234 800 55262 3316
rect 55318 3245 55370 3251
rect 55318 3187 55370 3193
rect 55330 800 55358 3187
rect 55426 800 55454 6961
rect 55522 3251 55550 9551
rect 55606 4355 55658 4361
rect 55606 4297 55658 4303
rect 55510 3245 55562 3251
rect 55510 3187 55562 3193
rect 55618 800 55646 4297
rect 55714 800 55742 10069
rect 55990 8943 56042 8949
rect 55990 8885 56042 8891
rect 55798 7685 55850 7691
rect 55798 7627 55850 7633
rect 55810 800 55838 7627
rect 56002 3917 56030 8885
rect 55990 3911 56042 3917
rect 55990 3853 56042 3859
rect 55894 3615 55946 3621
rect 55894 3557 55946 3563
rect 55906 800 55934 3557
rect 56098 800 56126 10069
rect 56182 7685 56234 7691
rect 56182 7627 56234 7633
rect 56194 800 56222 7627
rect 56278 6205 56330 6211
rect 56278 6147 56330 6153
rect 56290 4139 56318 6147
rect 56386 4213 56414 10883
rect 56470 10423 56522 10429
rect 56470 10365 56522 10371
rect 56374 4207 56426 4213
rect 56374 4149 56426 4155
rect 56278 4133 56330 4139
rect 56278 4075 56330 4081
rect 56278 3541 56330 3547
rect 56278 3483 56330 3489
rect 56290 800 56318 3483
rect 56482 800 56510 10365
rect 56662 7685 56714 7691
rect 56662 7627 56714 7633
rect 56674 5268 56702 7627
rect 56578 5240 56702 5268
rect 56578 800 56606 5240
rect 56662 4355 56714 4361
rect 56662 4297 56714 4303
rect 56674 800 56702 4297
rect 56770 800 56798 10883
rect 56854 9017 56906 9023
rect 56854 8959 56906 8965
rect 56866 4287 56894 8959
rect 56950 8351 57002 8357
rect 56950 8293 57002 8299
rect 56854 4281 56906 4287
rect 56854 4223 56906 4229
rect 56962 800 56990 8293
rect 57046 6945 57098 6951
rect 57046 6887 57098 6893
rect 57058 5841 57086 6887
rect 57046 5835 57098 5841
rect 57046 5777 57098 5783
rect 57046 5021 57098 5027
rect 57046 4963 57098 4969
rect 57058 800 57086 4963
rect 57154 800 57182 11697
rect 57238 9017 57290 9023
rect 57238 8959 57290 8965
rect 57250 800 57278 8959
rect 57442 5860 57470 17266
rect 57730 12974 57758 17266
rect 57730 12946 58238 12974
rect 57526 12273 57578 12279
rect 57526 12215 57578 12221
rect 57346 5832 57470 5860
rect 57346 4583 57374 5832
rect 57430 5687 57482 5693
rect 57430 5629 57482 5635
rect 57334 4577 57386 4583
rect 57334 4519 57386 4525
rect 57442 800 57470 5629
rect 57538 800 57566 12215
rect 57622 9683 57674 9689
rect 57622 9625 57674 9631
rect 57634 800 57662 9625
rect 58102 6353 58154 6359
rect 58102 6295 58154 6301
rect 57718 5835 57770 5841
rect 57718 5777 57770 5783
rect 57730 3177 57758 5777
rect 57814 4947 57866 4953
rect 57814 4889 57866 4895
rect 57718 3171 57770 3177
rect 57718 3113 57770 3119
rect 57826 800 57854 4889
rect 58006 4133 58058 4139
rect 58006 4075 58058 4081
rect 57910 3911 57962 3917
rect 57910 3853 57962 3859
rect 57922 800 57950 3853
rect 58018 800 58046 4075
rect 58114 800 58142 6295
rect 58210 3251 58238 12946
rect 59734 11829 59786 11835
rect 59734 11771 59786 11777
rect 58582 10201 58634 10207
rect 58582 10143 58634 10149
rect 58390 8277 58442 8283
rect 58390 8219 58442 8225
rect 58294 4207 58346 4213
rect 58294 4149 58346 4155
rect 58198 3245 58250 3251
rect 58198 3187 58250 3193
rect 58306 800 58334 4149
rect 58402 800 58430 8219
rect 58486 7019 58538 7025
rect 58486 6961 58538 6967
rect 58498 800 58526 6961
rect 58594 800 58622 10143
rect 58966 8129 59018 8135
rect 58966 8071 59018 8077
rect 58774 7611 58826 7617
rect 58774 7553 58826 7559
rect 58786 800 58814 7553
rect 58870 6279 58922 6285
rect 58870 6221 58922 6227
rect 58882 800 58910 6221
rect 58978 800 59006 8071
rect 59350 7833 59402 7839
rect 59350 7775 59402 7781
rect 59254 4873 59306 4879
rect 59254 4815 59306 4821
rect 59158 4281 59210 4287
rect 59158 4223 59210 4229
rect 59170 800 59198 4223
rect 59266 800 59294 4815
rect 59362 800 59390 7775
rect 59638 5613 59690 5619
rect 59638 5555 59690 5561
rect 59446 3171 59498 3177
rect 59446 3113 59498 3119
rect 59458 800 59486 3113
rect 59650 800 59678 5555
rect 59746 800 59774 11771
rect 59830 8203 59882 8209
rect 59830 8145 59882 8151
rect 59842 800 59870 8145
rect 20 0 76 800
rect 116 0 172 800
rect 212 0 268 800
rect 308 0 364 800
rect 500 0 556 800
rect 596 0 652 800
rect 692 0 748 800
rect 788 0 844 800
rect 980 0 1036 800
rect 1076 0 1132 800
rect 1172 0 1228 800
rect 1364 0 1420 800
rect 1460 0 1516 800
rect 1556 0 1612 800
rect 1652 0 1708 800
rect 1844 0 1900 800
rect 1940 0 1996 800
rect 2036 0 2092 800
rect 2132 0 2188 800
rect 2324 0 2380 800
rect 2420 0 2476 800
rect 2516 0 2572 800
rect 2708 0 2764 800
rect 2804 0 2860 800
rect 2900 0 2956 800
rect 2996 0 3052 800
rect 3188 0 3244 800
rect 3284 0 3340 800
rect 3380 0 3436 800
rect 3476 0 3532 800
rect 3668 0 3724 800
rect 3764 0 3820 800
rect 3860 0 3916 800
rect 4052 0 4108 800
rect 4148 0 4204 800
rect 4244 0 4300 800
rect 4340 0 4396 800
rect 4532 0 4588 800
rect 4628 0 4684 800
rect 4724 0 4780 800
rect 4916 0 4972 800
rect 5012 0 5068 800
rect 5108 0 5164 800
rect 5204 0 5260 800
rect 5396 0 5452 800
rect 5492 0 5548 800
rect 5588 0 5644 800
rect 5684 0 5740 800
rect 5876 0 5932 800
rect 5972 0 6028 800
rect 6068 0 6124 800
rect 6260 0 6316 800
rect 6356 0 6412 800
rect 6452 0 6508 800
rect 6548 0 6604 800
rect 6740 0 6796 800
rect 6836 0 6892 800
rect 6932 0 6988 800
rect 7028 0 7084 800
rect 7220 0 7276 800
rect 7316 0 7372 800
rect 7412 0 7468 800
rect 7604 0 7660 800
rect 7700 0 7756 800
rect 7796 0 7852 800
rect 7892 0 7948 800
rect 8084 0 8140 800
rect 8180 0 8236 800
rect 8276 0 8332 800
rect 8468 0 8524 800
rect 8564 0 8620 800
rect 8660 0 8716 800
rect 8756 0 8812 800
rect 8948 0 9004 800
rect 9044 0 9100 800
rect 9140 0 9196 800
rect 9236 0 9292 800
rect 9428 0 9484 800
rect 9524 0 9580 800
rect 9620 0 9676 800
rect 9812 0 9868 800
rect 9908 0 9964 800
rect 10004 0 10060 800
rect 10100 0 10156 800
rect 10292 0 10348 800
rect 10388 0 10444 800
rect 10484 0 10540 800
rect 10580 0 10636 800
rect 10772 0 10828 800
rect 10868 0 10924 800
rect 10964 0 11020 800
rect 11156 0 11212 800
rect 11252 0 11308 800
rect 11348 0 11404 800
rect 11444 0 11500 800
rect 11636 0 11692 800
rect 11732 0 11788 800
rect 11828 0 11884 800
rect 12020 0 12076 800
rect 12116 0 12172 800
rect 12212 0 12268 800
rect 12308 0 12364 800
rect 12500 0 12556 800
rect 12596 0 12652 800
rect 12692 0 12748 800
rect 12788 0 12844 800
rect 12980 0 13036 800
rect 13076 0 13132 800
rect 13172 0 13228 800
rect 13364 0 13420 800
rect 13460 0 13516 800
rect 13556 0 13612 800
rect 13652 0 13708 800
rect 13844 0 13900 800
rect 13940 0 13996 800
rect 14036 0 14092 800
rect 14132 0 14188 800
rect 14324 0 14380 800
rect 14420 0 14476 800
rect 14516 0 14572 800
rect 14708 0 14764 800
rect 14804 0 14860 800
rect 14900 0 14956 800
rect 14996 0 15052 800
rect 15188 0 15244 800
rect 15284 0 15340 800
rect 15380 0 15436 800
rect 15476 0 15532 800
rect 15668 0 15724 800
rect 15764 0 15820 800
rect 15860 0 15916 800
rect 16052 0 16108 800
rect 16148 0 16204 800
rect 16244 0 16300 800
rect 16340 0 16396 800
rect 16532 0 16588 800
rect 16628 0 16684 800
rect 16724 0 16780 800
rect 16916 0 16972 800
rect 17012 0 17068 800
rect 17108 0 17164 800
rect 17204 0 17260 800
rect 17396 0 17452 800
rect 17492 0 17548 800
rect 17588 0 17644 800
rect 17684 0 17740 800
rect 17876 0 17932 800
rect 17972 0 18028 800
rect 18068 0 18124 800
rect 18260 0 18316 800
rect 18356 0 18412 800
rect 18452 0 18508 800
rect 18548 0 18604 800
rect 18740 0 18796 800
rect 18836 0 18892 800
rect 18932 0 18988 800
rect 19028 0 19084 800
rect 19220 0 19276 800
rect 19316 0 19372 800
rect 19412 0 19468 800
rect 19604 0 19660 800
rect 19700 0 19756 800
rect 19796 0 19852 800
rect 19892 0 19948 800
rect 20084 0 20140 800
rect 20180 0 20236 800
rect 20276 0 20332 800
rect 20468 0 20524 800
rect 20564 0 20620 800
rect 20660 0 20716 800
rect 20756 0 20812 800
rect 20948 0 21004 800
rect 21044 0 21100 800
rect 21140 0 21196 800
rect 21236 0 21292 800
rect 21428 0 21484 800
rect 21524 0 21580 800
rect 21620 0 21676 800
rect 21812 0 21868 800
rect 21908 0 21964 800
rect 22004 0 22060 800
rect 22100 0 22156 800
rect 22292 0 22348 800
rect 22388 0 22444 800
rect 22484 0 22540 800
rect 22580 0 22636 800
rect 22772 0 22828 800
rect 22868 0 22924 800
rect 22964 0 23020 800
rect 23156 0 23212 800
rect 23252 0 23308 800
rect 23348 0 23404 800
rect 23444 0 23500 800
rect 23636 0 23692 800
rect 23732 0 23788 800
rect 23828 0 23884 800
rect 24020 0 24076 800
rect 24116 0 24172 800
rect 24212 0 24268 800
rect 24308 0 24364 800
rect 24500 0 24556 800
rect 24596 0 24652 800
rect 24692 0 24748 800
rect 24788 0 24844 800
rect 24980 0 25036 800
rect 25076 0 25132 800
rect 25172 0 25228 800
rect 25364 0 25420 800
rect 25460 0 25516 800
rect 25556 0 25612 800
rect 25652 0 25708 800
rect 25844 0 25900 800
rect 25940 0 25996 800
rect 26036 0 26092 800
rect 26132 0 26188 800
rect 26324 0 26380 800
rect 26420 0 26476 800
rect 26516 0 26572 800
rect 26708 0 26764 800
rect 26804 0 26860 800
rect 26900 0 26956 800
rect 26996 0 27052 800
rect 27188 0 27244 800
rect 27284 0 27340 800
rect 27380 0 27436 800
rect 27476 0 27532 800
rect 27668 0 27724 800
rect 27764 0 27820 800
rect 27860 0 27916 800
rect 28052 0 28108 800
rect 28148 0 28204 800
rect 28244 0 28300 800
rect 28340 0 28396 800
rect 28532 0 28588 800
rect 28628 0 28684 800
rect 28724 0 28780 800
rect 28916 0 28972 800
rect 29012 0 29068 800
rect 29108 0 29164 800
rect 29204 0 29260 800
rect 29396 0 29452 800
rect 29492 0 29548 800
rect 29588 0 29644 800
rect 29684 0 29740 800
rect 29876 0 29932 800
rect 29972 0 30028 800
rect 30068 0 30124 800
rect 30260 0 30316 800
rect 30356 0 30412 800
rect 30452 0 30508 800
rect 30548 0 30604 800
rect 30740 0 30796 800
rect 30836 0 30892 800
rect 30932 0 30988 800
rect 31028 0 31084 800
rect 31220 0 31276 800
rect 31316 0 31372 800
rect 31412 0 31468 800
rect 31604 0 31660 800
rect 31700 0 31756 800
rect 31796 0 31852 800
rect 31892 0 31948 800
rect 32084 0 32140 800
rect 32180 0 32236 800
rect 32276 0 32332 800
rect 32468 0 32524 800
rect 32564 0 32620 800
rect 32660 0 32716 800
rect 32756 0 32812 800
rect 32948 0 33004 800
rect 33044 0 33100 800
rect 33140 0 33196 800
rect 33236 0 33292 800
rect 33428 0 33484 800
rect 33524 0 33580 800
rect 33620 0 33676 800
rect 33812 0 33868 800
rect 33908 0 33964 800
rect 34004 0 34060 800
rect 34100 0 34156 800
rect 34292 0 34348 800
rect 34388 0 34444 800
rect 34484 0 34540 800
rect 34580 0 34636 800
rect 34772 0 34828 800
rect 34868 0 34924 800
rect 34964 0 35020 800
rect 35156 0 35212 800
rect 35252 0 35308 800
rect 35348 0 35404 800
rect 35444 0 35500 800
rect 35636 0 35692 800
rect 35732 0 35788 800
rect 35828 0 35884 800
rect 36020 0 36076 800
rect 36116 0 36172 800
rect 36212 0 36268 800
rect 36308 0 36364 800
rect 36500 0 36556 800
rect 36596 0 36652 800
rect 36692 0 36748 800
rect 36788 0 36844 800
rect 36980 0 37036 800
rect 37076 0 37132 800
rect 37172 0 37228 800
rect 37364 0 37420 800
rect 37460 0 37516 800
rect 37556 0 37612 800
rect 37652 0 37708 800
rect 37844 0 37900 800
rect 37940 0 37996 800
rect 38036 0 38092 800
rect 38132 0 38188 800
rect 38324 0 38380 800
rect 38420 0 38476 800
rect 38516 0 38572 800
rect 38708 0 38764 800
rect 38804 0 38860 800
rect 38900 0 38956 800
rect 38996 0 39052 800
rect 39188 0 39244 800
rect 39284 0 39340 800
rect 39380 0 39436 800
rect 39476 0 39532 800
rect 39668 0 39724 800
rect 39764 0 39820 800
rect 39860 0 39916 800
rect 40052 0 40108 800
rect 40148 0 40204 800
rect 40244 0 40300 800
rect 40340 0 40396 800
rect 40532 0 40588 800
rect 40628 0 40684 800
rect 40724 0 40780 800
rect 40916 0 40972 800
rect 41012 0 41068 800
rect 41108 0 41164 800
rect 41204 0 41260 800
rect 41396 0 41452 800
rect 41492 0 41548 800
rect 41588 0 41644 800
rect 41684 0 41740 800
rect 41876 0 41932 800
rect 41972 0 42028 800
rect 42068 0 42124 800
rect 42260 0 42316 800
rect 42356 0 42412 800
rect 42452 0 42508 800
rect 42548 0 42604 800
rect 42740 0 42796 800
rect 42836 0 42892 800
rect 42932 0 42988 800
rect 43028 0 43084 800
rect 43220 0 43276 800
rect 43316 0 43372 800
rect 43412 0 43468 800
rect 43604 0 43660 800
rect 43700 0 43756 800
rect 43796 0 43852 800
rect 43892 0 43948 800
rect 44084 0 44140 800
rect 44180 0 44236 800
rect 44276 0 44332 800
rect 44468 0 44524 800
rect 44564 0 44620 800
rect 44660 0 44716 800
rect 44756 0 44812 800
rect 44948 0 45004 800
rect 45044 0 45100 800
rect 45140 0 45196 800
rect 45236 0 45292 800
rect 45428 0 45484 800
rect 45524 0 45580 800
rect 45620 0 45676 800
rect 45812 0 45868 800
rect 45908 0 45964 800
rect 46004 0 46060 800
rect 46100 0 46156 800
rect 46292 0 46348 800
rect 46388 0 46444 800
rect 46484 0 46540 800
rect 46580 0 46636 800
rect 46772 0 46828 800
rect 46868 0 46924 800
rect 46964 0 47020 800
rect 47156 0 47212 800
rect 47252 0 47308 800
rect 47348 0 47404 800
rect 47444 0 47500 800
rect 47636 0 47692 800
rect 47732 0 47788 800
rect 47828 0 47884 800
rect 48020 0 48076 800
rect 48116 0 48172 800
rect 48212 0 48268 800
rect 48308 0 48364 800
rect 48500 0 48556 800
rect 48596 0 48652 800
rect 48692 0 48748 800
rect 48788 0 48844 800
rect 48980 0 49036 800
rect 49076 0 49132 800
rect 49172 0 49228 800
rect 49364 0 49420 800
rect 49460 0 49516 800
rect 49556 0 49612 800
rect 49652 0 49708 800
rect 49844 0 49900 800
rect 49940 0 49996 800
rect 50036 0 50092 800
rect 50132 0 50188 800
rect 50324 0 50380 800
rect 50420 0 50476 800
rect 50516 0 50572 800
rect 50708 0 50764 800
rect 50804 0 50860 800
rect 50900 0 50956 800
rect 50996 0 51052 800
rect 51188 0 51244 800
rect 51284 0 51340 800
rect 51380 0 51436 800
rect 51476 0 51532 800
rect 51668 0 51724 800
rect 51764 0 51820 800
rect 51860 0 51916 800
rect 52052 0 52108 800
rect 52148 0 52204 800
rect 52244 0 52300 800
rect 52340 0 52396 800
rect 52532 0 52588 800
rect 52628 0 52684 800
rect 52724 0 52780 800
rect 52916 0 52972 800
rect 53012 0 53068 800
rect 53108 0 53164 800
rect 53204 0 53260 800
rect 53396 0 53452 800
rect 53492 0 53548 800
rect 53588 0 53644 800
rect 53684 0 53740 800
rect 53876 0 53932 800
rect 53972 0 54028 800
rect 54068 0 54124 800
rect 54260 0 54316 800
rect 54356 0 54412 800
rect 54452 0 54508 800
rect 54548 0 54604 800
rect 54740 0 54796 800
rect 54836 0 54892 800
rect 54932 0 54988 800
rect 55028 0 55084 800
rect 55220 0 55276 800
rect 55316 0 55372 800
rect 55412 0 55468 800
rect 55604 0 55660 800
rect 55700 0 55756 800
rect 55796 0 55852 800
rect 55892 0 55948 800
rect 56084 0 56140 800
rect 56180 0 56236 800
rect 56276 0 56332 800
rect 56468 0 56524 800
rect 56564 0 56620 800
rect 56660 0 56716 800
rect 56756 0 56812 800
rect 56948 0 57004 800
rect 57044 0 57100 800
rect 57140 0 57196 800
rect 57236 0 57292 800
rect 57428 0 57484 800
rect 57524 0 57580 800
rect 57620 0 57676 800
rect 57812 0 57868 800
rect 57908 0 57964 800
rect 58004 0 58060 800
rect 58100 0 58156 800
rect 58292 0 58348 800
rect 58388 0 58444 800
rect 58484 0 58540 800
rect 58580 0 58636 800
rect 58772 0 58828 800
rect 58868 0 58924 800
rect 58964 0 59020 800
rect 59156 0 59212 800
rect 59252 0 59308 800
rect 59348 0 59404 800
rect 59444 0 59500 800
rect 59636 0 59692 800
rect 59732 0 59788 800
rect 59828 0 59884 800
<< via2 >>
rect 4268 57302 4324 57304
rect 4348 57302 4404 57304
rect 4428 57302 4484 57304
rect 4508 57302 4564 57304
rect 4268 57250 4294 57302
rect 4294 57250 4324 57302
rect 4348 57250 4358 57302
rect 4358 57250 4404 57302
rect 4428 57250 4474 57302
rect 4474 57250 4484 57302
rect 4508 57250 4538 57302
rect 4538 57250 4564 57302
rect 4268 57248 4324 57250
rect 4348 57248 4404 57250
rect 4428 57248 4484 57250
rect 4508 57248 4564 57250
rect 4268 55970 4324 55972
rect 4348 55970 4404 55972
rect 4428 55970 4484 55972
rect 4508 55970 4564 55972
rect 4268 55918 4294 55970
rect 4294 55918 4324 55970
rect 4348 55918 4358 55970
rect 4358 55918 4404 55970
rect 4428 55918 4474 55970
rect 4474 55918 4484 55970
rect 4508 55918 4538 55970
rect 4538 55918 4564 55970
rect 4268 55916 4324 55918
rect 4348 55916 4404 55918
rect 4428 55916 4484 55918
rect 4508 55916 4564 55918
rect 4268 54638 4324 54640
rect 4348 54638 4404 54640
rect 4428 54638 4484 54640
rect 4508 54638 4564 54640
rect 4268 54586 4294 54638
rect 4294 54586 4324 54638
rect 4348 54586 4358 54638
rect 4358 54586 4404 54638
rect 4428 54586 4474 54638
rect 4474 54586 4484 54638
rect 4508 54586 4538 54638
rect 4538 54586 4564 54638
rect 4268 54584 4324 54586
rect 4348 54584 4404 54586
rect 4428 54584 4484 54586
rect 4508 54584 4564 54586
rect 4268 53306 4324 53308
rect 4348 53306 4404 53308
rect 4428 53306 4484 53308
rect 4508 53306 4564 53308
rect 4268 53254 4294 53306
rect 4294 53254 4324 53306
rect 4348 53254 4358 53306
rect 4358 53254 4404 53306
rect 4428 53254 4474 53306
rect 4474 53254 4484 53306
rect 4508 53254 4538 53306
rect 4538 53254 4564 53306
rect 4268 53252 4324 53254
rect 4348 53252 4404 53254
rect 4428 53252 4484 53254
rect 4508 53252 4564 53254
rect 4268 51974 4324 51976
rect 4348 51974 4404 51976
rect 4428 51974 4484 51976
rect 4508 51974 4564 51976
rect 4268 51922 4294 51974
rect 4294 51922 4324 51974
rect 4348 51922 4358 51974
rect 4358 51922 4404 51974
rect 4428 51922 4474 51974
rect 4474 51922 4484 51974
rect 4508 51922 4538 51974
rect 4538 51922 4564 51974
rect 4268 51920 4324 51922
rect 4348 51920 4404 51922
rect 4428 51920 4484 51922
rect 4508 51920 4564 51922
rect 4268 50642 4324 50644
rect 4348 50642 4404 50644
rect 4428 50642 4484 50644
rect 4508 50642 4564 50644
rect 4268 50590 4294 50642
rect 4294 50590 4324 50642
rect 4348 50590 4358 50642
rect 4358 50590 4404 50642
rect 4428 50590 4474 50642
rect 4474 50590 4484 50642
rect 4508 50590 4538 50642
rect 4538 50590 4564 50642
rect 4268 50588 4324 50590
rect 4348 50588 4404 50590
rect 4428 50588 4484 50590
rect 4508 50588 4564 50590
rect 4268 49310 4324 49312
rect 4348 49310 4404 49312
rect 4428 49310 4484 49312
rect 4508 49310 4564 49312
rect 4268 49258 4294 49310
rect 4294 49258 4324 49310
rect 4348 49258 4358 49310
rect 4358 49258 4404 49310
rect 4428 49258 4474 49310
rect 4474 49258 4484 49310
rect 4508 49258 4538 49310
rect 4538 49258 4564 49310
rect 4268 49256 4324 49258
rect 4348 49256 4404 49258
rect 4428 49256 4484 49258
rect 4508 49256 4564 49258
rect 4268 47978 4324 47980
rect 4348 47978 4404 47980
rect 4428 47978 4484 47980
rect 4508 47978 4564 47980
rect 4268 47926 4294 47978
rect 4294 47926 4324 47978
rect 4348 47926 4358 47978
rect 4358 47926 4404 47978
rect 4428 47926 4474 47978
rect 4474 47926 4484 47978
rect 4508 47926 4538 47978
rect 4538 47926 4564 47978
rect 4268 47924 4324 47926
rect 4348 47924 4404 47926
rect 4428 47924 4484 47926
rect 4508 47924 4564 47926
rect 4268 46646 4324 46648
rect 4348 46646 4404 46648
rect 4428 46646 4484 46648
rect 4508 46646 4564 46648
rect 4268 46594 4294 46646
rect 4294 46594 4324 46646
rect 4348 46594 4358 46646
rect 4358 46594 4404 46646
rect 4428 46594 4474 46646
rect 4474 46594 4484 46646
rect 4508 46594 4538 46646
rect 4538 46594 4564 46646
rect 4268 46592 4324 46594
rect 4348 46592 4404 46594
rect 4428 46592 4484 46594
rect 4508 46592 4564 46594
rect 4268 45314 4324 45316
rect 4348 45314 4404 45316
rect 4428 45314 4484 45316
rect 4508 45314 4564 45316
rect 4268 45262 4294 45314
rect 4294 45262 4324 45314
rect 4348 45262 4358 45314
rect 4358 45262 4404 45314
rect 4428 45262 4474 45314
rect 4474 45262 4484 45314
rect 4508 45262 4538 45314
rect 4538 45262 4564 45314
rect 4268 45260 4324 45262
rect 4348 45260 4404 45262
rect 4428 45260 4484 45262
rect 4508 45260 4564 45262
rect 4268 43982 4324 43984
rect 4348 43982 4404 43984
rect 4428 43982 4484 43984
rect 4508 43982 4564 43984
rect 4268 43930 4294 43982
rect 4294 43930 4324 43982
rect 4348 43930 4358 43982
rect 4358 43930 4404 43982
rect 4428 43930 4474 43982
rect 4474 43930 4484 43982
rect 4508 43930 4538 43982
rect 4538 43930 4564 43982
rect 4268 43928 4324 43930
rect 4348 43928 4404 43930
rect 4428 43928 4484 43930
rect 4508 43928 4564 43930
rect 4268 42650 4324 42652
rect 4348 42650 4404 42652
rect 4428 42650 4484 42652
rect 4508 42650 4564 42652
rect 4268 42598 4294 42650
rect 4294 42598 4324 42650
rect 4348 42598 4358 42650
rect 4358 42598 4404 42650
rect 4428 42598 4474 42650
rect 4474 42598 4484 42650
rect 4508 42598 4538 42650
rect 4538 42598 4564 42650
rect 4268 42596 4324 42598
rect 4348 42596 4404 42598
rect 4428 42596 4484 42598
rect 4508 42596 4564 42598
rect 4268 41318 4324 41320
rect 4348 41318 4404 41320
rect 4428 41318 4484 41320
rect 4508 41318 4564 41320
rect 4268 41266 4294 41318
rect 4294 41266 4324 41318
rect 4348 41266 4358 41318
rect 4358 41266 4404 41318
rect 4428 41266 4474 41318
rect 4474 41266 4484 41318
rect 4508 41266 4538 41318
rect 4538 41266 4564 41318
rect 4268 41264 4324 41266
rect 4348 41264 4404 41266
rect 4428 41264 4484 41266
rect 4508 41264 4564 41266
rect 4268 39986 4324 39988
rect 4348 39986 4404 39988
rect 4428 39986 4484 39988
rect 4508 39986 4564 39988
rect 4268 39934 4294 39986
rect 4294 39934 4324 39986
rect 4348 39934 4358 39986
rect 4358 39934 4404 39986
rect 4428 39934 4474 39986
rect 4474 39934 4484 39986
rect 4508 39934 4538 39986
rect 4538 39934 4564 39986
rect 4268 39932 4324 39934
rect 4348 39932 4404 39934
rect 4428 39932 4484 39934
rect 4508 39932 4564 39934
rect 4268 38654 4324 38656
rect 4348 38654 4404 38656
rect 4428 38654 4484 38656
rect 4508 38654 4564 38656
rect 4268 38602 4294 38654
rect 4294 38602 4324 38654
rect 4348 38602 4358 38654
rect 4358 38602 4404 38654
rect 4428 38602 4474 38654
rect 4474 38602 4484 38654
rect 4508 38602 4538 38654
rect 4538 38602 4564 38654
rect 4268 38600 4324 38602
rect 4348 38600 4404 38602
rect 4428 38600 4484 38602
rect 4508 38600 4564 38602
rect 4268 37322 4324 37324
rect 4348 37322 4404 37324
rect 4428 37322 4484 37324
rect 4508 37322 4564 37324
rect 4268 37270 4294 37322
rect 4294 37270 4324 37322
rect 4348 37270 4358 37322
rect 4358 37270 4404 37322
rect 4428 37270 4474 37322
rect 4474 37270 4484 37322
rect 4508 37270 4538 37322
rect 4538 37270 4564 37322
rect 4268 37268 4324 37270
rect 4348 37268 4404 37270
rect 4428 37268 4484 37270
rect 4508 37268 4564 37270
rect 4268 35990 4324 35992
rect 4348 35990 4404 35992
rect 4428 35990 4484 35992
rect 4508 35990 4564 35992
rect 4268 35938 4294 35990
rect 4294 35938 4324 35990
rect 4348 35938 4358 35990
rect 4358 35938 4404 35990
rect 4428 35938 4474 35990
rect 4474 35938 4484 35990
rect 4508 35938 4538 35990
rect 4538 35938 4564 35990
rect 4268 35936 4324 35938
rect 4348 35936 4404 35938
rect 4428 35936 4484 35938
rect 4508 35936 4564 35938
rect 4268 34658 4324 34660
rect 4348 34658 4404 34660
rect 4428 34658 4484 34660
rect 4508 34658 4564 34660
rect 4268 34606 4294 34658
rect 4294 34606 4324 34658
rect 4348 34606 4358 34658
rect 4358 34606 4404 34658
rect 4428 34606 4474 34658
rect 4474 34606 4484 34658
rect 4508 34606 4538 34658
rect 4538 34606 4564 34658
rect 4268 34604 4324 34606
rect 4348 34604 4404 34606
rect 4428 34604 4484 34606
rect 4508 34604 4564 34606
rect 4268 33326 4324 33328
rect 4348 33326 4404 33328
rect 4428 33326 4484 33328
rect 4508 33326 4564 33328
rect 4268 33274 4294 33326
rect 4294 33274 4324 33326
rect 4348 33274 4358 33326
rect 4358 33274 4404 33326
rect 4428 33274 4474 33326
rect 4474 33274 4484 33326
rect 4508 33274 4538 33326
rect 4538 33274 4564 33326
rect 4268 33272 4324 33274
rect 4348 33272 4404 33274
rect 4428 33272 4484 33274
rect 4508 33272 4564 33274
rect 4268 31994 4324 31996
rect 4348 31994 4404 31996
rect 4428 31994 4484 31996
rect 4508 31994 4564 31996
rect 4268 31942 4294 31994
rect 4294 31942 4324 31994
rect 4348 31942 4358 31994
rect 4358 31942 4404 31994
rect 4428 31942 4474 31994
rect 4474 31942 4484 31994
rect 4508 31942 4538 31994
rect 4538 31942 4564 31994
rect 4268 31940 4324 31942
rect 4348 31940 4404 31942
rect 4428 31940 4484 31942
rect 4508 31940 4564 31942
rect 4268 30662 4324 30664
rect 4348 30662 4404 30664
rect 4428 30662 4484 30664
rect 4508 30662 4564 30664
rect 4268 30610 4294 30662
rect 4294 30610 4324 30662
rect 4348 30610 4358 30662
rect 4358 30610 4404 30662
rect 4428 30610 4474 30662
rect 4474 30610 4484 30662
rect 4508 30610 4538 30662
rect 4538 30610 4564 30662
rect 4268 30608 4324 30610
rect 4348 30608 4404 30610
rect 4428 30608 4484 30610
rect 4508 30608 4564 30610
rect 4268 29330 4324 29332
rect 4348 29330 4404 29332
rect 4428 29330 4484 29332
rect 4508 29330 4564 29332
rect 4268 29278 4294 29330
rect 4294 29278 4324 29330
rect 4348 29278 4358 29330
rect 4358 29278 4404 29330
rect 4428 29278 4474 29330
rect 4474 29278 4484 29330
rect 4508 29278 4538 29330
rect 4538 29278 4564 29330
rect 4268 29276 4324 29278
rect 4348 29276 4404 29278
rect 4428 29276 4484 29278
rect 4508 29276 4564 29278
rect 4268 27998 4324 28000
rect 4348 27998 4404 28000
rect 4428 27998 4484 28000
rect 4508 27998 4564 28000
rect 4268 27946 4294 27998
rect 4294 27946 4324 27998
rect 4348 27946 4358 27998
rect 4358 27946 4404 27998
rect 4428 27946 4474 27998
rect 4474 27946 4484 27998
rect 4508 27946 4538 27998
rect 4538 27946 4564 27998
rect 4268 27944 4324 27946
rect 4348 27944 4404 27946
rect 4428 27944 4484 27946
rect 4508 27944 4564 27946
rect 4268 26666 4324 26668
rect 4348 26666 4404 26668
rect 4428 26666 4484 26668
rect 4508 26666 4564 26668
rect 4268 26614 4294 26666
rect 4294 26614 4324 26666
rect 4348 26614 4358 26666
rect 4358 26614 4404 26666
rect 4428 26614 4474 26666
rect 4474 26614 4484 26666
rect 4508 26614 4538 26666
rect 4538 26614 4564 26666
rect 4268 26612 4324 26614
rect 4348 26612 4404 26614
rect 4428 26612 4484 26614
rect 4508 26612 4564 26614
rect 4268 25334 4324 25336
rect 4348 25334 4404 25336
rect 4428 25334 4484 25336
rect 4508 25334 4564 25336
rect 4268 25282 4294 25334
rect 4294 25282 4324 25334
rect 4348 25282 4358 25334
rect 4358 25282 4404 25334
rect 4428 25282 4474 25334
rect 4474 25282 4484 25334
rect 4508 25282 4538 25334
rect 4538 25282 4564 25334
rect 4268 25280 4324 25282
rect 4348 25280 4404 25282
rect 4428 25280 4484 25282
rect 4508 25280 4564 25282
rect 4268 24002 4324 24004
rect 4348 24002 4404 24004
rect 4428 24002 4484 24004
rect 4508 24002 4564 24004
rect 4268 23950 4294 24002
rect 4294 23950 4324 24002
rect 4348 23950 4358 24002
rect 4358 23950 4404 24002
rect 4428 23950 4474 24002
rect 4474 23950 4484 24002
rect 4508 23950 4538 24002
rect 4538 23950 4564 24002
rect 4268 23948 4324 23950
rect 4348 23948 4404 23950
rect 4428 23948 4484 23950
rect 4508 23948 4564 23950
rect 4268 22670 4324 22672
rect 4348 22670 4404 22672
rect 4428 22670 4484 22672
rect 4508 22670 4564 22672
rect 4268 22618 4294 22670
rect 4294 22618 4324 22670
rect 4348 22618 4358 22670
rect 4358 22618 4404 22670
rect 4428 22618 4474 22670
rect 4474 22618 4484 22670
rect 4508 22618 4538 22670
rect 4538 22618 4564 22670
rect 4268 22616 4324 22618
rect 4348 22616 4404 22618
rect 4428 22616 4484 22618
rect 4508 22616 4564 22618
rect 4268 21338 4324 21340
rect 4348 21338 4404 21340
rect 4428 21338 4484 21340
rect 4508 21338 4564 21340
rect 4268 21286 4294 21338
rect 4294 21286 4324 21338
rect 4348 21286 4358 21338
rect 4358 21286 4404 21338
rect 4428 21286 4474 21338
rect 4474 21286 4484 21338
rect 4508 21286 4538 21338
rect 4538 21286 4564 21338
rect 4268 21284 4324 21286
rect 4348 21284 4404 21286
rect 4428 21284 4484 21286
rect 4508 21284 4564 21286
rect 4268 20006 4324 20008
rect 4348 20006 4404 20008
rect 4428 20006 4484 20008
rect 4508 20006 4564 20008
rect 4268 19954 4294 20006
rect 4294 19954 4324 20006
rect 4348 19954 4358 20006
rect 4358 19954 4404 20006
rect 4428 19954 4474 20006
rect 4474 19954 4484 20006
rect 4508 19954 4538 20006
rect 4538 19954 4564 20006
rect 4268 19952 4324 19954
rect 4348 19952 4404 19954
rect 4428 19952 4484 19954
rect 4508 19952 4564 19954
rect 4268 18674 4324 18676
rect 4348 18674 4404 18676
rect 4428 18674 4484 18676
rect 4508 18674 4564 18676
rect 4268 18622 4294 18674
rect 4294 18622 4324 18674
rect 4348 18622 4358 18674
rect 4358 18622 4404 18674
rect 4428 18622 4474 18674
rect 4474 18622 4484 18674
rect 4508 18622 4538 18674
rect 4538 18622 4564 18674
rect 4268 18620 4324 18622
rect 4348 18620 4404 18622
rect 4428 18620 4484 18622
rect 4508 18620 4564 18622
rect 4268 17342 4324 17344
rect 4348 17342 4404 17344
rect 4428 17342 4484 17344
rect 4508 17342 4564 17344
rect 4268 17290 4294 17342
rect 4294 17290 4324 17342
rect 4348 17290 4358 17342
rect 4358 17290 4404 17342
rect 4428 17290 4474 17342
rect 4474 17290 4484 17342
rect 4508 17290 4538 17342
rect 4538 17290 4564 17342
rect 4268 17288 4324 17290
rect 4348 17288 4404 17290
rect 4428 17288 4484 17290
rect 4508 17288 4564 17290
rect 4268 16010 4324 16012
rect 4348 16010 4404 16012
rect 4428 16010 4484 16012
rect 4508 16010 4564 16012
rect 4268 15958 4294 16010
rect 4294 15958 4324 16010
rect 4348 15958 4358 16010
rect 4358 15958 4404 16010
rect 4428 15958 4474 16010
rect 4474 15958 4484 16010
rect 4508 15958 4538 16010
rect 4538 15958 4564 16010
rect 4268 15956 4324 15958
rect 4348 15956 4404 15958
rect 4428 15956 4484 15958
rect 4508 15956 4564 15958
rect 4268 14678 4324 14680
rect 4348 14678 4404 14680
rect 4428 14678 4484 14680
rect 4508 14678 4564 14680
rect 4268 14626 4294 14678
rect 4294 14626 4324 14678
rect 4348 14626 4358 14678
rect 4358 14626 4404 14678
rect 4428 14626 4474 14678
rect 4474 14626 4484 14678
rect 4508 14626 4538 14678
rect 4538 14626 4564 14678
rect 4268 14624 4324 14626
rect 4348 14624 4404 14626
rect 4428 14624 4484 14626
rect 4508 14624 4564 14626
rect 4268 13346 4324 13348
rect 4348 13346 4404 13348
rect 4428 13346 4484 13348
rect 4508 13346 4564 13348
rect 4268 13294 4294 13346
rect 4294 13294 4324 13346
rect 4348 13294 4358 13346
rect 4358 13294 4404 13346
rect 4428 13294 4474 13346
rect 4474 13294 4484 13346
rect 4508 13294 4538 13346
rect 4538 13294 4564 13346
rect 4268 13292 4324 13294
rect 4348 13292 4404 13294
rect 4428 13292 4484 13294
rect 4508 13292 4564 13294
rect 4268 12014 4324 12016
rect 4348 12014 4404 12016
rect 4428 12014 4484 12016
rect 4508 12014 4564 12016
rect 4268 11962 4294 12014
rect 4294 11962 4324 12014
rect 4348 11962 4358 12014
rect 4358 11962 4404 12014
rect 4428 11962 4474 12014
rect 4474 11962 4484 12014
rect 4508 11962 4538 12014
rect 4538 11962 4564 12014
rect 4268 11960 4324 11962
rect 4348 11960 4404 11962
rect 4428 11960 4484 11962
rect 4508 11960 4564 11962
rect 4268 10682 4324 10684
rect 4348 10682 4404 10684
rect 4428 10682 4484 10684
rect 4508 10682 4564 10684
rect 4268 10630 4294 10682
rect 4294 10630 4324 10682
rect 4348 10630 4358 10682
rect 4358 10630 4404 10682
rect 4428 10630 4474 10682
rect 4474 10630 4484 10682
rect 4508 10630 4538 10682
rect 4538 10630 4564 10682
rect 4268 10628 4324 10630
rect 4348 10628 4404 10630
rect 4428 10628 4484 10630
rect 4508 10628 4564 10630
rect 4268 9350 4324 9352
rect 4348 9350 4404 9352
rect 4428 9350 4484 9352
rect 4508 9350 4564 9352
rect 4268 9298 4294 9350
rect 4294 9298 4324 9350
rect 4348 9298 4358 9350
rect 4358 9298 4404 9350
rect 4428 9298 4474 9350
rect 4474 9298 4484 9350
rect 4508 9298 4538 9350
rect 4538 9298 4564 9350
rect 4268 9296 4324 9298
rect 4348 9296 4404 9298
rect 4428 9296 4484 9298
rect 4508 9296 4564 9298
rect 4268 8018 4324 8020
rect 4348 8018 4404 8020
rect 4428 8018 4484 8020
rect 4508 8018 4564 8020
rect 4268 7966 4294 8018
rect 4294 7966 4324 8018
rect 4348 7966 4358 8018
rect 4358 7966 4404 8018
rect 4428 7966 4474 8018
rect 4474 7966 4484 8018
rect 4508 7966 4538 8018
rect 4538 7966 4564 8018
rect 4268 7964 4324 7966
rect 4348 7964 4404 7966
rect 4428 7964 4484 7966
rect 4508 7964 4564 7966
rect 4268 6686 4324 6688
rect 4348 6686 4404 6688
rect 4428 6686 4484 6688
rect 4508 6686 4564 6688
rect 4268 6634 4294 6686
rect 4294 6634 4324 6686
rect 4348 6634 4358 6686
rect 4358 6634 4404 6686
rect 4428 6634 4474 6686
rect 4474 6634 4484 6686
rect 4508 6634 4538 6686
rect 4538 6634 4564 6686
rect 4268 6632 4324 6634
rect 4348 6632 4404 6634
rect 4428 6632 4484 6634
rect 4508 6632 4564 6634
rect 4268 5354 4324 5356
rect 4348 5354 4404 5356
rect 4428 5354 4484 5356
rect 4508 5354 4564 5356
rect 4268 5302 4294 5354
rect 4294 5302 4324 5354
rect 4348 5302 4358 5354
rect 4358 5302 4404 5354
rect 4428 5302 4474 5354
rect 4474 5302 4484 5354
rect 4508 5302 4538 5354
rect 4538 5302 4564 5354
rect 4268 5300 4324 5302
rect 4348 5300 4404 5302
rect 4428 5300 4484 5302
rect 4508 5300 4564 5302
rect 4268 4022 4324 4024
rect 4348 4022 4404 4024
rect 4428 4022 4484 4024
rect 4508 4022 4564 4024
rect 4268 3970 4294 4022
rect 4294 3970 4324 4022
rect 4348 3970 4358 4022
rect 4358 3970 4404 4022
rect 4428 3970 4474 4022
rect 4474 3970 4484 4022
rect 4508 3970 4538 4022
rect 4538 3970 4564 4022
rect 4268 3968 4324 3970
rect 4348 3968 4404 3970
rect 4428 3968 4484 3970
rect 4508 3968 4564 3970
rect 4268 2690 4324 2692
rect 4348 2690 4404 2692
rect 4428 2690 4484 2692
rect 4508 2690 4564 2692
rect 4268 2638 4294 2690
rect 4294 2638 4324 2690
rect 4348 2638 4358 2690
rect 4358 2638 4404 2690
rect 4428 2638 4474 2690
rect 4474 2638 4484 2690
rect 4508 2638 4538 2690
rect 4538 2638 4564 2690
rect 4268 2636 4324 2638
rect 4348 2636 4404 2638
rect 4428 2636 4484 2638
rect 4508 2636 4564 2638
rect 19628 56636 19684 56638
rect 19708 56636 19764 56638
rect 19788 56636 19844 56638
rect 19868 56636 19924 56638
rect 19628 56584 19654 56636
rect 19654 56584 19684 56636
rect 19708 56584 19718 56636
rect 19718 56584 19764 56636
rect 19788 56584 19834 56636
rect 19834 56584 19844 56636
rect 19868 56584 19898 56636
rect 19898 56584 19924 56636
rect 19628 56582 19684 56584
rect 19708 56582 19764 56584
rect 19788 56582 19844 56584
rect 19868 56582 19924 56584
rect 19628 55304 19684 55306
rect 19708 55304 19764 55306
rect 19788 55304 19844 55306
rect 19868 55304 19924 55306
rect 19628 55252 19654 55304
rect 19654 55252 19684 55304
rect 19708 55252 19718 55304
rect 19718 55252 19764 55304
rect 19788 55252 19834 55304
rect 19834 55252 19844 55304
rect 19868 55252 19898 55304
rect 19898 55252 19924 55304
rect 19628 55250 19684 55252
rect 19708 55250 19764 55252
rect 19788 55250 19844 55252
rect 19868 55250 19924 55252
rect 19628 53972 19684 53974
rect 19708 53972 19764 53974
rect 19788 53972 19844 53974
rect 19868 53972 19924 53974
rect 19628 53920 19654 53972
rect 19654 53920 19684 53972
rect 19708 53920 19718 53972
rect 19718 53920 19764 53972
rect 19788 53920 19834 53972
rect 19834 53920 19844 53972
rect 19868 53920 19898 53972
rect 19898 53920 19924 53972
rect 19628 53918 19684 53920
rect 19708 53918 19764 53920
rect 19788 53918 19844 53920
rect 19868 53918 19924 53920
rect 19628 52640 19684 52642
rect 19708 52640 19764 52642
rect 19788 52640 19844 52642
rect 19868 52640 19924 52642
rect 19628 52588 19654 52640
rect 19654 52588 19684 52640
rect 19708 52588 19718 52640
rect 19718 52588 19764 52640
rect 19788 52588 19834 52640
rect 19834 52588 19844 52640
rect 19868 52588 19898 52640
rect 19898 52588 19924 52640
rect 19628 52586 19684 52588
rect 19708 52586 19764 52588
rect 19788 52586 19844 52588
rect 19868 52586 19924 52588
rect 19628 51308 19684 51310
rect 19708 51308 19764 51310
rect 19788 51308 19844 51310
rect 19868 51308 19924 51310
rect 19628 51256 19654 51308
rect 19654 51256 19684 51308
rect 19708 51256 19718 51308
rect 19718 51256 19764 51308
rect 19788 51256 19834 51308
rect 19834 51256 19844 51308
rect 19868 51256 19898 51308
rect 19898 51256 19924 51308
rect 19628 51254 19684 51256
rect 19708 51254 19764 51256
rect 19788 51254 19844 51256
rect 19868 51254 19924 51256
rect 19628 49976 19684 49978
rect 19708 49976 19764 49978
rect 19788 49976 19844 49978
rect 19868 49976 19924 49978
rect 19628 49924 19654 49976
rect 19654 49924 19684 49976
rect 19708 49924 19718 49976
rect 19718 49924 19764 49976
rect 19788 49924 19834 49976
rect 19834 49924 19844 49976
rect 19868 49924 19898 49976
rect 19898 49924 19924 49976
rect 19628 49922 19684 49924
rect 19708 49922 19764 49924
rect 19788 49922 19844 49924
rect 19868 49922 19924 49924
rect 19628 48644 19684 48646
rect 19708 48644 19764 48646
rect 19788 48644 19844 48646
rect 19868 48644 19924 48646
rect 19628 48592 19654 48644
rect 19654 48592 19684 48644
rect 19708 48592 19718 48644
rect 19718 48592 19764 48644
rect 19788 48592 19834 48644
rect 19834 48592 19844 48644
rect 19868 48592 19898 48644
rect 19898 48592 19924 48644
rect 19628 48590 19684 48592
rect 19708 48590 19764 48592
rect 19788 48590 19844 48592
rect 19868 48590 19924 48592
rect 19628 47312 19684 47314
rect 19708 47312 19764 47314
rect 19788 47312 19844 47314
rect 19868 47312 19924 47314
rect 19628 47260 19654 47312
rect 19654 47260 19684 47312
rect 19708 47260 19718 47312
rect 19718 47260 19764 47312
rect 19788 47260 19834 47312
rect 19834 47260 19844 47312
rect 19868 47260 19898 47312
rect 19898 47260 19924 47312
rect 19628 47258 19684 47260
rect 19708 47258 19764 47260
rect 19788 47258 19844 47260
rect 19868 47258 19924 47260
rect 19628 45980 19684 45982
rect 19708 45980 19764 45982
rect 19788 45980 19844 45982
rect 19868 45980 19924 45982
rect 19628 45928 19654 45980
rect 19654 45928 19684 45980
rect 19708 45928 19718 45980
rect 19718 45928 19764 45980
rect 19788 45928 19834 45980
rect 19834 45928 19844 45980
rect 19868 45928 19898 45980
rect 19898 45928 19924 45980
rect 19628 45926 19684 45928
rect 19708 45926 19764 45928
rect 19788 45926 19844 45928
rect 19868 45926 19924 45928
rect 19628 44648 19684 44650
rect 19708 44648 19764 44650
rect 19788 44648 19844 44650
rect 19868 44648 19924 44650
rect 19628 44596 19654 44648
rect 19654 44596 19684 44648
rect 19708 44596 19718 44648
rect 19718 44596 19764 44648
rect 19788 44596 19834 44648
rect 19834 44596 19844 44648
rect 19868 44596 19898 44648
rect 19898 44596 19924 44648
rect 19628 44594 19684 44596
rect 19708 44594 19764 44596
rect 19788 44594 19844 44596
rect 19868 44594 19924 44596
rect 19628 43316 19684 43318
rect 19708 43316 19764 43318
rect 19788 43316 19844 43318
rect 19868 43316 19924 43318
rect 19628 43264 19654 43316
rect 19654 43264 19684 43316
rect 19708 43264 19718 43316
rect 19718 43264 19764 43316
rect 19788 43264 19834 43316
rect 19834 43264 19844 43316
rect 19868 43264 19898 43316
rect 19898 43264 19924 43316
rect 19628 43262 19684 43264
rect 19708 43262 19764 43264
rect 19788 43262 19844 43264
rect 19868 43262 19924 43264
rect 19628 41984 19684 41986
rect 19708 41984 19764 41986
rect 19788 41984 19844 41986
rect 19868 41984 19924 41986
rect 19628 41932 19654 41984
rect 19654 41932 19684 41984
rect 19708 41932 19718 41984
rect 19718 41932 19764 41984
rect 19788 41932 19834 41984
rect 19834 41932 19844 41984
rect 19868 41932 19898 41984
rect 19898 41932 19924 41984
rect 19628 41930 19684 41932
rect 19708 41930 19764 41932
rect 19788 41930 19844 41932
rect 19868 41930 19924 41932
rect 19628 40652 19684 40654
rect 19708 40652 19764 40654
rect 19788 40652 19844 40654
rect 19868 40652 19924 40654
rect 19628 40600 19654 40652
rect 19654 40600 19684 40652
rect 19708 40600 19718 40652
rect 19718 40600 19764 40652
rect 19788 40600 19834 40652
rect 19834 40600 19844 40652
rect 19868 40600 19898 40652
rect 19898 40600 19924 40652
rect 19628 40598 19684 40600
rect 19708 40598 19764 40600
rect 19788 40598 19844 40600
rect 19868 40598 19924 40600
rect 19628 39320 19684 39322
rect 19708 39320 19764 39322
rect 19788 39320 19844 39322
rect 19868 39320 19924 39322
rect 19628 39268 19654 39320
rect 19654 39268 19684 39320
rect 19708 39268 19718 39320
rect 19718 39268 19764 39320
rect 19788 39268 19834 39320
rect 19834 39268 19844 39320
rect 19868 39268 19898 39320
rect 19898 39268 19924 39320
rect 19628 39266 19684 39268
rect 19708 39266 19764 39268
rect 19788 39266 19844 39268
rect 19868 39266 19924 39268
rect 19628 37988 19684 37990
rect 19708 37988 19764 37990
rect 19788 37988 19844 37990
rect 19868 37988 19924 37990
rect 19628 37936 19654 37988
rect 19654 37936 19684 37988
rect 19708 37936 19718 37988
rect 19718 37936 19764 37988
rect 19788 37936 19834 37988
rect 19834 37936 19844 37988
rect 19868 37936 19898 37988
rect 19898 37936 19924 37988
rect 19628 37934 19684 37936
rect 19708 37934 19764 37936
rect 19788 37934 19844 37936
rect 19868 37934 19924 37936
rect 19628 36656 19684 36658
rect 19708 36656 19764 36658
rect 19788 36656 19844 36658
rect 19868 36656 19924 36658
rect 19628 36604 19654 36656
rect 19654 36604 19684 36656
rect 19708 36604 19718 36656
rect 19718 36604 19764 36656
rect 19788 36604 19834 36656
rect 19834 36604 19844 36656
rect 19868 36604 19898 36656
rect 19898 36604 19924 36656
rect 19628 36602 19684 36604
rect 19708 36602 19764 36604
rect 19788 36602 19844 36604
rect 19868 36602 19924 36604
rect 19628 35324 19684 35326
rect 19708 35324 19764 35326
rect 19788 35324 19844 35326
rect 19868 35324 19924 35326
rect 19628 35272 19654 35324
rect 19654 35272 19684 35324
rect 19708 35272 19718 35324
rect 19718 35272 19764 35324
rect 19788 35272 19834 35324
rect 19834 35272 19844 35324
rect 19868 35272 19898 35324
rect 19898 35272 19924 35324
rect 19628 35270 19684 35272
rect 19708 35270 19764 35272
rect 19788 35270 19844 35272
rect 19868 35270 19924 35272
rect 19628 33992 19684 33994
rect 19708 33992 19764 33994
rect 19788 33992 19844 33994
rect 19868 33992 19924 33994
rect 19628 33940 19654 33992
rect 19654 33940 19684 33992
rect 19708 33940 19718 33992
rect 19718 33940 19764 33992
rect 19788 33940 19834 33992
rect 19834 33940 19844 33992
rect 19868 33940 19898 33992
rect 19898 33940 19924 33992
rect 19628 33938 19684 33940
rect 19708 33938 19764 33940
rect 19788 33938 19844 33940
rect 19868 33938 19924 33940
rect 19628 32660 19684 32662
rect 19708 32660 19764 32662
rect 19788 32660 19844 32662
rect 19868 32660 19924 32662
rect 19628 32608 19654 32660
rect 19654 32608 19684 32660
rect 19708 32608 19718 32660
rect 19718 32608 19764 32660
rect 19788 32608 19834 32660
rect 19834 32608 19844 32660
rect 19868 32608 19898 32660
rect 19898 32608 19924 32660
rect 19628 32606 19684 32608
rect 19708 32606 19764 32608
rect 19788 32606 19844 32608
rect 19868 32606 19924 32608
rect 19628 31328 19684 31330
rect 19708 31328 19764 31330
rect 19788 31328 19844 31330
rect 19868 31328 19924 31330
rect 19628 31276 19654 31328
rect 19654 31276 19684 31328
rect 19708 31276 19718 31328
rect 19718 31276 19764 31328
rect 19788 31276 19834 31328
rect 19834 31276 19844 31328
rect 19868 31276 19898 31328
rect 19898 31276 19924 31328
rect 19628 31274 19684 31276
rect 19708 31274 19764 31276
rect 19788 31274 19844 31276
rect 19868 31274 19924 31276
rect 19628 29996 19684 29998
rect 19708 29996 19764 29998
rect 19788 29996 19844 29998
rect 19868 29996 19924 29998
rect 19628 29944 19654 29996
rect 19654 29944 19684 29996
rect 19708 29944 19718 29996
rect 19718 29944 19764 29996
rect 19788 29944 19834 29996
rect 19834 29944 19844 29996
rect 19868 29944 19898 29996
rect 19898 29944 19924 29996
rect 19628 29942 19684 29944
rect 19708 29942 19764 29944
rect 19788 29942 19844 29944
rect 19868 29942 19924 29944
rect 19628 28664 19684 28666
rect 19708 28664 19764 28666
rect 19788 28664 19844 28666
rect 19868 28664 19924 28666
rect 19628 28612 19654 28664
rect 19654 28612 19684 28664
rect 19708 28612 19718 28664
rect 19718 28612 19764 28664
rect 19788 28612 19834 28664
rect 19834 28612 19844 28664
rect 19868 28612 19898 28664
rect 19898 28612 19924 28664
rect 19628 28610 19684 28612
rect 19708 28610 19764 28612
rect 19788 28610 19844 28612
rect 19868 28610 19924 28612
rect 19628 27332 19684 27334
rect 19708 27332 19764 27334
rect 19788 27332 19844 27334
rect 19868 27332 19924 27334
rect 19628 27280 19654 27332
rect 19654 27280 19684 27332
rect 19708 27280 19718 27332
rect 19718 27280 19764 27332
rect 19788 27280 19834 27332
rect 19834 27280 19844 27332
rect 19868 27280 19898 27332
rect 19898 27280 19924 27332
rect 19628 27278 19684 27280
rect 19708 27278 19764 27280
rect 19788 27278 19844 27280
rect 19868 27278 19924 27280
rect 19628 26000 19684 26002
rect 19708 26000 19764 26002
rect 19788 26000 19844 26002
rect 19868 26000 19924 26002
rect 19628 25948 19654 26000
rect 19654 25948 19684 26000
rect 19708 25948 19718 26000
rect 19718 25948 19764 26000
rect 19788 25948 19834 26000
rect 19834 25948 19844 26000
rect 19868 25948 19898 26000
rect 19898 25948 19924 26000
rect 19628 25946 19684 25948
rect 19708 25946 19764 25948
rect 19788 25946 19844 25948
rect 19868 25946 19924 25948
rect 19628 24668 19684 24670
rect 19708 24668 19764 24670
rect 19788 24668 19844 24670
rect 19868 24668 19924 24670
rect 19628 24616 19654 24668
rect 19654 24616 19684 24668
rect 19708 24616 19718 24668
rect 19718 24616 19764 24668
rect 19788 24616 19834 24668
rect 19834 24616 19844 24668
rect 19868 24616 19898 24668
rect 19898 24616 19924 24668
rect 19628 24614 19684 24616
rect 19708 24614 19764 24616
rect 19788 24614 19844 24616
rect 19868 24614 19924 24616
rect 19628 23336 19684 23338
rect 19708 23336 19764 23338
rect 19788 23336 19844 23338
rect 19868 23336 19924 23338
rect 19628 23284 19654 23336
rect 19654 23284 19684 23336
rect 19708 23284 19718 23336
rect 19718 23284 19764 23336
rect 19788 23284 19834 23336
rect 19834 23284 19844 23336
rect 19868 23284 19898 23336
rect 19898 23284 19924 23336
rect 19628 23282 19684 23284
rect 19708 23282 19764 23284
rect 19788 23282 19844 23284
rect 19868 23282 19924 23284
rect 19628 22004 19684 22006
rect 19708 22004 19764 22006
rect 19788 22004 19844 22006
rect 19868 22004 19924 22006
rect 19628 21952 19654 22004
rect 19654 21952 19684 22004
rect 19708 21952 19718 22004
rect 19718 21952 19764 22004
rect 19788 21952 19834 22004
rect 19834 21952 19844 22004
rect 19868 21952 19898 22004
rect 19898 21952 19924 22004
rect 19628 21950 19684 21952
rect 19708 21950 19764 21952
rect 19788 21950 19844 21952
rect 19868 21950 19924 21952
rect 19628 20672 19684 20674
rect 19708 20672 19764 20674
rect 19788 20672 19844 20674
rect 19868 20672 19924 20674
rect 19628 20620 19654 20672
rect 19654 20620 19684 20672
rect 19708 20620 19718 20672
rect 19718 20620 19764 20672
rect 19788 20620 19834 20672
rect 19834 20620 19844 20672
rect 19868 20620 19898 20672
rect 19898 20620 19924 20672
rect 19628 20618 19684 20620
rect 19708 20618 19764 20620
rect 19788 20618 19844 20620
rect 19868 20618 19924 20620
rect 19628 19340 19684 19342
rect 19708 19340 19764 19342
rect 19788 19340 19844 19342
rect 19868 19340 19924 19342
rect 19628 19288 19654 19340
rect 19654 19288 19684 19340
rect 19708 19288 19718 19340
rect 19718 19288 19764 19340
rect 19788 19288 19834 19340
rect 19834 19288 19844 19340
rect 19868 19288 19898 19340
rect 19898 19288 19924 19340
rect 19628 19286 19684 19288
rect 19708 19286 19764 19288
rect 19788 19286 19844 19288
rect 19868 19286 19924 19288
rect 19628 18008 19684 18010
rect 19708 18008 19764 18010
rect 19788 18008 19844 18010
rect 19868 18008 19924 18010
rect 19628 17956 19654 18008
rect 19654 17956 19684 18008
rect 19708 17956 19718 18008
rect 19718 17956 19764 18008
rect 19788 17956 19834 18008
rect 19834 17956 19844 18008
rect 19868 17956 19898 18008
rect 19898 17956 19924 18008
rect 19628 17954 19684 17956
rect 19708 17954 19764 17956
rect 19788 17954 19844 17956
rect 19868 17954 19924 17956
rect 19628 16676 19684 16678
rect 19708 16676 19764 16678
rect 19788 16676 19844 16678
rect 19868 16676 19924 16678
rect 19628 16624 19654 16676
rect 19654 16624 19684 16676
rect 19708 16624 19718 16676
rect 19718 16624 19764 16676
rect 19788 16624 19834 16676
rect 19834 16624 19844 16676
rect 19868 16624 19898 16676
rect 19898 16624 19924 16676
rect 19628 16622 19684 16624
rect 19708 16622 19764 16624
rect 19788 16622 19844 16624
rect 19868 16622 19924 16624
rect 19628 15344 19684 15346
rect 19708 15344 19764 15346
rect 19788 15344 19844 15346
rect 19868 15344 19924 15346
rect 19628 15292 19654 15344
rect 19654 15292 19684 15344
rect 19708 15292 19718 15344
rect 19718 15292 19764 15344
rect 19788 15292 19834 15344
rect 19834 15292 19844 15344
rect 19868 15292 19898 15344
rect 19898 15292 19924 15344
rect 19628 15290 19684 15292
rect 19708 15290 19764 15292
rect 19788 15290 19844 15292
rect 19868 15290 19924 15292
rect 19628 14012 19684 14014
rect 19708 14012 19764 14014
rect 19788 14012 19844 14014
rect 19868 14012 19924 14014
rect 19628 13960 19654 14012
rect 19654 13960 19684 14012
rect 19708 13960 19718 14012
rect 19718 13960 19764 14012
rect 19788 13960 19834 14012
rect 19834 13960 19844 14012
rect 19868 13960 19898 14012
rect 19898 13960 19924 14012
rect 19628 13958 19684 13960
rect 19708 13958 19764 13960
rect 19788 13958 19844 13960
rect 19868 13958 19924 13960
rect 19628 12680 19684 12682
rect 19708 12680 19764 12682
rect 19788 12680 19844 12682
rect 19868 12680 19924 12682
rect 19628 12628 19654 12680
rect 19654 12628 19684 12680
rect 19708 12628 19718 12680
rect 19718 12628 19764 12680
rect 19788 12628 19834 12680
rect 19834 12628 19844 12680
rect 19868 12628 19898 12680
rect 19898 12628 19924 12680
rect 19628 12626 19684 12628
rect 19708 12626 19764 12628
rect 19788 12626 19844 12628
rect 19868 12626 19924 12628
rect 19628 11348 19684 11350
rect 19708 11348 19764 11350
rect 19788 11348 19844 11350
rect 19868 11348 19924 11350
rect 19628 11296 19654 11348
rect 19654 11296 19684 11348
rect 19708 11296 19718 11348
rect 19718 11296 19764 11348
rect 19788 11296 19834 11348
rect 19834 11296 19844 11348
rect 19868 11296 19898 11348
rect 19898 11296 19924 11348
rect 19628 11294 19684 11296
rect 19708 11294 19764 11296
rect 19788 11294 19844 11296
rect 19868 11294 19924 11296
rect 19628 10016 19684 10018
rect 19708 10016 19764 10018
rect 19788 10016 19844 10018
rect 19868 10016 19924 10018
rect 19628 9964 19654 10016
rect 19654 9964 19684 10016
rect 19708 9964 19718 10016
rect 19718 9964 19764 10016
rect 19788 9964 19834 10016
rect 19834 9964 19844 10016
rect 19868 9964 19898 10016
rect 19898 9964 19924 10016
rect 19628 9962 19684 9964
rect 19708 9962 19764 9964
rect 19788 9962 19844 9964
rect 19868 9962 19924 9964
rect 19628 8684 19684 8686
rect 19708 8684 19764 8686
rect 19788 8684 19844 8686
rect 19868 8684 19924 8686
rect 19628 8632 19654 8684
rect 19654 8632 19684 8684
rect 19708 8632 19718 8684
rect 19718 8632 19764 8684
rect 19788 8632 19834 8684
rect 19834 8632 19844 8684
rect 19868 8632 19898 8684
rect 19898 8632 19924 8684
rect 19628 8630 19684 8632
rect 19708 8630 19764 8632
rect 19788 8630 19844 8632
rect 19868 8630 19924 8632
rect 19628 7352 19684 7354
rect 19708 7352 19764 7354
rect 19788 7352 19844 7354
rect 19868 7352 19924 7354
rect 19628 7300 19654 7352
rect 19654 7300 19684 7352
rect 19708 7300 19718 7352
rect 19718 7300 19764 7352
rect 19788 7300 19834 7352
rect 19834 7300 19844 7352
rect 19868 7300 19898 7352
rect 19898 7300 19924 7352
rect 19628 7298 19684 7300
rect 19708 7298 19764 7300
rect 19788 7298 19844 7300
rect 19868 7298 19924 7300
rect 19628 6020 19684 6022
rect 19708 6020 19764 6022
rect 19788 6020 19844 6022
rect 19868 6020 19924 6022
rect 19628 5968 19654 6020
rect 19654 5968 19684 6020
rect 19708 5968 19718 6020
rect 19718 5968 19764 6020
rect 19788 5968 19834 6020
rect 19834 5968 19844 6020
rect 19868 5968 19898 6020
rect 19898 5968 19924 6020
rect 19628 5966 19684 5968
rect 19708 5966 19764 5968
rect 19788 5966 19844 5968
rect 19868 5966 19924 5968
rect 19628 4688 19684 4690
rect 19708 4688 19764 4690
rect 19788 4688 19844 4690
rect 19868 4688 19924 4690
rect 19628 4636 19654 4688
rect 19654 4636 19684 4688
rect 19708 4636 19718 4688
rect 19718 4636 19764 4688
rect 19788 4636 19834 4688
rect 19834 4636 19844 4688
rect 19868 4636 19898 4688
rect 19898 4636 19924 4688
rect 19628 4634 19684 4636
rect 19708 4634 19764 4636
rect 19788 4634 19844 4636
rect 19868 4634 19924 4636
rect 19628 3356 19684 3358
rect 19708 3356 19764 3358
rect 19788 3356 19844 3358
rect 19868 3356 19924 3358
rect 19628 3304 19654 3356
rect 19654 3304 19684 3356
rect 19708 3304 19718 3356
rect 19718 3304 19764 3356
rect 19788 3304 19834 3356
rect 19834 3304 19844 3356
rect 19868 3304 19898 3356
rect 19898 3304 19924 3356
rect 19628 3302 19684 3304
rect 19708 3302 19764 3304
rect 19788 3302 19844 3304
rect 19868 3302 19924 3304
rect 34988 57302 35044 57304
rect 35068 57302 35124 57304
rect 35148 57302 35204 57304
rect 35228 57302 35284 57304
rect 34988 57250 35014 57302
rect 35014 57250 35044 57302
rect 35068 57250 35078 57302
rect 35078 57250 35124 57302
rect 35148 57250 35194 57302
rect 35194 57250 35204 57302
rect 35228 57250 35258 57302
rect 35258 57250 35284 57302
rect 34988 57248 35044 57250
rect 35068 57248 35124 57250
rect 35148 57248 35204 57250
rect 35228 57248 35284 57250
rect 34988 55970 35044 55972
rect 35068 55970 35124 55972
rect 35148 55970 35204 55972
rect 35228 55970 35284 55972
rect 34988 55918 35014 55970
rect 35014 55918 35044 55970
rect 35068 55918 35078 55970
rect 35078 55918 35124 55970
rect 35148 55918 35194 55970
rect 35194 55918 35204 55970
rect 35228 55918 35258 55970
rect 35258 55918 35284 55970
rect 34988 55916 35044 55918
rect 35068 55916 35124 55918
rect 35148 55916 35204 55918
rect 35228 55916 35284 55918
rect 34988 54638 35044 54640
rect 35068 54638 35124 54640
rect 35148 54638 35204 54640
rect 35228 54638 35284 54640
rect 34988 54586 35014 54638
rect 35014 54586 35044 54638
rect 35068 54586 35078 54638
rect 35078 54586 35124 54638
rect 35148 54586 35194 54638
rect 35194 54586 35204 54638
rect 35228 54586 35258 54638
rect 35258 54586 35284 54638
rect 34988 54584 35044 54586
rect 35068 54584 35124 54586
rect 35148 54584 35204 54586
rect 35228 54584 35284 54586
rect 34988 53306 35044 53308
rect 35068 53306 35124 53308
rect 35148 53306 35204 53308
rect 35228 53306 35284 53308
rect 34988 53254 35014 53306
rect 35014 53254 35044 53306
rect 35068 53254 35078 53306
rect 35078 53254 35124 53306
rect 35148 53254 35194 53306
rect 35194 53254 35204 53306
rect 35228 53254 35258 53306
rect 35258 53254 35284 53306
rect 34988 53252 35044 53254
rect 35068 53252 35124 53254
rect 35148 53252 35204 53254
rect 35228 53252 35284 53254
rect 34988 51974 35044 51976
rect 35068 51974 35124 51976
rect 35148 51974 35204 51976
rect 35228 51974 35284 51976
rect 34988 51922 35014 51974
rect 35014 51922 35044 51974
rect 35068 51922 35078 51974
rect 35078 51922 35124 51974
rect 35148 51922 35194 51974
rect 35194 51922 35204 51974
rect 35228 51922 35258 51974
rect 35258 51922 35284 51974
rect 34988 51920 35044 51922
rect 35068 51920 35124 51922
rect 35148 51920 35204 51922
rect 35228 51920 35284 51922
rect 34988 50642 35044 50644
rect 35068 50642 35124 50644
rect 35148 50642 35204 50644
rect 35228 50642 35284 50644
rect 34988 50590 35014 50642
rect 35014 50590 35044 50642
rect 35068 50590 35078 50642
rect 35078 50590 35124 50642
rect 35148 50590 35194 50642
rect 35194 50590 35204 50642
rect 35228 50590 35258 50642
rect 35258 50590 35284 50642
rect 34988 50588 35044 50590
rect 35068 50588 35124 50590
rect 35148 50588 35204 50590
rect 35228 50588 35284 50590
rect 34988 49310 35044 49312
rect 35068 49310 35124 49312
rect 35148 49310 35204 49312
rect 35228 49310 35284 49312
rect 34988 49258 35014 49310
rect 35014 49258 35044 49310
rect 35068 49258 35078 49310
rect 35078 49258 35124 49310
rect 35148 49258 35194 49310
rect 35194 49258 35204 49310
rect 35228 49258 35258 49310
rect 35258 49258 35284 49310
rect 34988 49256 35044 49258
rect 35068 49256 35124 49258
rect 35148 49256 35204 49258
rect 35228 49256 35284 49258
rect 34988 47978 35044 47980
rect 35068 47978 35124 47980
rect 35148 47978 35204 47980
rect 35228 47978 35284 47980
rect 34988 47926 35014 47978
rect 35014 47926 35044 47978
rect 35068 47926 35078 47978
rect 35078 47926 35124 47978
rect 35148 47926 35194 47978
rect 35194 47926 35204 47978
rect 35228 47926 35258 47978
rect 35258 47926 35284 47978
rect 34988 47924 35044 47926
rect 35068 47924 35124 47926
rect 35148 47924 35204 47926
rect 35228 47924 35284 47926
rect 34988 46646 35044 46648
rect 35068 46646 35124 46648
rect 35148 46646 35204 46648
rect 35228 46646 35284 46648
rect 34988 46594 35014 46646
rect 35014 46594 35044 46646
rect 35068 46594 35078 46646
rect 35078 46594 35124 46646
rect 35148 46594 35194 46646
rect 35194 46594 35204 46646
rect 35228 46594 35258 46646
rect 35258 46594 35284 46646
rect 34988 46592 35044 46594
rect 35068 46592 35124 46594
rect 35148 46592 35204 46594
rect 35228 46592 35284 46594
rect 34988 45314 35044 45316
rect 35068 45314 35124 45316
rect 35148 45314 35204 45316
rect 35228 45314 35284 45316
rect 34988 45262 35014 45314
rect 35014 45262 35044 45314
rect 35068 45262 35078 45314
rect 35078 45262 35124 45314
rect 35148 45262 35194 45314
rect 35194 45262 35204 45314
rect 35228 45262 35258 45314
rect 35258 45262 35284 45314
rect 34988 45260 35044 45262
rect 35068 45260 35124 45262
rect 35148 45260 35204 45262
rect 35228 45260 35284 45262
rect 34988 43982 35044 43984
rect 35068 43982 35124 43984
rect 35148 43982 35204 43984
rect 35228 43982 35284 43984
rect 34988 43930 35014 43982
rect 35014 43930 35044 43982
rect 35068 43930 35078 43982
rect 35078 43930 35124 43982
rect 35148 43930 35194 43982
rect 35194 43930 35204 43982
rect 35228 43930 35258 43982
rect 35258 43930 35284 43982
rect 34988 43928 35044 43930
rect 35068 43928 35124 43930
rect 35148 43928 35204 43930
rect 35228 43928 35284 43930
rect 34988 42650 35044 42652
rect 35068 42650 35124 42652
rect 35148 42650 35204 42652
rect 35228 42650 35284 42652
rect 34988 42598 35014 42650
rect 35014 42598 35044 42650
rect 35068 42598 35078 42650
rect 35078 42598 35124 42650
rect 35148 42598 35194 42650
rect 35194 42598 35204 42650
rect 35228 42598 35258 42650
rect 35258 42598 35284 42650
rect 34988 42596 35044 42598
rect 35068 42596 35124 42598
rect 35148 42596 35204 42598
rect 35228 42596 35284 42598
rect 34988 41318 35044 41320
rect 35068 41318 35124 41320
rect 35148 41318 35204 41320
rect 35228 41318 35284 41320
rect 34988 41266 35014 41318
rect 35014 41266 35044 41318
rect 35068 41266 35078 41318
rect 35078 41266 35124 41318
rect 35148 41266 35194 41318
rect 35194 41266 35204 41318
rect 35228 41266 35258 41318
rect 35258 41266 35284 41318
rect 34988 41264 35044 41266
rect 35068 41264 35124 41266
rect 35148 41264 35204 41266
rect 35228 41264 35284 41266
rect 34988 39986 35044 39988
rect 35068 39986 35124 39988
rect 35148 39986 35204 39988
rect 35228 39986 35284 39988
rect 34988 39934 35014 39986
rect 35014 39934 35044 39986
rect 35068 39934 35078 39986
rect 35078 39934 35124 39986
rect 35148 39934 35194 39986
rect 35194 39934 35204 39986
rect 35228 39934 35258 39986
rect 35258 39934 35284 39986
rect 34988 39932 35044 39934
rect 35068 39932 35124 39934
rect 35148 39932 35204 39934
rect 35228 39932 35284 39934
rect 34988 38654 35044 38656
rect 35068 38654 35124 38656
rect 35148 38654 35204 38656
rect 35228 38654 35284 38656
rect 34988 38602 35014 38654
rect 35014 38602 35044 38654
rect 35068 38602 35078 38654
rect 35078 38602 35124 38654
rect 35148 38602 35194 38654
rect 35194 38602 35204 38654
rect 35228 38602 35258 38654
rect 35258 38602 35284 38654
rect 34988 38600 35044 38602
rect 35068 38600 35124 38602
rect 35148 38600 35204 38602
rect 35228 38600 35284 38602
rect 34988 37322 35044 37324
rect 35068 37322 35124 37324
rect 35148 37322 35204 37324
rect 35228 37322 35284 37324
rect 34988 37270 35014 37322
rect 35014 37270 35044 37322
rect 35068 37270 35078 37322
rect 35078 37270 35124 37322
rect 35148 37270 35194 37322
rect 35194 37270 35204 37322
rect 35228 37270 35258 37322
rect 35258 37270 35284 37322
rect 34988 37268 35044 37270
rect 35068 37268 35124 37270
rect 35148 37268 35204 37270
rect 35228 37268 35284 37270
rect 34988 35990 35044 35992
rect 35068 35990 35124 35992
rect 35148 35990 35204 35992
rect 35228 35990 35284 35992
rect 34988 35938 35014 35990
rect 35014 35938 35044 35990
rect 35068 35938 35078 35990
rect 35078 35938 35124 35990
rect 35148 35938 35194 35990
rect 35194 35938 35204 35990
rect 35228 35938 35258 35990
rect 35258 35938 35284 35990
rect 34988 35936 35044 35938
rect 35068 35936 35124 35938
rect 35148 35936 35204 35938
rect 35228 35936 35284 35938
rect 34988 34658 35044 34660
rect 35068 34658 35124 34660
rect 35148 34658 35204 34660
rect 35228 34658 35284 34660
rect 34988 34606 35014 34658
rect 35014 34606 35044 34658
rect 35068 34606 35078 34658
rect 35078 34606 35124 34658
rect 35148 34606 35194 34658
rect 35194 34606 35204 34658
rect 35228 34606 35258 34658
rect 35258 34606 35284 34658
rect 34988 34604 35044 34606
rect 35068 34604 35124 34606
rect 35148 34604 35204 34606
rect 35228 34604 35284 34606
rect 34988 33326 35044 33328
rect 35068 33326 35124 33328
rect 35148 33326 35204 33328
rect 35228 33326 35284 33328
rect 34988 33274 35014 33326
rect 35014 33274 35044 33326
rect 35068 33274 35078 33326
rect 35078 33274 35124 33326
rect 35148 33274 35194 33326
rect 35194 33274 35204 33326
rect 35228 33274 35258 33326
rect 35258 33274 35284 33326
rect 34988 33272 35044 33274
rect 35068 33272 35124 33274
rect 35148 33272 35204 33274
rect 35228 33272 35284 33274
rect 34988 31994 35044 31996
rect 35068 31994 35124 31996
rect 35148 31994 35204 31996
rect 35228 31994 35284 31996
rect 34988 31942 35014 31994
rect 35014 31942 35044 31994
rect 35068 31942 35078 31994
rect 35078 31942 35124 31994
rect 35148 31942 35194 31994
rect 35194 31942 35204 31994
rect 35228 31942 35258 31994
rect 35258 31942 35284 31994
rect 34988 31940 35044 31942
rect 35068 31940 35124 31942
rect 35148 31940 35204 31942
rect 35228 31940 35284 31942
rect 34988 30662 35044 30664
rect 35068 30662 35124 30664
rect 35148 30662 35204 30664
rect 35228 30662 35284 30664
rect 34988 30610 35014 30662
rect 35014 30610 35044 30662
rect 35068 30610 35078 30662
rect 35078 30610 35124 30662
rect 35148 30610 35194 30662
rect 35194 30610 35204 30662
rect 35228 30610 35258 30662
rect 35258 30610 35284 30662
rect 34988 30608 35044 30610
rect 35068 30608 35124 30610
rect 35148 30608 35204 30610
rect 35228 30608 35284 30610
rect 34988 29330 35044 29332
rect 35068 29330 35124 29332
rect 35148 29330 35204 29332
rect 35228 29330 35284 29332
rect 34988 29278 35014 29330
rect 35014 29278 35044 29330
rect 35068 29278 35078 29330
rect 35078 29278 35124 29330
rect 35148 29278 35194 29330
rect 35194 29278 35204 29330
rect 35228 29278 35258 29330
rect 35258 29278 35284 29330
rect 34988 29276 35044 29278
rect 35068 29276 35124 29278
rect 35148 29276 35204 29278
rect 35228 29276 35284 29278
rect 34988 27998 35044 28000
rect 35068 27998 35124 28000
rect 35148 27998 35204 28000
rect 35228 27998 35284 28000
rect 34988 27946 35014 27998
rect 35014 27946 35044 27998
rect 35068 27946 35078 27998
rect 35078 27946 35124 27998
rect 35148 27946 35194 27998
rect 35194 27946 35204 27998
rect 35228 27946 35258 27998
rect 35258 27946 35284 27998
rect 34988 27944 35044 27946
rect 35068 27944 35124 27946
rect 35148 27944 35204 27946
rect 35228 27944 35284 27946
rect 34988 26666 35044 26668
rect 35068 26666 35124 26668
rect 35148 26666 35204 26668
rect 35228 26666 35284 26668
rect 34988 26614 35014 26666
rect 35014 26614 35044 26666
rect 35068 26614 35078 26666
rect 35078 26614 35124 26666
rect 35148 26614 35194 26666
rect 35194 26614 35204 26666
rect 35228 26614 35258 26666
rect 35258 26614 35284 26666
rect 34988 26612 35044 26614
rect 35068 26612 35124 26614
rect 35148 26612 35204 26614
rect 35228 26612 35284 26614
rect 34988 25334 35044 25336
rect 35068 25334 35124 25336
rect 35148 25334 35204 25336
rect 35228 25334 35284 25336
rect 34988 25282 35014 25334
rect 35014 25282 35044 25334
rect 35068 25282 35078 25334
rect 35078 25282 35124 25334
rect 35148 25282 35194 25334
rect 35194 25282 35204 25334
rect 35228 25282 35258 25334
rect 35258 25282 35284 25334
rect 34988 25280 35044 25282
rect 35068 25280 35124 25282
rect 35148 25280 35204 25282
rect 35228 25280 35284 25282
rect 34988 24002 35044 24004
rect 35068 24002 35124 24004
rect 35148 24002 35204 24004
rect 35228 24002 35284 24004
rect 34988 23950 35014 24002
rect 35014 23950 35044 24002
rect 35068 23950 35078 24002
rect 35078 23950 35124 24002
rect 35148 23950 35194 24002
rect 35194 23950 35204 24002
rect 35228 23950 35258 24002
rect 35258 23950 35284 24002
rect 34988 23948 35044 23950
rect 35068 23948 35124 23950
rect 35148 23948 35204 23950
rect 35228 23948 35284 23950
rect 34988 22670 35044 22672
rect 35068 22670 35124 22672
rect 35148 22670 35204 22672
rect 35228 22670 35284 22672
rect 34988 22618 35014 22670
rect 35014 22618 35044 22670
rect 35068 22618 35078 22670
rect 35078 22618 35124 22670
rect 35148 22618 35194 22670
rect 35194 22618 35204 22670
rect 35228 22618 35258 22670
rect 35258 22618 35284 22670
rect 34988 22616 35044 22618
rect 35068 22616 35124 22618
rect 35148 22616 35204 22618
rect 35228 22616 35284 22618
rect 34988 21338 35044 21340
rect 35068 21338 35124 21340
rect 35148 21338 35204 21340
rect 35228 21338 35284 21340
rect 34988 21286 35014 21338
rect 35014 21286 35044 21338
rect 35068 21286 35078 21338
rect 35078 21286 35124 21338
rect 35148 21286 35194 21338
rect 35194 21286 35204 21338
rect 35228 21286 35258 21338
rect 35258 21286 35284 21338
rect 34988 21284 35044 21286
rect 35068 21284 35124 21286
rect 35148 21284 35204 21286
rect 35228 21284 35284 21286
rect 34988 20006 35044 20008
rect 35068 20006 35124 20008
rect 35148 20006 35204 20008
rect 35228 20006 35284 20008
rect 34988 19954 35014 20006
rect 35014 19954 35044 20006
rect 35068 19954 35078 20006
rect 35078 19954 35124 20006
rect 35148 19954 35194 20006
rect 35194 19954 35204 20006
rect 35228 19954 35258 20006
rect 35258 19954 35284 20006
rect 34988 19952 35044 19954
rect 35068 19952 35124 19954
rect 35148 19952 35204 19954
rect 35228 19952 35284 19954
rect 34988 18674 35044 18676
rect 35068 18674 35124 18676
rect 35148 18674 35204 18676
rect 35228 18674 35284 18676
rect 34988 18622 35014 18674
rect 35014 18622 35044 18674
rect 35068 18622 35078 18674
rect 35078 18622 35124 18674
rect 35148 18622 35194 18674
rect 35194 18622 35204 18674
rect 35228 18622 35258 18674
rect 35258 18622 35284 18674
rect 34988 18620 35044 18622
rect 35068 18620 35124 18622
rect 35148 18620 35204 18622
rect 35228 18620 35284 18622
rect 34988 17342 35044 17344
rect 35068 17342 35124 17344
rect 35148 17342 35204 17344
rect 35228 17342 35284 17344
rect 34988 17290 35014 17342
rect 35014 17290 35044 17342
rect 35068 17290 35078 17342
rect 35078 17290 35124 17342
rect 35148 17290 35194 17342
rect 35194 17290 35204 17342
rect 35228 17290 35258 17342
rect 35258 17290 35284 17342
rect 34988 17288 35044 17290
rect 35068 17288 35124 17290
rect 35148 17288 35204 17290
rect 35228 17288 35284 17290
rect 34988 16010 35044 16012
rect 35068 16010 35124 16012
rect 35148 16010 35204 16012
rect 35228 16010 35284 16012
rect 34988 15958 35014 16010
rect 35014 15958 35044 16010
rect 35068 15958 35078 16010
rect 35078 15958 35124 16010
rect 35148 15958 35194 16010
rect 35194 15958 35204 16010
rect 35228 15958 35258 16010
rect 35258 15958 35284 16010
rect 34988 15956 35044 15958
rect 35068 15956 35124 15958
rect 35148 15956 35204 15958
rect 35228 15956 35284 15958
rect 34988 14678 35044 14680
rect 35068 14678 35124 14680
rect 35148 14678 35204 14680
rect 35228 14678 35284 14680
rect 34988 14626 35014 14678
rect 35014 14626 35044 14678
rect 35068 14626 35078 14678
rect 35078 14626 35124 14678
rect 35148 14626 35194 14678
rect 35194 14626 35204 14678
rect 35228 14626 35258 14678
rect 35258 14626 35284 14678
rect 34988 14624 35044 14626
rect 35068 14624 35124 14626
rect 35148 14624 35204 14626
rect 35228 14624 35284 14626
rect 34988 13346 35044 13348
rect 35068 13346 35124 13348
rect 35148 13346 35204 13348
rect 35228 13346 35284 13348
rect 34988 13294 35014 13346
rect 35014 13294 35044 13346
rect 35068 13294 35078 13346
rect 35078 13294 35124 13346
rect 35148 13294 35194 13346
rect 35194 13294 35204 13346
rect 35228 13294 35258 13346
rect 35258 13294 35284 13346
rect 34988 13292 35044 13294
rect 35068 13292 35124 13294
rect 35148 13292 35204 13294
rect 35228 13292 35284 13294
rect 34988 12014 35044 12016
rect 35068 12014 35124 12016
rect 35148 12014 35204 12016
rect 35228 12014 35284 12016
rect 34988 11962 35014 12014
rect 35014 11962 35044 12014
rect 35068 11962 35078 12014
rect 35078 11962 35124 12014
rect 35148 11962 35194 12014
rect 35194 11962 35204 12014
rect 35228 11962 35258 12014
rect 35258 11962 35284 12014
rect 34988 11960 35044 11962
rect 35068 11960 35124 11962
rect 35148 11960 35204 11962
rect 35228 11960 35284 11962
rect 34988 10682 35044 10684
rect 35068 10682 35124 10684
rect 35148 10682 35204 10684
rect 35228 10682 35284 10684
rect 34988 10630 35014 10682
rect 35014 10630 35044 10682
rect 35068 10630 35078 10682
rect 35078 10630 35124 10682
rect 35148 10630 35194 10682
rect 35194 10630 35204 10682
rect 35228 10630 35258 10682
rect 35258 10630 35284 10682
rect 34988 10628 35044 10630
rect 35068 10628 35124 10630
rect 35148 10628 35204 10630
rect 35228 10628 35284 10630
rect 34988 9350 35044 9352
rect 35068 9350 35124 9352
rect 35148 9350 35204 9352
rect 35228 9350 35284 9352
rect 34988 9298 35014 9350
rect 35014 9298 35044 9350
rect 35068 9298 35078 9350
rect 35078 9298 35124 9350
rect 35148 9298 35194 9350
rect 35194 9298 35204 9350
rect 35228 9298 35258 9350
rect 35258 9298 35284 9350
rect 34988 9296 35044 9298
rect 35068 9296 35124 9298
rect 35148 9296 35204 9298
rect 35228 9296 35284 9298
rect 34988 8018 35044 8020
rect 35068 8018 35124 8020
rect 35148 8018 35204 8020
rect 35228 8018 35284 8020
rect 34988 7966 35014 8018
rect 35014 7966 35044 8018
rect 35068 7966 35078 8018
rect 35078 7966 35124 8018
rect 35148 7966 35194 8018
rect 35194 7966 35204 8018
rect 35228 7966 35258 8018
rect 35258 7966 35284 8018
rect 34988 7964 35044 7966
rect 35068 7964 35124 7966
rect 35148 7964 35204 7966
rect 35228 7964 35284 7966
rect 34988 6686 35044 6688
rect 35068 6686 35124 6688
rect 35148 6686 35204 6688
rect 35228 6686 35284 6688
rect 34988 6634 35014 6686
rect 35014 6634 35044 6686
rect 35068 6634 35078 6686
rect 35078 6634 35124 6686
rect 35148 6634 35194 6686
rect 35194 6634 35204 6686
rect 35228 6634 35258 6686
rect 35258 6634 35284 6686
rect 34988 6632 35044 6634
rect 35068 6632 35124 6634
rect 35148 6632 35204 6634
rect 35228 6632 35284 6634
rect 34988 5354 35044 5356
rect 35068 5354 35124 5356
rect 35148 5354 35204 5356
rect 35228 5354 35284 5356
rect 34988 5302 35014 5354
rect 35014 5302 35044 5354
rect 35068 5302 35078 5354
rect 35078 5302 35124 5354
rect 35148 5302 35194 5354
rect 35194 5302 35204 5354
rect 35228 5302 35258 5354
rect 35258 5302 35284 5354
rect 34988 5300 35044 5302
rect 35068 5300 35124 5302
rect 35148 5300 35204 5302
rect 35228 5300 35284 5302
rect 34988 4022 35044 4024
rect 35068 4022 35124 4024
rect 35148 4022 35204 4024
rect 35228 4022 35284 4024
rect 34988 3970 35014 4022
rect 35014 3970 35044 4022
rect 35068 3970 35078 4022
rect 35078 3970 35124 4022
rect 35148 3970 35194 4022
rect 35194 3970 35204 4022
rect 35228 3970 35258 4022
rect 35258 3970 35284 4022
rect 34988 3968 35044 3970
rect 35068 3968 35124 3970
rect 35148 3968 35204 3970
rect 35228 3968 35284 3970
rect 34988 2690 35044 2692
rect 35068 2690 35124 2692
rect 35148 2690 35204 2692
rect 35228 2690 35284 2692
rect 34988 2638 35014 2690
rect 35014 2638 35044 2690
rect 35068 2638 35078 2690
rect 35078 2638 35124 2690
rect 35148 2638 35194 2690
rect 35194 2638 35204 2690
rect 35228 2638 35258 2690
rect 35258 2638 35284 2690
rect 34988 2636 35044 2638
rect 35068 2636 35124 2638
rect 35148 2636 35204 2638
rect 35228 2636 35284 2638
rect 41780 3006 41836 3062
rect 44372 3006 44428 3062
rect 50348 56636 50404 56638
rect 50428 56636 50484 56638
rect 50508 56636 50564 56638
rect 50588 56636 50644 56638
rect 50348 56584 50374 56636
rect 50374 56584 50404 56636
rect 50428 56584 50438 56636
rect 50438 56584 50484 56636
rect 50508 56584 50554 56636
rect 50554 56584 50564 56636
rect 50588 56584 50618 56636
rect 50618 56584 50644 56636
rect 50348 56582 50404 56584
rect 50428 56582 50484 56584
rect 50508 56582 50564 56584
rect 50588 56582 50644 56584
rect 50348 55304 50404 55306
rect 50428 55304 50484 55306
rect 50508 55304 50564 55306
rect 50588 55304 50644 55306
rect 50348 55252 50374 55304
rect 50374 55252 50404 55304
rect 50428 55252 50438 55304
rect 50438 55252 50484 55304
rect 50508 55252 50554 55304
rect 50554 55252 50564 55304
rect 50588 55252 50618 55304
rect 50618 55252 50644 55304
rect 50348 55250 50404 55252
rect 50428 55250 50484 55252
rect 50508 55250 50564 55252
rect 50588 55250 50644 55252
rect 50348 53972 50404 53974
rect 50428 53972 50484 53974
rect 50508 53972 50564 53974
rect 50588 53972 50644 53974
rect 50348 53920 50374 53972
rect 50374 53920 50404 53972
rect 50428 53920 50438 53972
rect 50438 53920 50484 53972
rect 50508 53920 50554 53972
rect 50554 53920 50564 53972
rect 50588 53920 50618 53972
rect 50618 53920 50644 53972
rect 50348 53918 50404 53920
rect 50428 53918 50484 53920
rect 50508 53918 50564 53920
rect 50588 53918 50644 53920
rect 50348 52640 50404 52642
rect 50428 52640 50484 52642
rect 50508 52640 50564 52642
rect 50588 52640 50644 52642
rect 50348 52588 50374 52640
rect 50374 52588 50404 52640
rect 50428 52588 50438 52640
rect 50438 52588 50484 52640
rect 50508 52588 50554 52640
rect 50554 52588 50564 52640
rect 50588 52588 50618 52640
rect 50618 52588 50644 52640
rect 50348 52586 50404 52588
rect 50428 52586 50484 52588
rect 50508 52586 50564 52588
rect 50588 52586 50644 52588
rect 50348 51308 50404 51310
rect 50428 51308 50484 51310
rect 50508 51308 50564 51310
rect 50588 51308 50644 51310
rect 50348 51256 50374 51308
rect 50374 51256 50404 51308
rect 50428 51256 50438 51308
rect 50438 51256 50484 51308
rect 50508 51256 50554 51308
rect 50554 51256 50564 51308
rect 50588 51256 50618 51308
rect 50618 51256 50644 51308
rect 50348 51254 50404 51256
rect 50428 51254 50484 51256
rect 50508 51254 50564 51256
rect 50588 51254 50644 51256
rect 50348 49976 50404 49978
rect 50428 49976 50484 49978
rect 50508 49976 50564 49978
rect 50588 49976 50644 49978
rect 50348 49924 50374 49976
rect 50374 49924 50404 49976
rect 50428 49924 50438 49976
rect 50438 49924 50484 49976
rect 50508 49924 50554 49976
rect 50554 49924 50564 49976
rect 50588 49924 50618 49976
rect 50618 49924 50644 49976
rect 50348 49922 50404 49924
rect 50428 49922 50484 49924
rect 50508 49922 50564 49924
rect 50588 49922 50644 49924
rect 50348 48644 50404 48646
rect 50428 48644 50484 48646
rect 50508 48644 50564 48646
rect 50588 48644 50644 48646
rect 50348 48592 50374 48644
rect 50374 48592 50404 48644
rect 50428 48592 50438 48644
rect 50438 48592 50484 48644
rect 50508 48592 50554 48644
rect 50554 48592 50564 48644
rect 50588 48592 50618 48644
rect 50618 48592 50644 48644
rect 50348 48590 50404 48592
rect 50428 48590 50484 48592
rect 50508 48590 50564 48592
rect 50588 48590 50644 48592
rect 50348 47312 50404 47314
rect 50428 47312 50484 47314
rect 50508 47312 50564 47314
rect 50588 47312 50644 47314
rect 50348 47260 50374 47312
rect 50374 47260 50404 47312
rect 50428 47260 50438 47312
rect 50438 47260 50484 47312
rect 50508 47260 50554 47312
rect 50554 47260 50564 47312
rect 50588 47260 50618 47312
rect 50618 47260 50644 47312
rect 50348 47258 50404 47260
rect 50428 47258 50484 47260
rect 50508 47258 50564 47260
rect 50588 47258 50644 47260
rect 50348 45980 50404 45982
rect 50428 45980 50484 45982
rect 50508 45980 50564 45982
rect 50588 45980 50644 45982
rect 50348 45928 50374 45980
rect 50374 45928 50404 45980
rect 50428 45928 50438 45980
rect 50438 45928 50484 45980
rect 50508 45928 50554 45980
rect 50554 45928 50564 45980
rect 50588 45928 50618 45980
rect 50618 45928 50644 45980
rect 50348 45926 50404 45928
rect 50428 45926 50484 45928
rect 50508 45926 50564 45928
rect 50588 45926 50644 45928
rect 50348 44648 50404 44650
rect 50428 44648 50484 44650
rect 50508 44648 50564 44650
rect 50588 44648 50644 44650
rect 50348 44596 50374 44648
rect 50374 44596 50404 44648
rect 50428 44596 50438 44648
rect 50438 44596 50484 44648
rect 50508 44596 50554 44648
rect 50554 44596 50564 44648
rect 50588 44596 50618 44648
rect 50618 44596 50644 44648
rect 50348 44594 50404 44596
rect 50428 44594 50484 44596
rect 50508 44594 50564 44596
rect 50588 44594 50644 44596
rect 50348 43316 50404 43318
rect 50428 43316 50484 43318
rect 50508 43316 50564 43318
rect 50588 43316 50644 43318
rect 50348 43264 50374 43316
rect 50374 43264 50404 43316
rect 50428 43264 50438 43316
rect 50438 43264 50484 43316
rect 50508 43264 50554 43316
rect 50554 43264 50564 43316
rect 50588 43264 50618 43316
rect 50618 43264 50644 43316
rect 50348 43262 50404 43264
rect 50428 43262 50484 43264
rect 50508 43262 50564 43264
rect 50588 43262 50644 43264
rect 50348 41984 50404 41986
rect 50428 41984 50484 41986
rect 50508 41984 50564 41986
rect 50588 41984 50644 41986
rect 50348 41932 50374 41984
rect 50374 41932 50404 41984
rect 50428 41932 50438 41984
rect 50438 41932 50484 41984
rect 50508 41932 50554 41984
rect 50554 41932 50564 41984
rect 50588 41932 50618 41984
rect 50618 41932 50644 41984
rect 50348 41930 50404 41932
rect 50428 41930 50484 41932
rect 50508 41930 50564 41932
rect 50588 41930 50644 41932
rect 50348 40652 50404 40654
rect 50428 40652 50484 40654
rect 50508 40652 50564 40654
rect 50588 40652 50644 40654
rect 50348 40600 50374 40652
rect 50374 40600 50404 40652
rect 50428 40600 50438 40652
rect 50438 40600 50484 40652
rect 50508 40600 50554 40652
rect 50554 40600 50564 40652
rect 50588 40600 50618 40652
rect 50618 40600 50644 40652
rect 50348 40598 50404 40600
rect 50428 40598 50484 40600
rect 50508 40598 50564 40600
rect 50588 40598 50644 40600
rect 50348 39320 50404 39322
rect 50428 39320 50484 39322
rect 50508 39320 50564 39322
rect 50588 39320 50644 39322
rect 50348 39268 50374 39320
rect 50374 39268 50404 39320
rect 50428 39268 50438 39320
rect 50438 39268 50484 39320
rect 50508 39268 50554 39320
rect 50554 39268 50564 39320
rect 50588 39268 50618 39320
rect 50618 39268 50644 39320
rect 50348 39266 50404 39268
rect 50428 39266 50484 39268
rect 50508 39266 50564 39268
rect 50588 39266 50644 39268
rect 50348 37988 50404 37990
rect 50428 37988 50484 37990
rect 50508 37988 50564 37990
rect 50588 37988 50644 37990
rect 50348 37936 50374 37988
rect 50374 37936 50404 37988
rect 50428 37936 50438 37988
rect 50438 37936 50484 37988
rect 50508 37936 50554 37988
rect 50554 37936 50564 37988
rect 50588 37936 50618 37988
rect 50618 37936 50644 37988
rect 50348 37934 50404 37936
rect 50428 37934 50484 37936
rect 50508 37934 50564 37936
rect 50588 37934 50644 37936
rect 50348 36656 50404 36658
rect 50428 36656 50484 36658
rect 50508 36656 50564 36658
rect 50588 36656 50644 36658
rect 50348 36604 50374 36656
rect 50374 36604 50404 36656
rect 50428 36604 50438 36656
rect 50438 36604 50484 36656
rect 50508 36604 50554 36656
rect 50554 36604 50564 36656
rect 50588 36604 50618 36656
rect 50618 36604 50644 36656
rect 50348 36602 50404 36604
rect 50428 36602 50484 36604
rect 50508 36602 50564 36604
rect 50588 36602 50644 36604
rect 50348 35324 50404 35326
rect 50428 35324 50484 35326
rect 50508 35324 50564 35326
rect 50588 35324 50644 35326
rect 50348 35272 50374 35324
rect 50374 35272 50404 35324
rect 50428 35272 50438 35324
rect 50438 35272 50484 35324
rect 50508 35272 50554 35324
rect 50554 35272 50564 35324
rect 50588 35272 50618 35324
rect 50618 35272 50644 35324
rect 50348 35270 50404 35272
rect 50428 35270 50484 35272
rect 50508 35270 50564 35272
rect 50588 35270 50644 35272
rect 50348 33992 50404 33994
rect 50428 33992 50484 33994
rect 50508 33992 50564 33994
rect 50588 33992 50644 33994
rect 50348 33940 50374 33992
rect 50374 33940 50404 33992
rect 50428 33940 50438 33992
rect 50438 33940 50484 33992
rect 50508 33940 50554 33992
rect 50554 33940 50564 33992
rect 50588 33940 50618 33992
rect 50618 33940 50644 33992
rect 50348 33938 50404 33940
rect 50428 33938 50484 33940
rect 50508 33938 50564 33940
rect 50588 33938 50644 33940
rect 50348 32660 50404 32662
rect 50428 32660 50484 32662
rect 50508 32660 50564 32662
rect 50588 32660 50644 32662
rect 50348 32608 50374 32660
rect 50374 32608 50404 32660
rect 50428 32608 50438 32660
rect 50438 32608 50484 32660
rect 50508 32608 50554 32660
rect 50554 32608 50564 32660
rect 50588 32608 50618 32660
rect 50618 32608 50644 32660
rect 50348 32606 50404 32608
rect 50428 32606 50484 32608
rect 50508 32606 50564 32608
rect 50588 32606 50644 32608
rect 50348 31328 50404 31330
rect 50428 31328 50484 31330
rect 50508 31328 50564 31330
rect 50588 31328 50644 31330
rect 50348 31276 50374 31328
rect 50374 31276 50404 31328
rect 50428 31276 50438 31328
rect 50438 31276 50484 31328
rect 50508 31276 50554 31328
rect 50554 31276 50564 31328
rect 50588 31276 50618 31328
rect 50618 31276 50644 31328
rect 50348 31274 50404 31276
rect 50428 31274 50484 31276
rect 50508 31274 50564 31276
rect 50588 31274 50644 31276
rect 50348 29996 50404 29998
rect 50428 29996 50484 29998
rect 50508 29996 50564 29998
rect 50588 29996 50644 29998
rect 50348 29944 50374 29996
rect 50374 29944 50404 29996
rect 50428 29944 50438 29996
rect 50438 29944 50484 29996
rect 50508 29944 50554 29996
rect 50554 29944 50564 29996
rect 50588 29944 50618 29996
rect 50618 29944 50644 29996
rect 50348 29942 50404 29944
rect 50428 29942 50484 29944
rect 50508 29942 50564 29944
rect 50588 29942 50644 29944
rect 50348 28664 50404 28666
rect 50428 28664 50484 28666
rect 50508 28664 50564 28666
rect 50588 28664 50644 28666
rect 50348 28612 50374 28664
rect 50374 28612 50404 28664
rect 50428 28612 50438 28664
rect 50438 28612 50484 28664
rect 50508 28612 50554 28664
rect 50554 28612 50564 28664
rect 50588 28612 50618 28664
rect 50618 28612 50644 28664
rect 50348 28610 50404 28612
rect 50428 28610 50484 28612
rect 50508 28610 50564 28612
rect 50588 28610 50644 28612
rect 50348 27332 50404 27334
rect 50428 27332 50484 27334
rect 50508 27332 50564 27334
rect 50588 27332 50644 27334
rect 50348 27280 50374 27332
rect 50374 27280 50404 27332
rect 50428 27280 50438 27332
rect 50438 27280 50484 27332
rect 50508 27280 50554 27332
rect 50554 27280 50564 27332
rect 50588 27280 50618 27332
rect 50618 27280 50644 27332
rect 50348 27278 50404 27280
rect 50428 27278 50484 27280
rect 50508 27278 50564 27280
rect 50588 27278 50644 27280
rect 50348 26000 50404 26002
rect 50428 26000 50484 26002
rect 50508 26000 50564 26002
rect 50588 26000 50644 26002
rect 50348 25948 50374 26000
rect 50374 25948 50404 26000
rect 50428 25948 50438 26000
rect 50438 25948 50484 26000
rect 50508 25948 50554 26000
rect 50554 25948 50564 26000
rect 50588 25948 50618 26000
rect 50618 25948 50644 26000
rect 50348 25946 50404 25948
rect 50428 25946 50484 25948
rect 50508 25946 50564 25948
rect 50588 25946 50644 25948
rect 50348 24668 50404 24670
rect 50428 24668 50484 24670
rect 50508 24668 50564 24670
rect 50588 24668 50644 24670
rect 50348 24616 50374 24668
rect 50374 24616 50404 24668
rect 50428 24616 50438 24668
rect 50438 24616 50484 24668
rect 50508 24616 50554 24668
rect 50554 24616 50564 24668
rect 50588 24616 50618 24668
rect 50618 24616 50644 24668
rect 50348 24614 50404 24616
rect 50428 24614 50484 24616
rect 50508 24614 50564 24616
rect 50588 24614 50644 24616
rect 50348 23336 50404 23338
rect 50428 23336 50484 23338
rect 50508 23336 50564 23338
rect 50588 23336 50644 23338
rect 50348 23284 50374 23336
rect 50374 23284 50404 23336
rect 50428 23284 50438 23336
rect 50438 23284 50484 23336
rect 50508 23284 50554 23336
rect 50554 23284 50564 23336
rect 50588 23284 50618 23336
rect 50618 23284 50644 23336
rect 50348 23282 50404 23284
rect 50428 23282 50484 23284
rect 50508 23282 50564 23284
rect 50588 23282 50644 23284
rect 50348 22004 50404 22006
rect 50428 22004 50484 22006
rect 50508 22004 50564 22006
rect 50588 22004 50644 22006
rect 50348 21952 50374 22004
rect 50374 21952 50404 22004
rect 50428 21952 50438 22004
rect 50438 21952 50484 22004
rect 50508 21952 50554 22004
rect 50554 21952 50564 22004
rect 50588 21952 50618 22004
rect 50618 21952 50644 22004
rect 50348 21950 50404 21952
rect 50428 21950 50484 21952
rect 50508 21950 50564 21952
rect 50588 21950 50644 21952
rect 50348 20672 50404 20674
rect 50428 20672 50484 20674
rect 50508 20672 50564 20674
rect 50588 20672 50644 20674
rect 50348 20620 50374 20672
rect 50374 20620 50404 20672
rect 50428 20620 50438 20672
rect 50438 20620 50484 20672
rect 50508 20620 50554 20672
rect 50554 20620 50564 20672
rect 50588 20620 50618 20672
rect 50618 20620 50644 20672
rect 50348 20618 50404 20620
rect 50428 20618 50484 20620
rect 50508 20618 50564 20620
rect 50588 20618 50644 20620
rect 50348 19340 50404 19342
rect 50428 19340 50484 19342
rect 50508 19340 50564 19342
rect 50588 19340 50644 19342
rect 50348 19288 50374 19340
rect 50374 19288 50404 19340
rect 50428 19288 50438 19340
rect 50438 19288 50484 19340
rect 50508 19288 50554 19340
rect 50554 19288 50564 19340
rect 50588 19288 50618 19340
rect 50618 19288 50644 19340
rect 50348 19286 50404 19288
rect 50428 19286 50484 19288
rect 50508 19286 50564 19288
rect 50588 19286 50644 19288
rect 50348 18008 50404 18010
rect 50428 18008 50484 18010
rect 50508 18008 50564 18010
rect 50588 18008 50644 18010
rect 50348 17956 50374 18008
rect 50374 17956 50404 18008
rect 50428 17956 50438 18008
rect 50438 17956 50484 18008
rect 50508 17956 50554 18008
rect 50554 17956 50564 18008
rect 50588 17956 50618 18008
rect 50618 17956 50644 18008
rect 50348 17954 50404 17956
rect 50428 17954 50484 17956
rect 50508 17954 50564 17956
rect 50588 17954 50644 17956
rect 50348 16676 50404 16678
rect 50428 16676 50484 16678
rect 50508 16676 50564 16678
rect 50588 16676 50644 16678
rect 50348 16624 50374 16676
rect 50374 16624 50404 16676
rect 50428 16624 50438 16676
rect 50438 16624 50484 16676
rect 50508 16624 50554 16676
rect 50554 16624 50564 16676
rect 50588 16624 50618 16676
rect 50618 16624 50644 16676
rect 50348 16622 50404 16624
rect 50428 16622 50484 16624
rect 50508 16622 50564 16624
rect 50588 16622 50644 16624
rect 50348 15344 50404 15346
rect 50428 15344 50484 15346
rect 50508 15344 50564 15346
rect 50588 15344 50644 15346
rect 50348 15292 50374 15344
rect 50374 15292 50404 15344
rect 50428 15292 50438 15344
rect 50438 15292 50484 15344
rect 50508 15292 50554 15344
rect 50554 15292 50564 15344
rect 50588 15292 50618 15344
rect 50618 15292 50644 15344
rect 50348 15290 50404 15292
rect 50428 15290 50484 15292
rect 50508 15290 50564 15292
rect 50588 15290 50644 15292
rect 50348 14012 50404 14014
rect 50428 14012 50484 14014
rect 50508 14012 50564 14014
rect 50588 14012 50644 14014
rect 50348 13960 50374 14012
rect 50374 13960 50404 14012
rect 50428 13960 50438 14012
rect 50438 13960 50484 14012
rect 50508 13960 50554 14012
rect 50554 13960 50564 14012
rect 50588 13960 50618 14012
rect 50618 13960 50644 14012
rect 50348 13958 50404 13960
rect 50428 13958 50484 13960
rect 50508 13958 50564 13960
rect 50588 13958 50644 13960
rect 50348 12680 50404 12682
rect 50428 12680 50484 12682
rect 50508 12680 50564 12682
rect 50588 12680 50644 12682
rect 50348 12628 50374 12680
rect 50374 12628 50404 12680
rect 50428 12628 50438 12680
rect 50438 12628 50484 12680
rect 50508 12628 50554 12680
rect 50554 12628 50564 12680
rect 50588 12628 50618 12680
rect 50618 12628 50644 12680
rect 50348 12626 50404 12628
rect 50428 12626 50484 12628
rect 50508 12626 50564 12628
rect 50588 12626 50644 12628
rect 50348 11348 50404 11350
rect 50428 11348 50484 11350
rect 50508 11348 50564 11350
rect 50588 11348 50644 11350
rect 50348 11296 50374 11348
rect 50374 11296 50404 11348
rect 50428 11296 50438 11348
rect 50438 11296 50484 11348
rect 50508 11296 50554 11348
rect 50554 11296 50564 11348
rect 50588 11296 50618 11348
rect 50618 11296 50644 11348
rect 50348 11294 50404 11296
rect 50428 11294 50484 11296
rect 50508 11294 50564 11296
rect 50588 11294 50644 11296
rect 50348 10016 50404 10018
rect 50428 10016 50484 10018
rect 50508 10016 50564 10018
rect 50588 10016 50644 10018
rect 50348 9964 50374 10016
rect 50374 9964 50404 10016
rect 50428 9964 50438 10016
rect 50438 9964 50484 10016
rect 50508 9964 50554 10016
rect 50554 9964 50564 10016
rect 50588 9964 50618 10016
rect 50618 9964 50644 10016
rect 50348 9962 50404 9964
rect 50428 9962 50484 9964
rect 50508 9962 50564 9964
rect 50588 9962 50644 9964
rect 50348 8684 50404 8686
rect 50428 8684 50484 8686
rect 50508 8684 50564 8686
rect 50588 8684 50644 8686
rect 50348 8632 50374 8684
rect 50374 8632 50404 8684
rect 50428 8632 50438 8684
rect 50438 8632 50484 8684
rect 50508 8632 50554 8684
rect 50554 8632 50564 8684
rect 50588 8632 50618 8684
rect 50618 8632 50644 8684
rect 50348 8630 50404 8632
rect 50428 8630 50484 8632
rect 50508 8630 50564 8632
rect 50588 8630 50644 8632
rect 50348 7352 50404 7354
rect 50428 7352 50484 7354
rect 50508 7352 50564 7354
rect 50588 7352 50644 7354
rect 50348 7300 50374 7352
rect 50374 7300 50404 7352
rect 50428 7300 50438 7352
rect 50438 7300 50484 7352
rect 50508 7300 50554 7352
rect 50554 7300 50564 7352
rect 50588 7300 50618 7352
rect 50618 7300 50644 7352
rect 50348 7298 50404 7300
rect 50428 7298 50484 7300
rect 50508 7298 50564 7300
rect 50588 7298 50644 7300
rect 50348 6020 50404 6022
rect 50428 6020 50484 6022
rect 50508 6020 50564 6022
rect 50588 6020 50644 6022
rect 50348 5968 50374 6020
rect 50374 5968 50404 6020
rect 50428 5968 50438 6020
rect 50438 5968 50484 6020
rect 50508 5968 50554 6020
rect 50554 5968 50564 6020
rect 50588 5968 50618 6020
rect 50618 5968 50644 6020
rect 50348 5966 50404 5968
rect 50428 5966 50484 5968
rect 50508 5966 50564 5968
rect 50588 5966 50644 5968
rect 50348 4688 50404 4690
rect 50428 4688 50484 4690
rect 50508 4688 50564 4690
rect 50588 4688 50644 4690
rect 50348 4636 50374 4688
rect 50374 4636 50404 4688
rect 50428 4636 50438 4688
rect 50438 4636 50484 4688
rect 50508 4636 50554 4688
rect 50554 4636 50564 4688
rect 50588 4636 50618 4688
rect 50618 4636 50644 4688
rect 50348 4634 50404 4636
rect 50428 4634 50484 4636
rect 50508 4634 50564 4636
rect 50588 4634 50644 4636
rect 50348 3356 50404 3358
rect 50428 3356 50484 3358
rect 50508 3356 50564 3358
rect 50588 3356 50644 3358
rect 50348 3304 50374 3356
rect 50374 3304 50404 3356
rect 50428 3304 50438 3356
rect 50438 3304 50484 3356
rect 50508 3304 50554 3356
rect 50554 3304 50564 3356
rect 50588 3304 50618 3356
rect 50618 3304 50644 3356
rect 50348 3302 50404 3304
rect 50428 3302 50484 3304
rect 50508 3302 50564 3304
rect 50588 3302 50644 3304
<< metal3 >>
rect 4256 57308 4576 57309
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 57243 4576 57244
rect 34976 57308 35296 57309
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 57243 35296 57244
rect 19616 56642 19936 56643
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 56577 19936 56578
rect 50336 56642 50656 56643
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 56577 50656 56578
rect 4256 55976 4576 55977
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 55911 4576 55912
rect 34976 55976 35296 55977
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 55911 35296 55912
rect 19616 55310 19936 55311
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 55245 19936 55246
rect 50336 55310 50656 55311
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 55245 50656 55246
rect 4256 54644 4576 54645
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 54579 4576 54580
rect 34976 54644 35296 54645
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 54579 35296 54580
rect 19616 53978 19936 53979
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 53913 19936 53914
rect 50336 53978 50656 53979
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 53913 50656 53914
rect 4256 53312 4576 53313
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 53247 4576 53248
rect 34976 53312 35296 53313
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 53247 35296 53248
rect 19616 52646 19936 52647
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 52581 19936 52582
rect 50336 52646 50656 52647
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 52581 50656 52582
rect 4256 51980 4576 51981
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 51915 4576 51916
rect 34976 51980 35296 51981
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 51915 35296 51916
rect 19616 51314 19936 51315
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 51249 19936 51250
rect 50336 51314 50656 51315
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 51249 50656 51250
rect 4256 50648 4576 50649
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 50583 4576 50584
rect 34976 50648 35296 50649
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 50583 35296 50584
rect 19616 49982 19936 49983
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 49917 19936 49918
rect 50336 49982 50656 49983
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 49917 50656 49918
rect 4256 49316 4576 49317
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 49251 4576 49252
rect 34976 49316 35296 49317
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 49251 35296 49252
rect 19616 48650 19936 48651
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 48585 19936 48586
rect 50336 48650 50656 48651
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 48585 50656 48586
rect 4256 47984 4576 47985
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 47919 4576 47920
rect 34976 47984 35296 47985
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 47919 35296 47920
rect 19616 47318 19936 47319
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 47253 19936 47254
rect 50336 47318 50656 47319
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 47253 50656 47254
rect 4256 46652 4576 46653
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 46587 4576 46588
rect 34976 46652 35296 46653
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 46587 35296 46588
rect 19616 45986 19936 45987
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 45921 19936 45922
rect 50336 45986 50656 45987
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 45921 50656 45922
rect 4256 45320 4576 45321
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 45255 4576 45256
rect 34976 45320 35296 45321
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 45255 35296 45256
rect 19616 44654 19936 44655
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 44589 19936 44590
rect 50336 44654 50656 44655
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 44589 50656 44590
rect 4256 43988 4576 43989
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 43923 4576 43924
rect 34976 43988 35296 43989
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 43923 35296 43924
rect 19616 43322 19936 43323
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 43257 19936 43258
rect 50336 43322 50656 43323
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 43257 50656 43258
rect 4256 42656 4576 42657
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 42591 4576 42592
rect 34976 42656 35296 42657
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 42591 35296 42592
rect 19616 41990 19936 41991
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 41925 19936 41926
rect 50336 41990 50656 41991
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 41925 50656 41926
rect 4256 41324 4576 41325
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 41259 4576 41260
rect 34976 41324 35296 41325
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 41259 35296 41260
rect 19616 40658 19936 40659
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 40593 19936 40594
rect 50336 40658 50656 40659
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 40593 50656 40594
rect 4256 39992 4576 39993
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 39927 4576 39928
rect 34976 39992 35296 39993
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 39927 35296 39928
rect 19616 39326 19936 39327
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 39261 19936 39262
rect 50336 39326 50656 39327
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 39261 50656 39262
rect 4256 38660 4576 38661
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 38595 4576 38596
rect 34976 38660 35296 38661
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 38595 35296 38596
rect 19616 37994 19936 37995
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 37929 19936 37930
rect 50336 37994 50656 37995
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 37929 50656 37930
rect 4256 37328 4576 37329
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 37263 4576 37264
rect 34976 37328 35296 37329
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 37263 35296 37264
rect 19616 36662 19936 36663
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 36597 19936 36598
rect 50336 36662 50656 36663
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 36597 50656 36598
rect 4256 35996 4576 35997
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 35931 4576 35932
rect 34976 35996 35296 35997
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 35931 35296 35932
rect 19616 35330 19936 35331
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 35265 19936 35266
rect 50336 35330 50656 35331
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 35265 50656 35266
rect 4256 34664 4576 34665
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 34599 4576 34600
rect 34976 34664 35296 34665
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 34599 35296 34600
rect 19616 33998 19936 33999
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 33933 19936 33934
rect 50336 33998 50656 33999
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 33933 50656 33934
rect 4256 33332 4576 33333
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 33267 4576 33268
rect 34976 33332 35296 33333
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 33267 35296 33268
rect 19616 32666 19936 32667
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 32601 19936 32602
rect 50336 32666 50656 32667
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 32601 50656 32602
rect 4256 32000 4576 32001
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 31935 4576 31936
rect 34976 32000 35296 32001
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 31935 35296 31936
rect 19616 31334 19936 31335
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 31269 19936 31270
rect 50336 31334 50656 31335
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 31269 50656 31270
rect 4256 30668 4576 30669
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 30603 4576 30604
rect 34976 30668 35296 30669
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 30603 35296 30604
rect 19616 30002 19936 30003
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 29937 19936 29938
rect 50336 30002 50656 30003
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 29937 50656 29938
rect 4256 29336 4576 29337
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 29271 4576 29272
rect 34976 29336 35296 29337
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 29271 35296 29272
rect 19616 28670 19936 28671
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 28605 19936 28606
rect 50336 28670 50656 28671
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 28605 50656 28606
rect 4256 28004 4576 28005
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 27939 4576 27940
rect 34976 28004 35296 28005
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 27939 35296 27940
rect 19616 27338 19936 27339
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 27273 19936 27274
rect 50336 27338 50656 27339
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 27273 50656 27274
rect 4256 26672 4576 26673
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 26607 4576 26608
rect 34976 26672 35296 26673
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 26607 35296 26608
rect 19616 26006 19936 26007
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 25941 19936 25942
rect 50336 26006 50656 26007
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 25941 50656 25942
rect 4256 25340 4576 25341
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 25275 4576 25276
rect 34976 25340 35296 25341
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 25275 35296 25276
rect 19616 24674 19936 24675
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 24609 19936 24610
rect 50336 24674 50656 24675
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 24609 50656 24610
rect 4256 24008 4576 24009
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 23943 4576 23944
rect 34976 24008 35296 24009
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 23943 35296 23944
rect 19616 23342 19936 23343
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 23277 19936 23278
rect 50336 23342 50656 23343
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 23277 50656 23278
rect 4256 22676 4576 22677
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 22611 4576 22612
rect 34976 22676 35296 22677
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 22611 35296 22612
rect 19616 22010 19936 22011
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 21945 19936 21946
rect 50336 22010 50656 22011
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 21945 50656 21946
rect 4256 21344 4576 21345
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 21279 4576 21280
rect 34976 21344 35296 21345
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 21279 35296 21280
rect 19616 20678 19936 20679
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 20613 19936 20614
rect 50336 20678 50656 20679
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 20613 50656 20614
rect 4256 20012 4576 20013
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 19947 4576 19948
rect 34976 20012 35296 20013
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 19947 35296 19948
rect 19616 19346 19936 19347
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 19281 19936 19282
rect 50336 19346 50656 19347
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 19281 50656 19282
rect 4256 18680 4576 18681
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 18615 4576 18616
rect 34976 18680 35296 18681
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 18615 35296 18616
rect 19616 18014 19936 18015
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 17949 19936 17950
rect 50336 18014 50656 18015
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 17949 50656 17950
rect 4256 17348 4576 17349
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 17283 4576 17284
rect 34976 17348 35296 17349
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 17283 35296 17284
rect 19616 16682 19936 16683
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 16617 19936 16618
rect 50336 16682 50656 16683
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 16617 50656 16618
rect 4256 16016 4576 16017
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 15951 4576 15952
rect 34976 16016 35296 16017
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 15951 35296 15952
rect 19616 15350 19936 15351
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 15285 19936 15286
rect 50336 15350 50656 15351
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 15285 50656 15286
rect 4256 14684 4576 14685
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 14619 4576 14620
rect 34976 14684 35296 14685
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 14619 35296 14620
rect 19616 14018 19936 14019
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 13953 19936 13954
rect 50336 14018 50656 14019
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 13953 50656 13954
rect 4256 13352 4576 13353
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 13287 4576 13288
rect 34976 13352 35296 13353
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 13287 35296 13288
rect 19616 12686 19936 12687
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 12621 19936 12622
rect 50336 12686 50656 12687
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 12621 50656 12622
rect 4256 12020 4576 12021
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 11955 4576 11956
rect 34976 12020 35296 12021
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 11955 35296 11956
rect 19616 11354 19936 11355
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 11289 19936 11290
rect 50336 11354 50656 11355
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 11289 50656 11290
rect 4256 10688 4576 10689
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 10623 4576 10624
rect 34976 10688 35296 10689
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 10623 35296 10624
rect 19616 10022 19936 10023
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 9957 19936 9958
rect 50336 10022 50656 10023
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 9957 50656 9958
rect 4256 9356 4576 9357
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 9291 4576 9292
rect 34976 9356 35296 9357
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 9291 35296 9292
rect 19616 8690 19936 8691
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 8625 19936 8626
rect 50336 8690 50656 8691
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 8625 50656 8626
rect 4256 8024 4576 8025
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 7959 4576 7960
rect 34976 8024 35296 8025
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 7959 35296 7960
rect 19616 7358 19936 7359
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 7293 19936 7294
rect 50336 7358 50656 7359
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 7293 50656 7294
rect 4256 6692 4576 6693
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 6627 4576 6628
rect 34976 6692 35296 6693
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 6627 35296 6628
rect 19616 6026 19936 6027
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 5961 19936 5962
rect 50336 6026 50656 6027
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 5961 50656 5962
rect 4256 5360 4576 5361
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 5295 4576 5296
rect 34976 5360 35296 5361
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 5295 35296 5296
rect 19616 4694 19936 4695
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 4629 19936 4630
rect 50336 4694 50656 4695
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 4629 50656 4630
rect 4256 4028 4576 4029
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 3963 4576 3964
rect 34976 4028 35296 4029
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 3963 35296 3964
rect 19616 3362 19936 3363
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 19616 3297 19936 3298
rect 50336 3362 50656 3363
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 50336 3297 50656 3298
rect 41775 3064 41841 3067
rect 44367 3064 44433 3067
rect 41775 3062 44433 3064
rect 41775 3006 41780 3062
rect 41836 3006 44372 3062
rect 44428 3006 44433 3062
rect 41775 3004 44433 3006
rect 41775 3001 41841 3004
rect 44367 3001 44433 3004
rect 4256 2696 4576 2697
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4256 2631 4576 2632
rect 34976 2696 35296 2697
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 34976 2631 35296 2632
<< via3 >>
rect 4264 57304 4328 57308
rect 4264 57248 4268 57304
rect 4268 57248 4324 57304
rect 4324 57248 4328 57304
rect 4264 57244 4328 57248
rect 4344 57304 4408 57308
rect 4344 57248 4348 57304
rect 4348 57248 4404 57304
rect 4404 57248 4408 57304
rect 4344 57244 4408 57248
rect 4424 57304 4488 57308
rect 4424 57248 4428 57304
rect 4428 57248 4484 57304
rect 4484 57248 4488 57304
rect 4424 57244 4488 57248
rect 4504 57304 4568 57308
rect 4504 57248 4508 57304
rect 4508 57248 4564 57304
rect 4564 57248 4568 57304
rect 4504 57244 4568 57248
rect 34984 57304 35048 57308
rect 34984 57248 34988 57304
rect 34988 57248 35044 57304
rect 35044 57248 35048 57304
rect 34984 57244 35048 57248
rect 35064 57304 35128 57308
rect 35064 57248 35068 57304
rect 35068 57248 35124 57304
rect 35124 57248 35128 57304
rect 35064 57244 35128 57248
rect 35144 57304 35208 57308
rect 35144 57248 35148 57304
rect 35148 57248 35204 57304
rect 35204 57248 35208 57304
rect 35144 57244 35208 57248
rect 35224 57304 35288 57308
rect 35224 57248 35228 57304
rect 35228 57248 35284 57304
rect 35284 57248 35288 57304
rect 35224 57244 35288 57248
rect 19624 56638 19688 56642
rect 19624 56582 19628 56638
rect 19628 56582 19684 56638
rect 19684 56582 19688 56638
rect 19624 56578 19688 56582
rect 19704 56638 19768 56642
rect 19704 56582 19708 56638
rect 19708 56582 19764 56638
rect 19764 56582 19768 56638
rect 19704 56578 19768 56582
rect 19784 56638 19848 56642
rect 19784 56582 19788 56638
rect 19788 56582 19844 56638
rect 19844 56582 19848 56638
rect 19784 56578 19848 56582
rect 19864 56638 19928 56642
rect 19864 56582 19868 56638
rect 19868 56582 19924 56638
rect 19924 56582 19928 56638
rect 19864 56578 19928 56582
rect 50344 56638 50408 56642
rect 50344 56582 50348 56638
rect 50348 56582 50404 56638
rect 50404 56582 50408 56638
rect 50344 56578 50408 56582
rect 50424 56638 50488 56642
rect 50424 56582 50428 56638
rect 50428 56582 50484 56638
rect 50484 56582 50488 56638
rect 50424 56578 50488 56582
rect 50504 56638 50568 56642
rect 50504 56582 50508 56638
rect 50508 56582 50564 56638
rect 50564 56582 50568 56638
rect 50504 56578 50568 56582
rect 50584 56638 50648 56642
rect 50584 56582 50588 56638
rect 50588 56582 50644 56638
rect 50644 56582 50648 56638
rect 50584 56578 50648 56582
rect 4264 55972 4328 55976
rect 4264 55916 4268 55972
rect 4268 55916 4324 55972
rect 4324 55916 4328 55972
rect 4264 55912 4328 55916
rect 4344 55972 4408 55976
rect 4344 55916 4348 55972
rect 4348 55916 4404 55972
rect 4404 55916 4408 55972
rect 4344 55912 4408 55916
rect 4424 55972 4488 55976
rect 4424 55916 4428 55972
rect 4428 55916 4484 55972
rect 4484 55916 4488 55972
rect 4424 55912 4488 55916
rect 4504 55972 4568 55976
rect 4504 55916 4508 55972
rect 4508 55916 4564 55972
rect 4564 55916 4568 55972
rect 4504 55912 4568 55916
rect 34984 55972 35048 55976
rect 34984 55916 34988 55972
rect 34988 55916 35044 55972
rect 35044 55916 35048 55972
rect 34984 55912 35048 55916
rect 35064 55972 35128 55976
rect 35064 55916 35068 55972
rect 35068 55916 35124 55972
rect 35124 55916 35128 55972
rect 35064 55912 35128 55916
rect 35144 55972 35208 55976
rect 35144 55916 35148 55972
rect 35148 55916 35204 55972
rect 35204 55916 35208 55972
rect 35144 55912 35208 55916
rect 35224 55972 35288 55976
rect 35224 55916 35228 55972
rect 35228 55916 35284 55972
rect 35284 55916 35288 55972
rect 35224 55912 35288 55916
rect 19624 55306 19688 55310
rect 19624 55250 19628 55306
rect 19628 55250 19684 55306
rect 19684 55250 19688 55306
rect 19624 55246 19688 55250
rect 19704 55306 19768 55310
rect 19704 55250 19708 55306
rect 19708 55250 19764 55306
rect 19764 55250 19768 55306
rect 19704 55246 19768 55250
rect 19784 55306 19848 55310
rect 19784 55250 19788 55306
rect 19788 55250 19844 55306
rect 19844 55250 19848 55306
rect 19784 55246 19848 55250
rect 19864 55306 19928 55310
rect 19864 55250 19868 55306
rect 19868 55250 19924 55306
rect 19924 55250 19928 55306
rect 19864 55246 19928 55250
rect 50344 55306 50408 55310
rect 50344 55250 50348 55306
rect 50348 55250 50404 55306
rect 50404 55250 50408 55306
rect 50344 55246 50408 55250
rect 50424 55306 50488 55310
rect 50424 55250 50428 55306
rect 50428 55250 50484 55306
rect 50484 55250 50488 55306
rect 50424 55246 50488 55250
rect 50504 55306 50568 55310
rect 50504 55250 50508 55306
rect 50508 55250 50564 55306
rect 50564 55250 50568 55306
rect 50504 55246 50568 55250
rect 50584 55306 50648 55310
rect 50584 55250 50588 55306
rect 50588 55250 50644 55306
rect 50644 55250 50648 55306
rect 50584 55246 50648 55250
rect 4264 54640 4328 54644
rect 4264 54584 4268 54640
rect 4268 54584 4324 54640
rect 4324 54584 4328 54640
rect 4264 54580 4328 54584
rect 4344 54640 4408 54644
rect 4344 54584 4348 54640
rect 4348 54584 4404 54640
rect 4404 54584 4408 54640
rect 4344 54580 4408 54584
rect 4424 54640 4488 54644
rect 4424 54584 4428 54640
rect 4428 54584 4484 54640
rect 4484 54584 4488 54640
rect 4424 54580 4488 54584
rect 4504 54640 4568 54644
rect 4504 54584 4508 54640
rect 4508 54584 4564 54640
rect 4564 54584 4568 54640
rect 4504 54580 4568 54584
rect 34984 54640 35048 54644
rect 34984 54584 34988 54640
rect 34988 54584 35044 54640
rect 35044 54584 35048 54640
rect 34984 54580 35048 54584
rect 35064 54640 35128 54644
rect 35064 54584 35068 54640
rect 35068 54584 35124 54640
rect 35124 54584 35128 54640
rect 35064 54580 35128 54584
rect 35144 54640 35208 54644
rect 35144 54584 35148 54640
rect 35148 54584 35204 54640
rect 35204 54584 35208 54640
rect 35144 54580 35208 54584
rect 35224 54640 35288 54644
rect 35224 54584 35228 54640
rect 35228 54584 35284 54640
rect 35284 54584 35288 54640
rect 35224 54580 35288 54584
rect 19624 53974 19688 53978
rect 19624 53918 19628 53974
rect 19628 53918 19684 53974
rect 19684 53918 19688 53974
rect 19624 53914 19688 53918
rect 19704 53974 19768 53978
rect 19704 53918 19708 53974
rect 19708 53918 19764 53974
rect 19764 53918 19768 53974
rect 19704 53914 19768 53918
rect 19784 53974 19848 53978
rect 19784 53918 19788 53974
rect 19788 53918 19844 53974
rect 19844 53918 19848 53974
rect 19784 53914 19848 53918
rect 19864 53974 19928 53978
rect 19864 53918 19868 53974
rect 19868 53918 19924 53974
rect 19924 53918 19928 53974
rect 19864 53914 19928 53918
rect 50344 53974 50408 53978
rect 50344 53918 50348 53974
rect 50348 53918 50404 53974
rect 50404 53918 50408 53974
rect 50344 53914 50408 53918
rect 50424 53974 50488 53978
rect 50424 53918 50428 53974
rect 50428 53918 50484 53974
rect 50484 53918 50488 53974
rect 50424 53914 50488 53918
rect 50504 53974 50568 53978
rect 50504 53918 50508 53974
rect 50508 53918 50564 53974
rect 50564 53918 50568 53974
rect 50504 53914 50568 53918
rect 50584 53974 50648 53978
rect 50584 53918 50588 53974
rect 50588 53918 50644 53974
rect 50644 53918 50648 53974
rect 50584 53914 50648 53918
rect 4264 53308 4328 53312
rect 4264 53252 4268 53308
rect 4268 53252 4324 53308
rect 4324 53252 4328 53308
rect 4264 53248 4328 53252
rect 4344 53308 4408 53312
rect 4344 53252 4348 53308
rect 4348 53252 4404 53308
rect 4404 53252 4408 53308
rect 4344 53248 4408 53252
rect 4424 53308 4488 53312
rect 4424 53252 4428 53308
rect 4428 53252 4484 53308
rect 4484 53252 4488 53308
rect 4424 53248 4488 53252
rect 4504 53308 4568 53312
rect 4504 53252 4508 53308
rect 4508 53252 4564 53308
rect 4564 53252 4568 53308
rect 4504 53248 4568 53252
rect 34984 53308 35048 53312
rect 34984 53252 34988 53308
rect 34988 53252 35044 53308
rect 35044 53252 35048 53308
rect 34984 53248 35048 53252
rect 35064 53308 35128 53312
rect 35064 53252 35068 53308
rect 35068 53252 35124 53308
rect 35124 53252 35128 53308
rect 35064 53248 35128 53252
rect 35144 53308 35208 53312
rect 35144 53252 35148 53308
rect 35148 53252 35204 53308
rect 35204 53252 35208 53308
rect 35144 53248 35208 53252
rect 35224 53308 35288 53312
rect 35224 53252 35228 53308
rect 35228 53252 35284 53308
rect 35284 53252 35288 53308
rect 35224 53248 35288 53252
rect 19624 52642 19688 52646
rect 19624 52586 19628 52642
rect 19628 52586 19684 52642
rect 19684 52586 19688 52642
rect 19624 52582 19688 52586
rect 19704 52642 19768 52646
rect 19704 52586 19708 52642
rect 19708 52586 19764 52642
rect 19764 52586 19768 52642
rect 19704 52582 19768 52586
rect 19784 52642 19848 52646
rect 19784 52586 19788 52642
rect 19788 52586 19844 52642
rect 19844 52586 19848 52642
rect 19784 52582 19848 52586
rect 19864 52642 19928 52646
rect 19864 52586 19868 52642
rect 19868 52586 19924 52642
rect 19924 52586 19928 52642
rect 19864 52582 19928 52586
rect 50344 52642 50408 52646
rect 50344 52586 50348 52642
rect 50348 52586 50404 52642
rect 50404 52586 50408 52642
rect 50344 52582 50408 52586
rect 50424 52642 50488 52646
rect 50424 52586 50428 52642
rect 50428 52586 50484 52642
rect 50484 52586 50488 52642
rect 50424 52582 50488 52586
rect 50504 52642 50568 52646
rect 50504 52586 50508 52642
rect 50508 52586 50564 52642
rect 50564 52586 50568 52642
rect 50504 52582 50568 52586
rect 50584 52642 50648 52646
rect 50584 52586 50588 52642
rect 50588 52586 50644 52642
rect 50644 52586 50648 52642
rect 50584 52582 50648 52586
rect 4264 51976 4328 51980
rect 4264 51920 4268 51976
rect 4268 51920 4324 51976
rect 4324 51920 4328 51976
rect 4264 51916 4328 51920
rect 4344 51976 4408 51980
rect 4344 51920 4348 51976
rect 4348 51920 4404 51976
rect 4404 51920 4408 51976
rect 4344 51916 4408 51920
rect 4424 51976 4488 51980
rect 4424 51920 4428 51976
rect 4428 51920 4484 51976
rect 4484 51920 4488 51976
rect 4424 51916 4488 51920
rect 4504 51976 4568 51980
rect 4504 51920 4508 51976
rect 4508 51920 4564 51976
rect 4564 51920 4568 51976
rect 4504 51916 4568 51920
rect 34984 51976 35048 51980
rect 34984 51920 34988 51976
rect 34988 51920 35044 51976
rect 35044 51920 35048 51976
rect 34984 51916 35048 51920
rect 35064 51976 35128 51980
rect 35064 51920 35068 51976
rect 35068 51920 35124 51976
rect 35124 51920 35128 51976
rect 35064 51916 35128 51920
rect 35144 51976 35208 51980
rect 35144 51920 35148 51976
rect 35148 51920 35204 51976
rect 35204 51920 35208 51976
rect 35144 51916 35208 51920
rect 35224 51976 35288 51980
rect 35224 51920 35228 51976
rect 35228 51920 35284 51976
rect 35284 51920 35288 51976
rect 35224 51916 35288 51920
rect 19624 51310 19688 51314
rect 19624 51254 19628 51310
rect 19628 51254 19684 51310
rect 19684 51254 19688 51310
rect 19624 51250 19688 51254
rect 19704 51310 19768 51314
rect 19704 51254 19708 51310
rect 19708 51254 19764 51310
rect 19764 51254 19768 51310
rect 19704 51250 19768 51254
rect 19784 51310 19848 51314
rect 19784 51254 19788 51310
rect 19788 51254 19844 51310
rect 19844 51254 19848 51310
rect 19784 51250 19848 51254
rect 19864 51310 19928 51314
rect 19864 51254 19868 51310
rect 19868 51254 19924 51310
rect 19924 51254 19928 51310
rect 19864 51250 19928 51254
rect 50344 51310 50408 51314
rect 50344 51254 50348 51310
rect 50348 51254 50404 51310
rect 50404 51254 50408 51310
rect 50344 51250 50408 51254
rect 50424 51310 50488 51314
rect 50424 51254 50428 51310
rect 50428 51254 50484 51310
rect 50484 51254 50488 51310
rect 50424 51250 50488 51254
rect 50504 51310 50568 51314
rect 50504 51254 50508 51310
rect 50508 51254 50564 51310
rect 50564 51254 50568 51310
rect 50504 51250 50568 51254
rect 50584 51310 50648 51314
rect 50584 51254 50588 51310
rect 50588 51254 50644 51310
rect 50644 51254 50648 51310
rect 50584 51250 50648 51254
rect 4264 50644 4328 50648
rect 4264 50588 4268 50644
rect 4268 50588 4324 50644
rect 4324 50588 4328 50644
rect 4264 50584 4328 50588
rect 4344 50644 4408 50648
rect 4344 50588 4348 50644
rect 4348 50588 4404 50644
rect 4404 50588 4408 50644
rect 4344 50584 4408 50588
rect 4424 50644 4488 50648
rect 4424 50588 4428 50644
rect 4428 50588 4484 50644
rect 4484 50588 4488 50644
rect 4424 50584 4488 50588
rect 4504 50644 4568 50648
rect 4504 50588 4508 50644
rect 4508 50588 4564 50644
rect 4564 50588 4568 50644
rect 4504 50584 4568 50588
rect 34984 50644 35048 50648
rect 34984 50588 34988 50644
rect 34988 50588 35044 50644
rect 35044 50588 35048 50644
rect 34984 50584 35048 50588
rect 35064 50644 35128 50648
rect 35064 50588 35068 50644
rect 35068 50588 35124 50644
rect 35124 50588 35128 50644
rect 35064 50584 35128 50588
rect 35144 50644 35208 50648
rect 35144 50588 35148 50644
rect 35148 50588 35204 50644
rect 35204 50588 35208 50644
rect 35144 50584 35208 50588
rect 35224 50644 35288 50648
rect 35224 50588 35228 50644
rect 35228 50588 35284 50644
rect 35284 50588 35288 50644
rect 35224 50584 35288 50588
rect 19624 49978 19688 49982
rect 19624 49922 19628 49978
rect 19628 49922 19684 49978
rect 19684 49922 19688 49978
rect 19624 49918 19688 49922
rect 19704 49978 19768 49982
rect 19704 49922 19708 49978
rect 19708 49922 19764 49978
rect 19764 49922 19768 49978
rect 19704 49918 19768 49922
rect 19784 49978 19848 49982
rect 19784 49922 19788 49978
rect 19788 49922 19844 49978
rect 19844 49922 19848 49978
rect 19784 49918 19848 49922
rect 19864 49978 19928 49982
rect 19864 49922 19868 49978
rect 19868 49922 19924 49978
rect 19924 49922 19928 49978
rect 19864 49918 19928 49922
rect 50344 49978 50408 49982
rect 50344 49922 50348 49978
rect 50348 49922 50404 49978
rect 50404 49922 50408 49978
rect 50344 49918 50408 49922
rect 50424 49978 50488 49982
rect 50424 49922 50428 49978
rect 50428 49922 50484 49978
rect 50484 49922 50488 49978
rect 50424 49918 50488 49922
rect 50504 49978 50568 49982
rect 50504 49922 50508 49978
rect 50508 49922 50564 49978
rect 50564 49922 50568 49978
rect 50504 49918 50568 49922
rect 50584 49978 50648 49982
rect 50584 49922 50588 49978
rect 50588 49922 50644 49978
rect 50644 49922 50648 49978
rect 50584 49918 50648 49922
rect 4264 49312 4328 49316
rect 4264 49256 4268 49312
rect 4268 49256 4324 49312
rect 4324 49256 4328 49312
rect 4264 49252 4328 49256
rect 4344 49312 4408 49316
rect 4344 49256 4348 49312
rect 4348 49256 4404 49312
rect 4404 49256 4408 49312
rect 4344 49252 4408 49256
rect 4424 49312 4488 49316
rect 4424 49256 4428 49312
rect 4428 49256 4484 49312
rect 4484 49256 4488 49312
rect 4424 49252 4488 49256
rect 4504 49312 4568 49316
rect 4504 49256 4508 49312
rect 4508 49256 4564 49312
rect 4564 49256 4568 49312
rect 4504 49252 4568 49256
rect 34984 49312 35048 49316
rect 34984 49256 34988 49312
rect 34988 49256 35044 49312
rect 35044 49256 35048 49312
rect 34984 49252 35048 49256
rect 35064 49312 35128 49316
rect 35064 49256 35068 49312
rect 35068 49256 35124 49312
rect 35124 49256 35128 49312
rect 35064 49252 35128 49256
rect 35144 49312 35208 49316
rect 35144 49256 35148 49312
rect 35148 49256 35204 49312
rect 35204 49256 35208 49312
rect 35144 49252 35208 49256
rect 35224 49312 35288 49316
rect 35224 49256 35228 49312
rect 35228 49256 35284 49312
rect 35284 49256 35288 49312
rect 35224 49252 35288 49256
rect 19624 48646 19688 48650
rect 19624 48590 19628 48646
rect 19628 48590 19684 48646
rect 19684 48590 19688 48646
rect 19624 48586 19688 48590
rect 19704 48646 19768 48650
rect 19704 48590 19708 48646
rect 19708 48590 19764 48646
rect 19764 48590 19768 48646
rect 19704 48586 19768 48590
rect 19784 48646 19848 48650
rect 19784 48590 19788 48646
rect 19788 48590 19844 48646
rect 19844 48590 19848 48646
rect 19784 48586 19848 48590
rect 19864 48646 19928 48650
rect 19864 48590 19868 48646
rect 19868 48590 19924 48646
rect 19924 48590 19928 48646
rect 19864 48586 19928 48590
rect 50344 48646 50408 48650
rect 50344 48590 50348 48646
rect 50348 48590 50404 48646
rect 50404 48590 50408 48646
rect 50344 48586 50408 48590
rect 50424 48646 50488 48650
rect 50424 48590 50428 48646
rect 50428 48590 50484 48646
rect 50484 48590 50488 48646
rect 50424 48586 50488 48590
rect 50504 48646 50568 48650
rect 50504 48590 50508 48646
rect 50508 48590 50564 48646
rect 50564 48590 50568 48646
rect 50504 48586 50568 48590
rect 50584 48646 50648 48650
rect 50584 48590 50588 48646
rect 50588 48590 50644 48646
rect 50644 48590 50648 48646
rect 50584 48586 50648 48590
rect 4264 47980 4328 47984
rect 4264 47924 4268 47980
rect 4268 47924 4324 47980
rect 4324 47924 4328 47980
rect 4264 47920 4328 47924
rect 4344 47980 4408 47984
rect 4344 47924 4348 47980
rect 4348 47924 4404 47980
rect 4404 47924 4408 47980
rect 4344 47920 4408 47924
rect 4424 47980 4488 47984
rect 4424 47924 4428 47980
rect 4428 47924 4484 47980
rect 4484 47924 4488 47980
rect 4424 47920 4488 47924
rect 4504 47980 4568 47984
rect 4504 47924 4508 47980
rect 4508 47924 4564 47980
rect 4564 47924 4568 47980
rect 4504 47920 4568 47924
rect 34984 47980 35048 47984
rect 34984 47924 34988 47980
rect 34988 47924 35044 47980
rect 35044 47924 35048 47980
rect 34984 47920 35048 47924
rect 35064 47980 35128 47984
rect 35064 47924 35068 47980
rect 35068 47924 35124 47980
rect 35124 47924 35128 47980
rect 35064 47920 35128 47924
rect 35144 47980 35208 47984
rect 35144 47924 35148 47980
rect 35148 47924 35204 47980
rect 35204 47924 35208 47980
rect 35144 47920 35208 47924
rect 35224 47980 35288 47984
rect 35224 47924 35228 47980
rect 35228 47924 35284 47980
rect 35284 47924 35288 47980
rect 35224 47920 35288 47924
rect 19624 47314 19688 47318
rect 19624 47258 19628 47314
rect 19628 47258 19684 47314
rect 19684 47258 19688 47314
rect 19624 47254 19688 47258
rect 19704 47314 19768 47318
rect 19704 47258 19708 47314
rect 19708 47258 19764 47314
rect 19764 47258 19768 47314
rect 19704 47254 19768 47258
rect 19784 47314 19848 47318
rect 19784 47258 19788 47314
rect 19788 47258 19844 47314
rect 19844 47258 19848 47314
rect 19784 47254 19848 47258
rect 19864 47314 19928 47318
rect 19864 47258 19868 47314
rect 19868 47258 19924 47314
rect 19924 47258 19928 47314
rect 19864 47254 19928 47258
rect 50344 47314 50408 47318
rect 50344 47258 50348 47314
rect 50348 47258 50404 47314
rect 50404 47258 50408 47314
rect 50344 47254 50408 47258
rect 50424 47314 50488 47318
rect 50424 47258 50428 47314
rect 50428 47258 50484 47314
rect 50484 47258 50488 47314
rect 50424 47254 50488 47258
rect 50504 47314 50568 47318
rect 50504 47258 50508 47314
rect 50508 47258 50564 47314
rect 50564 47258 50568 47314
rect 50504 47254 50568 47258
rect 50584 47314 50648 47318
rect 50584 47258 50588 47314
rect 50588 47258 50644 47314
rect 50644 47258 50648 47314
rect 50584 47254 50648 47258
rect 4264 46648 4328 46652
rect 4264 46592 4268 46648
rect 4268 46592 4324 46648
rect 4324 46592 4328 46648
rect 4264 46588 4328 46592
rect 4344 46648 4408 46652
rect 4344 46592 4348 46648
rect 4348 46592 4404 46648
rect 4404 46592 4408 46648
rect 4344 46588 4408 46592
rect 4424 46648 4488 46652
rect 4424 46592 4428 46648
rect 4428 46592 4484 46648
rect 4484 46592 4488 46648
rect 4424 46588 4488 46592
rect 4504 46648 4568 46652
rect 4504 46592 4508 46648
rect 4508 46592 4564 46648
rect 4564 46592 4568 46648
rect 4504 46588 4568 46592
rect 34984 46648 35048 46652
rect 34984 46592 34988 46648
rect 34988 46592 35044 46648
rect 35044 46592 35048 46648
rect 34984 46588 35048 46592
rect 35064 46648 35128 46652
rect 35064 46592 35068 46648
rect 35068 46592 35124 46648
rect 35124 46592 35128 46648
rect 35064 46588 35128 46592
rect 35144 46648 35208 46652
rect 35144 46592 35148 46648
rect 35148 46592 35204 46648
rect 35204 46592 35208 46648
rect 35144 46588 35208 46592
rect 35224 46648 35288 46652
rect 35224 46592 35228 46648
rect 35228 46592 35284 46648
rect 35284 46592 35288 46648
rect 35224 46588 35288 46592
rect 19624 45982 19688 45986
rect 19624 45926 19628 45982
rect 19628 45926 19684 45982
rect 19684 45926 19688 45982
rect 19624 45922 19688 45926
rect 19704 45982 19768 45986
rect 19704 45926 19708 45982
rect 19708 45926 19764 45982
rect 19764 45926 19768 45982
rect 19704 45922 19768 45926
rect 19784 45982 19848 45986
rect 19784 45926 19788 45982
rect 19788 45926 19844 45982
rect 19844 45926 19848 45982
rect 19784 45922 19848 45926
rect 19864 45982 19928 45986
rect 19864 45926 19868 45982
rect 19868 45926 19924 45982
rect 19924 45926 19928 45982
rect 19864 45922 19928 45926
rect 50344 45982 50408 45986
rect 50344 45926 50348 45982
rect 50348 45926 50404 45982
rect 50404 45926 50408 45982
rect 50344 45922 50408 45926
rect 50424 45982 50488 45986
rect 50424 45926 50428 45982
rect 50428 45926 50484 45982
rect 50484 45926 50488 45982
rect 50424 45922 50488 45926
rect 50504 45982 50568 45986
rect 50504 45926 50508 45982
rect 50508 45926 50564 45982
rect 50564 45926 50568 45982
rect 50504 45922 50568 45926
rect 50584 45982 50648 45986
rect 50584 45926 50588 45982
rect 50588 45926 50644 45982
rect 50644 45926 50648 45982
rect 50584 45922 50648 45926
rect 4264 45316 4328 45320
rect 4264 45260 4268 45316
rect 4268 45260 4324 45316
rect 4324 45260 4328 45316
rect 4264 45256 4328 45260
rect 4344 45316 4408 45320
rect 4344 45260 4348 45316
rect 4348 45260 4404 45316
rect 4404 45260 4408 45316
rect 4344 45256 4408 45260
rect 4424 45316 4488 45320
rect 4424 45260 4428 45316
rect 4428 45260 4484 45316
rect 4484 45260 4488 45316
rect 4424 45256 4488 45260
rect 4504 45316 4568 45320
rect 4504 45260 4508 45316
rect 4508 45260 4564 45316
rect 4564 45260 4568 45316
rect 4504 45256 4568 45260
rect 34984 45316 35048 45320
rect 34984 45260 34988 45316
rect 34988 45260 35044 45316
rect 35044 45260 35048 45316
rect 34984 45256 35048 45260
rect 35064 45316 35128 45320
rect 35064 45260 35068 45316
rect 35068 45260 35124 45316
rect 35124 45260 35128 45316
rect 35064 45256 35128 45260
rect 35144 45316 35208 45320
rect 35144 45260 35148 45316
rect 35148 45260 35204 45316
rect 35204 45260 35208 45316
rect 35144 45256 35208 45260
rect 35224 45316 35288 45320
rect 35224 45260 35228 45316
rect 35228 45260 35284 45316
rect 35284 45260 35288 45316
rect 35224 45256 35288 45260
rect 19624 44650 19688 44654
rect 19624 44594 19628 44650
rect 19628 44594 19684 44650
rect 19684 44594 19688 44650
rect 19624 44590 19688 44594
rect 19704 44650 19768 44654
rect 19704 44594 19708 44650
rect 19708 44594 19764 44650
rect 19764 44594 19768 44650
rect 19704 44590 19768 44594
rect 19784 44650 19848 44654
rect 19784 44594 19788 44650
rect 19788 44594 19844 44650
rect 19844 44594 19848 44650
rect 19784 44590 19848 44594
rect 19864 44650 19928 44654
rect 19864 44594 19868 44650
rect 19868 44594 19924 44650
rect 19924 44594 19928 44650
rect 19864 44590 19928 44594
rect 50344 44650 50408 44654
rect 50344 44594 50348 44650
rect 50348 44594 50404 44650
rect 50404 44594 50408 44650
rect 50344 44590 50408 44594
rect 50424 44650 50488 44654
rect 50424 44594 50428 44650
rect 50428 44594 50484 44650
rect 50484 44594 50488 44650
rect 50424 44590 50488 44594
rect 50504 44650 50568 44654
rect 50504 44594 50508 44650
rect 50508 44594 50564 44650
rect 50564 44594 50568 44650
rect 50504 44590 50568 44594
rect 50584 44650 50648 44654
rect 50584 44594 50588 44650
rect 50588 44594 50644 44650
rect 50644 44594 50648 44650
rect 50584 44590 50648 44594
rect 4264 43984 4328 43988
rect 4264 43928 4268 43984
rect 4268 43928 4324 43984
rect 4324 43928 4328 43984
rect 4264 43924 4328 43928
rect 4344 43984 4408 43988
rect 4344 43928 4348 43984
rect 4348 43928 4404 43984
rect 4404 43928 4408 43984
rect 4344 43924 4408 43928
rect 4424 43984 4488 43988
rect 4424 43928 4428 43984
rect 4428 43928 4484 43984
rect 4484 43928 4488 43984
rect 4424 43924 4488 43928
rect 4504 43984 4568 43988
rect 4504 43928 4508 43984
rect 4508 43928 4564 43984
rect 4564 43928 4568 43984
rect 4504 43924 4568 43928
rect 34984 43984 35048 43988
rect 34984 43928 34988 43984
rect 34988 43928 35044 43984
rect 35044 43928 35048 43984
rect 34984 43924 35048 43928
rect 35064 43984 35128 43988
rect 35064 43928 35068 43984
rect 35068 43928 35124 43984
rect 35124 43928 35128 43984
rect 35064 43924 35128 43928
rect 35144 43984 35208 43988
rect 35144 43928 35148 43984
rect 35148 43928 35204 43984
rect 35204 43928 35208 43984
rect 35144 43924 35208 43928
rect 35224 43984 35288 43988
rect 35224 43928 35228 43984
rect 35228 43928 35284 43984
rect 35284 43928 35288 43984
rect 35224 43924 35288 43928
rect 19624 43318 19688 43322
rect 19624 43262 19628 43318
rect 19628 43262 19684 43318
rect 19684 43262 19688 43318
rect 19624 43258 19688 43262
rect 19704 43318 19768 43322
rect 19704 43262 19708 43318
rect 19708 43262 19764 43318
rect 19764 43262 19768 43318
rect 19704 43258 19768 43262
rect 19784 43318 19848 43322
rect 19784 43262 19788 43318
rect 19788 43262 19844 43318
rect 19844 43262 19848 43318
rect 19784 43258 19848 43262
rect 19864 43318 19928 43322
rect 19864 43262 19868 43318
rect 19868 43262 19924 43318
rect 19924 43262 19928 43318
rect 19864 43258 19928 43262
rect 50344 43318 50408 43322
rect 50344 43262 50348 43318
rect 50348 43262 50404 43318
rect 50404 43262 50408 43318
rect 50344 43258 50408 43262
rect 50424 43318 50488 43322
rect 50424 43262 50428 43318
rect 50428 43262 50484 43318
rect 50484 43262 50488 43318
rect 50424 43258 50488 43262
rect 50504 43318 50568 43322
rect 50504 43262 50508 43318
rect 50508 43262 50564 43318
rect 50564 43262 50568 43318
rect 50504 43258 50568 43262
rect 50584 43318 50648 43322
rect 50584 43262 50588 43318
rect 50588 43262 50644 43318
rect 50644 43262 50648 43318
rect 50584 43258 50648 43262
rect 4264 42652 4328 42656
rect 4264 42596 4268 42652
rect 4268 42596 4324 42652
rect 4324 42596 4328 42652
rect 4264 42592 4328 42596
rect 4344 42652 4408 42656
rect 4344 42596 4348 42652
rect 4348 42596 4404 42652
rect 4404 42596 4408 42652
rect 4344 42592 4408 42596
rect 4424 42652 4488 42656
rect 4424 42596 4428 42652
rect 4428 42596 4484 42652
rect 4484 42596 4488 42652
rect 4424 42592 4488 42596
rect 4504 42652 4568 42656
rect 4504 42596 4508 42652
rect 4508 42596 4564 42652
rect 4564 42596 4568 42652
rect 4504 42592 4568 42596
rect 34984 42652 35048 42656
rect 34984 42596 34988 42652
rect 34988 42596 35044 42652
rect 35044 42596 35048 42652
rect 34984 42592 35048 42596
rect 35064 42652 35128 42656
rect 35064 42596 35068 42652
rect 35068 42596 35124 42652
rect 35124 42596 35128 42652
rect 35064 42592 35128 42596
rect 35144 42652 35208 42656
rect 35144 42596 35148 42652
rect 35148 42596 35204 42652
rect 35204 42596 35208 42652
rect 35144 42592 35208 42596
rect 35224 42652 35288 42656
rect 35224 42596 35228 42652
rect 35228 42596 35284 42652
rect 35284 42596 35288 42652
rect 35224 42592 35288 42596
rect 19624 41986 19688 41990
rect 19624 41930 19628 41986
rect 19628 41930 19684 41986
rect 19684 41930 19688 41986
rect 19624 41926 19688 41930
rect 19704 41986 19768 41990
rect 19704 41930 19708 41986
rect 19708 41930 19764 41986
rect 19764 41930 19768 41986
rect 19704 41926 19768 41930
rect 19784 41986 19848 41990
rect 19784 41930 19788 41986
rect 19788 41930 19844 41986
rect 19844 41930 19848 41986
rect 19784 41926 19848 41930
rect 19864 41986 19928 41990
rect 19864 41930 19868 41986
rect 19868 41930 19924 41986
rect 19924 41930 19928 41986
rect 19864 41926 19928 41930
rect 50344 41986 50408 41990
rect 50344 41930 50348 41986
rect 50348 41930 50404 41986
rect 50404 41930 50408 41986
rect 50344 41926 50408 41930
rect 50424 41986 50488 41990
rect 50424 41930 50428 41986
rect 50428 41930 50484 41986
rect 50484 41930 50488 41986
rect 50424 41926 50488 41930
rect 50504 41986 50568 41990
rect 50504 41930 50508 41986
rect 50508 41930 50564 41986
rect 50564 41930 50568 41986
rect 50504 41926 50568 41930
rect 50584 41986 50648 41990
rect 50584 41930 50588 41986
rect 50588 41930 50644 41986
rect 50644 41930 50648 41986
rect 50584 41926 50648 41930
rect 4264 41320 4328 41324
rect 4264 41264 4268 41320
rect 4268 41264 4324 41320
rect 4324 41264 4328 41320
rect 4264 41260 4328 41264
rect 4344 41320 4408 41324
rect 4344 41264 4348 41320
rect 4348 41264 4404 41320
rect 4404 41264 4408 41320
rect 4344 41260 4408 41264
rect 4424 41320 4488 41324
rect 4424 41264 4428 41320
rect 4428 41264 4484 41320
rect 4484 41264 4488 41320
rect 4424 41260 4488 41264
rect 4504 41320 4568 41324
rect 4504 41264 4508 41320
rect 4508 41264 4564 41320
rect 4564 41264 4568 41320
rect 4504 41260 4568 41264
rect 34984 41320 35048 41324
rect 34984 41264 34988 41320
rect 34988 41264 35044 41320
rect 35044 41264 35048 41320
rect 34984 41260 35048 41264
rect 35064 41320 35128 41324
rect 35064 41264 35068 41320
rect 35068 41264 35124 41320
rect 35124 41264 35128 41320
rect 35064 41260 35128 41264
rect 35144 41320 35208 41324
rect 35144 41264 35148 41320
rect 35148 41264 35204 41320
rect 35204 41264 35208 41320
rect 35144 41260 35208 41264
rect 35224 41320 35288 41324
rect 35224 41264 35228 41320
rect 35228 41264 35284 41320
rect 35284 41264 35288 41320
rect 35224 41260 35288 41264
rect 19624 40654 19688 40658
rect 19624 40598 19628 40654
rect 19628 40598 19684 40654
rect 19684 40598 19688 40654
rect 19624 40594 19688 40598
rect 19704 40654 19768 40658
rect 19704 40598 19708 40654
rect 19708 40598 19764 40654
rect 19764 40598 19768 40654
rect 19704 40594 19768 40598
rect 19784 40654 19848 40658
rect 19784 40598 19788 40654
rect 19788 40598 19844 40654
rect 19844 40598 19848 40654
rect 19784 40594 19848 40598
rect 19864 40654 19928 40658
rect 19864 40598 19868 40654
rect 19868 40598 19924 40654
rect 19924 40598 19928 40654
rect 19864 40594 19928 40598
rect 50344 40654 50408 40658
rect 50344 40598 50348 40654
rect 50348 40598 50404 40654
rect 50404 40598 50408 40654
rect 50344 40594 50408 40598
rect 50424 40654 50488 40658
rect 50424 40598 50428 40654
rect 50428 40598 50484 40654
rect 50484 40598 50488 40654
rect 50424 40594 50488 40598
rect 50504 40654 50568 40658
rect 50504 40598 50508 40654
rect 50508 40598 50564 40654
rect 50564 40598 50568 40654
rect 50504 40594 50568 40598
rect 50584 40654 50648 40658
rect 50584 40598 50588 40654
rect 50588 40598 50644 40654
rect 50644 40598 50648 40654
rect 50584 40594 50648 40598
rect 4264 39988 4328 39992
rect 4264 39932 4268 39988
rect 4268 39932 4324 39988
rect 4324 39932 4328 39988
rect 4264 39928 4328 39932
rect 4344 39988 4408 39992
rect 4344 39932 4348 39988
rect 4348 39932 4404 39988
rect 4404 39932 4408 39988
rect 4344 39928 4408 39932
rect 4424 39988 4488 39992
rect 4424 39932 4428 39988
rect 4428 39932 4484 39988
rect 4484 39932 4488 39988
rect 4424 39928 4488 39932
rect 4504 39988 4568 39992
rect 4504 39932 4508 39988
rect 4508 39932 4564 39988
rect 4564 39932 4568 39988
rect 4504 39928 4568 39932
rect 34984 39988 35048 39992
rect 34984 39932 34988 39988
rect 34988 39932 35044 39988
rect 35044 39932 35048 39988
rect 34984 39928 35048 39932
rect 35064 39988 35128 39992
rect 35064 39932 35068 39988
rect 35068 39932 35124 39988
rect 35124 39932 35128 39988
rect 35064 39928 35128 39932
rect 35144 39988 35208 39992
rect 35144 39932 35148 39988
rect 35148 39932 35204 39988
rect 35204 39932 35208 39988
rect 35144 39928 35208 39932
rect 35224 39988 35288 39992
rect 35224 39932 35228 39988
rect 35228 39932 35284 39988
rect 35284 39932 35288 39988
rect 35224 39928 35288 39932
rect 19624 39322 19688 39326
rect 19624 39266 19628 39322
rect 19628 39266 19684 39322
rect 19684 39266 19688 39322
rect 19624 39262 19688 39266
rect 19704 39322 19768 39326
rect 19704 39266 19708 39322
rect 19708 39266 19764 39322
rect 19764 39266 19768 39322
rect 19704 39262 19768 39266
rect 19784 39322 19848 39326
rect 19784 39266 19788 39322
rect 19788 39266 19844 39322
rect 19844 39266 19848 39322
rect 19784 39262 19848 39266
rect 19864 39322 19928 39326
rect 19864 39266 19868 39322
rect 19868 39266 19924 39322
rect 19924 39266 19928 39322
rect 19864 39262 19928 39266
rect 50344 39322 50408 39326
rect 50344 39266 50348 39322
rect 50348 39266 50404 39322
rect 50404 39266 50408 39322
rect 50344 39262 50408 39266
rect 50424 39322 50488 39326
rect 50424 39266 50428 39322
rect 50428 39266 50484 39322
rect 50484 39266 50488 39322
rect 50424 39262 50488 39266
rect 50504 39322 50568 39326
rect 50504 39266 50508 39322
rect 50508 39266 50564 39322
rect 50564 39266 50568 39322
rect 50504 39262 50568 39266
rect 50584 39322 50648 39326
rect 50584 39266 50588 39322
rect 50588 39266 50644 39322
rect 50644 39266 50648 39322
rect 50584 39262 50648 39266
rect 4264 38656 4328 38660
rect 4264 38600 4268 38656
rect 4268 38600 4324 38656
rect 4324 38600 4328 38656
rect 4264 38596 4328 38600
rect 4344 38656 4408 38660
rect 4344 38600 4348 38656
rect 4348 38600 4404 38656
rect 4404 38600 4408 38656
rect 4344 38596 4408 38600
rect 4424 38656 4488 38660
rect 4424 38600 4428 38656
rect 4428 38600 4484 38656
rect 4484 38600 4488 38656
rect 4424 38596 4488 38600
rect 4504 38656 4568 38660
rect 4504 38600 4508 38656
rect 4508 38600 4564 38656
rect 4564 38600 4568 38656
rect 4504 38596 4568 38600
rect 34984 38656 35048 38660
rect 34984 38600 34988 38656
rect 34988 38600 35044 38656
rect 35044 38600 35048 38656
rect 34984 38596 35048 38600
rect 35064 38656 35128 38660
rect 35064 38600 35068 38656
rect 35068 38600 35124 38656
rect 35124 38600 35128 38656
rect 35064 38596 35128 38600
rect 35144 38656 35208 38660
rect 35144 38600 35148 38656
rect 35148 38600 35204 38656
rect 35204 38600 35208 38656
rect 35144 38596 35208 38600
rect 35224 38656 35288 38660
rect 35224 38600 35228 38656
rect 35228 38600 35284 38656
rect 35284 38600 35288 38656
rect 35224 38596 35288 38600
rect 19624 37990 19688 37994
rect 19624 37934 19628 37990
rect 19628 37934 19684 37990
rect 19684 37934 19688 37990
rect 19624 37930 19688 37934
rect 19704 37990 19768 37994
rect 19704 37934 19708 37990
rect 19708 37934 19764 37990
rect 19764 37934 19768 37990
rect 19704 37930 19768 37934
rect 19784 37990 19848 37994
rect 19784 37934 19788 37990
rect 19788 37934 19844 37990
rect 19844 37934 19848 37990
rect 19784 37930 19848 37934
rect 19864 37990 19928 37994
rect 19864 37934 19868 37990
rect 19868 37934 19924 37990
rect 19924 37934 19928 37990
rect 19864 37930 19928 37934
rect 50344 37990 50408 37994
rect 50344 37934 50348 37990
rect 50348 37934 50404 37990
rect 50404 37934 50408 37990
rect 50344 37930 50408 37934
rect 50424 37990 50488 37994
rect 50424 37934 50428 37990
rect 50428 37934 50484 37990
rect 50484 37934 50488 37990
rect 50424 37930 50488 37934
rect 50504 37990 50568 37994
rect 50504 37934 50508 37990
rect 50508 37934 50564 37990
rect 50564 37934 50568 37990
rect 50504 37930 50568 37934
rect 50584 37990 50648 37994
rect 50584 37934 50588 37990
rect 50588 37934 50644 37990
rect 50644 37934 50648 37990
rect 50584 37930 50648 37934
rect 4264 37324 4328 37328
rect 4264 37268 4268 37324
rect 4268 37268 4324 37324
rect 4324 37268 4328 37324
rect 4264 37264 4328 37268
rect 4344 37324 4408 37328
rect 4344 37268 4348 37324
rect 4348 37268 4404 37324
rect 4404 37268 4408 37324
rect 4344 37264 4408 37268
rect 4424 37324 4488 37328
rect 4424 37268 4428 37324
rect 4428 37268 4484 37324
rect 4484 37268 4488 37324
rect 4424 37264 4488 37268
rect 4504 37324 4568 37328
rect 4504 37268 4508 37324
rect 4508 37268 4564 37324
rect 4564 37268 4568 37324
rect 4504 37264 4568 37268
rect 34984 37324 35048 37328
rect 34984 37268 34988 37324
rect 34988 37268 35044 37324
rect 35044 37268 35048 37324
rect 34984 37264 35048 37268
rect 35064 37324 35128 37328
rect 35064 37268 35068 37324
rect 35068 37268 35124 37324
rect 35124 37268 35128 37324
rect 35064 37264 35128 37268
rect 35144 37324 35208 37328
rect 35144 37268 35148 37324
rect 35148 37268 35204 37324
rect 35204 37268 35208 37324
rect 35144 37264 35208 37268
rect 35224 37324 35288 37328
rect 35224 37268 35228 37324
rect 35228 37268 35284 37324
rect 35284 37268 35288 37324
rect 35224 37264 35288 37268
rect 19624 36658 19688 36662
rect 19624 36602 19628 36658
rect 19628 36602 19684 36658
rect 19684 36602 19688 36658
rect 19624 36598 19688 36602
rect 19704 36658 19768 36662
rect 19704 36602 19708 36658
rect 19708 36602 19764 36658
rect 19764 36602 19768 36658
rect 19704 36598 19768 36602
rect 19784 36658 19848 36662
rect 19784 36602 19788 36658
rect 19788 36602 19844 36658
rect 19844 36602 19848 36658
rect 19784 36598 19848 36602
rect 19864 36658 19928 36662
rect 19864 36602 19868 36658
rect 19868 36602 19924 36658
rect 19924 36602 19928 36658
rect 19864 36598 19928 36602
rect 50344 36658 50408 36662
rect 50344 36602 50348 36658
rect 50348 36602 50404 36658
rect 50404 36602 50408 36658
rect 50344 36598 50408 36602
rect 50424 36658 50488 36662
rect 50424 36602 50428 36658
rect 50428 36602 50484 36658
rect 50484 36602 50488 36658
rect 50424 36598 50488 36602
rect 50504 36658 50568 36662
rect 50504 36602 50508 36658
rect 50508 36602 50564 36658
rect 50564 36602 50568 36658
rect 50504 36598 50568 36602
rect 50584 36658 50648 36662
rect 50584 36602 50588 36658
rect 50588 36602 50644 36658
rect 50644 36602 50648 36658
rect 50584 36598 50648 36602
rect 4264 35992 4328 35996
rect 4264 35936 4268 35992
rect 4268 35936 4324 35992
rect 4324 35936 4328 35992
rect 4264 35932 4328 35936
rect 4344 35992 4408 35996
rect 4344 35936 4348 35992
rect 4348 35936 4404 35992
rect 4404 35936 4408 35992
rect 4344 35932 4408 35936
rect 4424 35992 4488 35996
rect 4424 35936 4428 35992
rect 4428 35936 4484 35992
rect 4484 35936 4488 35992
rect 4424 35932 4488 35936
rect 4504 35992 4568 35996
rect 4504 35936 4508 35992
rect 4508 35936 4564 35992
rect 4564 35936 4568 35992
rect 4504 35932 4568 35936
rect 34984 35992 35048 35996
rect 34984 35936 34988 35992
rect 34988 35936 35044 35992
rect 35044 35936 35048 35992
rect 34984 35932 35048 35936
rect 35064 35992 35128 35996
rect 35064 35936 35068 35992
rect 35068 35936 35124 35992
rect 35124 35936 35128 35992
rect 35064 35932 35128 35936
rect 35144 35992 35208 35996
rect 35144 35936 35148 35992
rect 35148 35936 35204 35992
rect 35204 35936 35208 35992
rect 35144 35932 35208 35936
rect 35224 35992 35288 35996
rect 35224 35936 35228 35992
rect 35228 35936 35284 35992
rect 35284 35936 35288 35992
rect 35224 35932 35288 35936
rect 19624 35326 19688 35330
rect 19624 35270 19628 35326
rect 19628 35270 19684 35326
rect 19684 35270 19688 35326
rect 19624 35266 19688 35270
rect 19704 35326 19768 35330
rect 19704 35270 19708 35326
rect 19708 35270 19764 35326
rect 19764 35270 19768 35326
rect 19704 35266 19768 35270
rect 19784 35326 19848 35330
rect 19784 35270 19788 35326
rect 19788 35270 19844 35326
rect 19844 35270 19848 35326
rect 19784 35266 19848 35270
rect 19864 35326 19928 35330
rect 19864 35270 19868 35326
rect 19868 35270 19924 35326
rect 19924 35270 19928 35326
rect 19864 35266 19928 35270
rect 50344 35326 50408 35330
rect 50344 35270 50348 35326
rect 50348 35270 50404 35326
rect 50404 35270 50408 35326
rect 50344 35266 50408 35270
rect 50424 35326 50488 35330
rect 50424 35270 50428 35326
rect 50428 35270 50484 35326
rect 50484 35270 50488 35326
rect 50424 35266 50488 35270
rect 50504 35326 50568 35330
rect 50504 35270 50508 35326
rect 50508 35270 50564 35326
rect 50564 35270 50568 35326
rect 50504 35266 50568 35270
rect 50584 35326 50648 35330
rect 50584 35270 50588 35326
rect 50588 35270 50644 35326
rect 50644 35270 50648 35326
rect 50584 35266 50648 35270
rect 4264 34660 4328 34664
rect 4264 34604 4268 34660
rect 4268 34604 4324 34660
rect 4324 34604 4328 34660
rect 4264 34600 4328 34604
rect 4344 34660 4408 34664
rect 4344 34604 4348 34660
rect 4348 34604 4404 34660
rect 4404 34604 4408 34660
rect 4344 34600 4408 34604
rect 4424 34660 4488 34664
rect 4424 34604 4428 34660
rect 4428 34604 4484 34660
rect 4484 34604 4488 34660
rect 4424 34600 4488 34604
rect 4504 34660 4568 34664
rect 4504 34604 4508 34660
rect 4508 34604 4564 34660
rect 4564 34604 4568 34660
rect 4504 34600 4568 34604
rect 34984 34660 35048 34664
rect 34984 34604 34988 34660
rect 34988 34604 35044 34660
rect 35044 34604 35048 34660
rect 34984 34600 35048 34604
rect 35064 34660 35128 34664
rect 35064 34604 35068 34660
rect 35068 34604 35124 34660
rect 35124 34604 35128 34660
rect 35064 34600 35128 34604
rect 35144 34660 35208 34664
rect 35144 34604 35148 34660
rect 35148 34604 35204 34660
rect 35204 34604 35208 34660
rect 35144 34600 35208 34604
rect 35224 34660 35288 34664
rect 35224 34604 35228 34660
rect 35228 34604 35284 34660
rect 35284 34604 35288 34660
rect 35224 34600 35288 34604
rect 19624 33994 19688 33998
rect 19624 33938 19628 33994
rect 19628 33938 19684 33994
rect 19684 33938 19688 33994
rect 19624 33934 19688 33938
rect 19704 33994 19768 33998
rect 19704 33938 19708 33994
rect 19708 33938 19764 33994
rect 19764 33938 19768 33994
rect 19704 33934 19768 33938
rect 19784 33994 19848 33998
rect 19784 33938 19788 33994
rect 19788 33938 19844 33994
rect 19844 33938 19848 33994
rect 19784 33934 19848 33938
rect 19864 33994 19928 33998
rect 19864 33938 19868 33994
rect 19868 33938 19924 33994
rect 19924 33938 19928 33994
rect 19864 33934 19928 33938
rect 50344 33994 50408 33998
rect 50344 33938 50348 33994
rect 50348 33938 50404 33994
rect 50404 33938 50408 33994
rect 50344 33934 50408 33938
rect 50424 33994 50488 33998
rect 50424 33938 50428 33994
rect 50428 33938 50484 33994
rect 50484 33938 50488 33994
rect 50424 33934 50488 33938
rect 50504 33994 50568 33998
rect 50504 33938 50508 33994
rect 50508 33938 50564 33994
rect 50564 33938 50568 33994
rect 50504 33934 50568 33938
rect 50584 33994 50648 33998
rect 50584 33938 50588 33994
rect 50588 33938 50644 33994
rect 50644 33938 50648 33994
rect 50584 33934 50648 33938
rect 4264 33328 4328 33332
rect 4264 33272 4268 33328
rect 4268 33272 4324 33328
rect 4324 33272 4328 33328
rect 4264 33268 4328 33272
rect 4344 33328 4408 33332
rect 4344 33272 4348 33328
rect 4348 33272 4404 33328
rect 4404 33272 4408 33328
rect 4344 33268 4408 33272
rect 4424 33328 4488 33332
rect 4424 33272 4428 33328
rect 4428 33272 4484 33328
rect 4484 33272 4488 33328
rect 4424 33268 4488 33272
rect 4504 33328 4568 33332
rect 4504 33272 4508 33328
rect 4508 33272 4564 33328
rect 4564 33272 4568 33328
rect 4504 33268 4568 33272
rect 34984 33328 35048 33332
rect 34984 33272 34988 33328
rect 34988 33272 35044 33328
rect 35044 33272 35048 33328
rect 34984 33268 35048 33272
rect 35064 33328 35128 33332
rect 35064 33272 35068 33328
rect 35068 33272 35124 33328
rect 35124 33272 35128 33328
rect 35064 33268 35128 33272
rect 35144 33328 35208 33332
rect 35144 33272 35148 33328
rect 35148 33272 35204 33328
rect 35204 33272 35208 33328
rect 35144 33268 35208 33272
rect 35224 33328 35288 33332
rect 35224 33272 35228 33328
rect 35228 33272 35284 33328
rect 35284 33272 35288 33328
rect 35224 33268 35288 33272
rect 19624 32662 19688 32666
rect 19624 32606 19628 32662
rect 19628 32606 19684 32662
rect 19684 32606 19688 32662
rect 19624 32602 19688 32606
rect 19704 32662 19768 32666
rect 19704 32606 19708 32662
rect 19708 32606 19764 32662
rect 19764 32606 19768 32662
rect 19704 32602 19768 32606
rect 19784 32662 19848 32666
rect 19784 32606 19788 32662
rect 19788 32606 19844 32662
rect 19844 32606 19848 32662
rect 19784 32602 19848 32606
rect 19864 32662 19928 32666
rect 19864 32606 19868 32662
rect 19868 32606 19924 32662
rect 19924 32606 19928 32662
rect 19864 32602 19928 32606
rect 50344 32662 50408 32666
rect 50344 32606 50348 32662
rect 50348 32606 50404 32662
rect 50404 32606 50408 32662
rect 50344 32602 50408 32606
rect 50424 32662 50488 32666
rect 50424 32606 50428 32662
rect 50428 32606 50484 32662
rect 50484 32606 50488 32662
rect 50424 32602 50488 32606
rect 50504 32662 50568 32666
rect 50504 32606 50508 32662
rect 50508 32606 50564 32662
rect 50564 32606 50568 32662
rect 50504 32602 50568 32606
rect 50584 32662 50648 32666
rect 50584 32606 50588 32662
rect 50588 32606 50644 32662
rect 50644 32606 50648 32662
rect 50584 32602 50648 32606
rect 4264 31996 4328 32000
rect 4264 31940 4268 31996
rect 4268 31940 4324 31996
rect 4324 31940 4328 31996
rect 4264 31936 4328 31940
rect 4344 31996 4408 32000
rect 4344 31940 4348 31996
rect 4348 31940 4404 31996
rect 4404 31940 4408 31996
rect 4344 31936 4408 31940
rect 4424 31996 4488 32000
rect 4424 31940 4428 31996
rect 4428 31940 4484 31996
rect 4484 31940 4488 31996
rect 4424 31936 4488 31940
rect 4504 31996 4568 32000
rect 4504 31940 4508 31996
rect 4508 31940 4564 31996
rect 4564 31940 4568 31996
rect 4504 31936 4568 31940
rect 34984 31996 35048 32000
rect 34984 31940 34988 31996
rect 34988 31940 35044 31996
rect 35044 31940 35048 31996
rect 34984 31936 35048 31940
rect 35064 31996 35128 32000
rect 35064 31940 35068 31996
rect 35068 31940 35124 31996
rect 35124 31940 35128 31996
rect 35064 31936 35128 31940
rect 35144 31996 35208 32000
rect 35144 31940 35148 31996
rect 35148 31940 35204 31996
rect 35204 31940 35208 31996
rect 35144 31936 35208 31940
rect 35224 31996 35288 32000
rect 35224 31940 35228 31996
rect 35228 31940 35284 31996
rect 35284 31940 35288 31996
rect 35224 31936 35288 31940
rect 19624 31330 19688 31334
rect 19624 31274 19628 31330
rect 19628 31274 19684 31330
rect 19684 31274 19688 31330
rect 19624 31270 19688 31274
rect 19704 31330 19768 31334
rect 19704 31274 19708 31330
rect 19708 31274 19764 31330
rect 19764 31274 19768 31330
rect 19704 31270 19768 31274
rect 19784 31330 19848 31334
rect 19784 31274 19788 31330
rect 19788 31274 19844 31330
rect 19844 31274 19848 31330
rect 19784 31270 19848 31274
rect 19864 31330 19928 31334
rect 19864 31274 19868 31330
rect 19868 31274 19924 31330
rect 19924 31274 19928 31330
rect 19864 31270 19928 31274
rect 50344 31330 50408 31334
rect 50344 31274 50348 31330
rect 50348 31274 50404 31330
rect 50404 31274 50408 31330
rect 50344 31270 50408 31274
rect 50424 31330 50488 31334
rect 50424 31274 50428 31330
rect 50428 31274 50484 31330
rect 50484 31274 50488 31330
rect 50424 31270 50488 31274
rect 50504 31330 50568 31334
rect 50504 31274 50508 31330
rect 50508 31274 50564 31330
rect 50564 31274 50568 31330
rect 50504 31270 50568 31274
rect 50584 31330 50648 31334
rect 50584 31274 50588 31330
rect 50588 31274 50644 31330
rect 50644 31274 50648 31330
rect 50584 31270 50648 31274
rect 4264 30664 4328 30668
rect 4264 30608 4268 30664
rect 4268 30608 4324 30664
rect 4324 30608 4328 30664
rect 4264 30604 4328 30608
rect 4344 30664 4408 30668
rect 4344 30608 4348 30664
rect 4348 30608 4404 30664
rect 4404 30608 4408 30664
rect 4344 30604 4408 30608
rect 4424 30664 4488 30668
rect 4424 30608 4428 30664
rect 4428 30608 4484 30664
rect 4484 30608 4488 30664
rect 4424 30604 4488 30608
rect 4504 30664 4568 30668
rect 4504 30608 4508 30664
rect 4508 30608 4564 30664
rect 4564 30608 4568 30664
rect 4504 30604 4568 30608
rect 34984 30664 35048 30668
rect 34984 30608 34988 30664
rect 34988 30608 35044 30664
rect 35044 30608 35048 30664
rect 34984 30604 35048 30608
rect 35064 30664 35128 30668
rect 35064 30608 35068 30664
rect 35068 30608 35124 30664
rect 35124 30608 35128 30664
rect 35064 30604 35128 30608
rect 35144 30664 35208 30668
rect 35144 30608 35148 30664
rect 35148 30608 35204 30664
rect 35204 30608 35208 30664
rect 35144 30604 35208 30608
rect 35224 30664 35288 30668
rect 35224 30608 35228 30664
rect 35228 30608 35284 30664
rect 35284 30608 35288 30664
rect 35224 30604 35288 30608
rect 19624 29998 19688 30002
rect 19624 29942 19628 29998
rect 19628 29942 19684 29998
rect 19684 29942 19688 29998
rect 19624 29938 19688 29942
rect 19704 29998 19768 30002
rect 19704 29942 19708 29998
rect 19708 29942 19764 29998
rect 19764 29942 19768 29998
rect 19704 29938 19768 29942
rect 19784 29998 19848 30002
rect 19784 29942 19788 29998
rect 19788 29942 19844 29998
rect 19844 29942 19848 29998
rect 19784 29938 19848 29942
rect 19864 29998 19928 30002
rect 19864 29942 19868 29998
rect 19868 29942 19924 29998
rect 19924 29942 19928 29998
rect 19864 29938 19928 29942
rect 50344 29998 50408 30002
rect 50344 29942 50348 29998
rect 50348 29942 50404 29998
rect 50404 29942 50408 29998
rect 50344 29938 50408 29942
rect 50424 29998 50488 30002
rect 50424 29942 50428 29998
rect 50428 29942 50484 29998
rect 50484 29942 50488 29998
rect 50424 29938 50488 29942
rect 50504 29998 50568 30002
rect 50504 29942 50508 29998
rect 50508 29942 50564 29998
rect 50564 29942 50568 29998
rect 50504 29938 50568 29942
rect 50584 29998 50648 30002
rect 50584 29942 50588 29998
rect 50588 29942 50644 29998
rect 50644 29942 50648 29998
rect 50584 29938 50648 29942
rect 4264 29332 4328 29336
rect 4264 29276 4268 29332
rect 4268 29276 4324 29332
rect 4324 29276 4328 29332
rect 4264 29272 4328 29276
rect 4344 29332 4408 29336
rect 4344 29276 4348 29332
rect 4348 29276 4404 29332
rect 4404 29276 4408 29332
rect 4344 29272 4408 29276
rect 4424 29332 4488 29336
rect 4424 29276 4428 29332
rect 4428 29276 4484 29332
rect 4484 29276 4488 29332
rect 4424 29272 4488 29276
rect 4504 29332 4568 29336
rect 4504 29276 4508 29332
rect 4508 29276 4564 29332
rect 4564 29276 4568 29332
rect 4504 29272 4568 29276
rect 34984 29332 35048 29336
rect 34984 29276 34988 29332
rect 34988 29276 35044 29332
rect 35044 29276 35048 29332
rect 34984 29272 35048 29276
rect 35064 29332 35128 29336
rect 35064 29276 35068 29332
rect 35068 29276 35124 29332
rect 35124 29276 35128 29332
rect 35064 29272 35128 29276
rect 35144 29332 35208 29336
rect 35144 29276 35148 29332
rect 35148 29276 35204 29332
rect 35204 29276 35208 29332
rect 35144 29272 35208 29276
rect 35224 29332 35288 29336
rect 35224 29276 35228 29332
rect 35228 29276 35284 29332
rect 35284 29276 35288 29332
rect 35224 29272 35288 29276
rect 19624 28666 19688 28670
rect 19624 28610 19628 28666
rect 19628 28610 19684 28666
rect 19684 28610 19688 28666
rect 19624 28606 19688 28610
rect 19704 28666 19768 28670
rect 19704 28610 19708 28666
rect 19708 28610 19764 28666
rect 19764 28610 19768 28666
rect 19704 28606 19768 28610
rect 19784 28666 19848 28670
rect 19784 28610 19788 28666
rect 19788 28610 19844 28666
rect 19844 28610 19848 28666
rect 19784 28606 19848 28610
rect 19864 28666 19928 28670
rect 19864 28610 19868 28666
rect 19868 28610 19924 28666
rect 19924 28610 19928 28666
rect 19864 28606 19928 28610
rect 50344 28666 50408 28670
rect 50344 28610 50348 28666
rect 50348 28610 50404 28666
rect 50404 28610 50408 28666
rect 50344 28606 50408 28610
rect 50424 28666 50488 28670
rect 50424 28610 50428 28666
rect 50428 28610 50484 28666
rect 50484 28610 50488 28666
rect 50424 28606 50488 28610
rect 50504 28666 50568 28670
rect 50504 28610 50508 28666
rect 50508 28610 50564 28666
rect 50564 28610 50568 28666
rect 50504 28606 50568 28610
rect 50584 28666 50648 28670
rect 50584 28610 50588 28666
rect 50588 28610 50644 28666
rect 50644 28610 50648 28666
rect 50584 28606 50648 28610
rect 4264 28000 4328 28004
rect 4264 27944 4268 28000
rect 4268 27944 4324 28000
rect 4324 27944 4328 28000
rect 4264 27940 4328 27944
rect 4344 28000 4408 28004
rect 4344 27944 4348 28000
rect 4348 27944 4404 28000
rect 4404 27944 4408 28000
rect 4344 27940 4408 27944
rect 4424 28000 4488 28004
rect 4424 27944 4428 28000
rect 4428 27944 4484 28000
rect 4484 27944 4488 28000
rect 4424 27940 4488 27944
rect 4504 28000 4568 28004
rect 4504 27944 4508 28000
rect 4508 27944 4564 28000
rect 4564 27944 4568 28000
rect 4504 27940 4568 27944
rect 34984 28000 35048 28004
rect 34984 27944 34988 28000
rect 34988 27944 35044 28000
rect 35044 27944 35048 28000
rect 34984 27940 35048 27944
rect 35064 28000 35128 28004
rect 35064 27944 35068 28000
rect 35068 27944 35124 28000
rect 35124 27944 35128 28000
rect 35064 27940 35128 27944
rect 35144 28000 35208 28004
rect 35144 27944 35148 28000
rect 35148 27944 35204 28000
rect 35204 27944 35208 28000
rect 35144 27940 35208 27944
rect 35224 28000 35288 28004
rect 35224 27944 35228 28000
rect 35228 27944 35284 28000
rect 35284 27944 35288 28000
rect 35224 27940 35288 27944
rect 19624 27334 19688 27338
rect 19624 27278 19628 27334
rect 19628 27278 19684 27334
rect 19684 27278 19688 27334
rect 19624 27274 19688 27278
rect 19704 27334 19768 27338
rect 19704 27278 19708 27334
rect 19708 27278 19764 27334
rect 19764 27278 19768 27334
rect 19704 27274 19768 27278
rect 19784 27334 19848 27338
rect 19784 27278 19788 27334
rect 19788 27278 19844 27334
rect 19844 27278 19848 27334
rect 19784 27274 19848 27278
rect 19864 27334 19928 27338
rect 19864 27278 19868 27334
rect 19868 27278 19924 27334
rect 19924 27278 19928 27334
rect 19864 27274 19928 27278
rect 50344 27334 50408 27338
rect 50344 27278 50348 27334
rect 50348 27278 50404 27334
rect 50404 27278 50408 27334
rect 50344 27274 50408 27278
rect 50424 27334 50488 27338
rect 50424 27278 50428 27334
rect 50428 27278 50484 27334
rect 50484 27278 50488 27334
rect 50424 27274 50488 27278
rect 50504 27334 50568 27338
rect 50504 27278 50508 27334
rect 50508 27278 50564 27334
rect 50564 27278 50568 27334
rect 50504 27274 50568 27278
rect 50584 27334 50648 27338
rect 50584 27278 50588 27334
rect 50588 27278 50644 27334
rect 50644 27278 50648 27334
rect 50584 27274 50648 27278
rect 4264 26668 4328 26672
rect 4264 26612 4268 26668
rect 4268 26612 4324 26668
rect 4324 26612 4328 26668
rect 4264 26608 4328 26612
rect 4344 26668 4408 26672
rect 4344 26612 4348 26668
rect 4348 26612 4404 26668
rect 4404 26612 4408 26668
rect 4344 26608 4408 26612
rect 4424 26668 4488 26672
rect 4424 26612 4428 26668
rect 4428 26612 4484 26668
rect 4484 26612 4488 26668
rect 4424 26608 4488 26612
rect 4504 26668 4568 26672
rect 4504 26612 4508 26668
rect 4508 26612 4564 26668
rect 4564 26612 4568 26668
rect 4504 26608 4568 26612
rect 34984 26668 35048 26672
rect 34984 26612 34988 26668
rect 34988 26612 35044 26668
rect 35044 26612 35048 26668
rect 34984 26608 35048 26612
rect 35064 26668 35128 26672
rect 35064 26612 35068 26668
rect 35068 26612 35124 26668
rect 35124 26612 35128 26668
rect 35064 26608 35128 26612
rect 35144 26668 35208 26672
rect 35144 26612 35148 26668
rect 35148 26612 35204 26668
rect 35204 26612 35208 26668
rect 35144 26608 35208 26612
rect 35224 26668 35288 26672
rect 35224 26612 35228 26668
rect 35228 26612 35284 26668
rect 35284 26612 35288 26668
rect 35224 26608 35288 26612
rect 19624 26002 19688 26006
rect 19624 25946 19628 26002
rect 19628 25946 19684 26002
rect 19684 25946 19688 26002
rect 19624 25942 19688 25946
rect 19704 26002 19768 26006
rect 19704 25946 19708 26002
rect 19708 25946 19764 26002
rect 19764 25946 19768 26002
rect 19704 25942 19768 25946
rect 19784 26002 19848 26006
rect 19784 25946 19788 26002
rect 19788 25946 19844 26002
rect 19844 25946 19848 26002
rect 19784 25942 19848 25946
rect 19864 26002 19928 26006
rect 19864 25946 19868 26002
rect 19868 25946 19924 26002
rect 19924 25946 19928 26002
rect 19864 25942 19928 25946
rect 50344 26002 50408 26006
rect 50344 25946 50348 26002
rect 50348 25946 50404 26002
rect 50404 25946 50408 26002
rect 50344 25942 50408 25946
rect 50424 26002 50488 26006
rect 50424 25946 50428 26002
rect 50428 25946 50484 26002
rect 50484 25946 50488 26002
rect 50424 25942 50488 25946
rect 50504 26002 50568 26006
rect 50504 25946 50508 26002
rect 50508 25946 50564 26002
rect 50564 25946 50568 26002
rect 50504 25942 50568 25946
rect 50584 26002 50648 26006
rect 50584 25946 50588 26002
rect 50588 25946 50644 26002
rect 50644 25946 50648 26002
rect 50584 25942 50648 25946
rect 4264 25336 4328 25340
rect 4264 25280 4268 25336
rect 4268 25280 4324 25336
rect 4324 25280 4328 25336
rect 4264 25276 4328 25280
rect 4344 25336 4408 25340
rect 4344 25280 4348 25336
rect 4348 25280 4404 25336
rect 4404 25280 4408 25336
rect 4344 25276 4408 25280
rect 4424 25336 4488 25340
rect 4424 25280 4428 25336
rect 4428 25280 4484 25336
rect 4484 25280 4488 25336
rect 4424 25276 4488 25280
rect 4504 25336 4568 25340
rect 4504 25280 4508 25336
rect 4508 25280 4564 25336
rect 4564 25280 4568 25336
rect 4504 25276 4568 25280
rect 34984 25336 35048 25340
rect 34984 25280 34988 25336
rect 34988 25280 35044 25336
rect 35044 25280 35048 25336
rect 34984 25276 35048 25280
rect 35064 25336 35128 25340
rect 35064 25280 35068 25336
rect 35068 25280 35124 25336
rect 35124 25280 35128 25336
rect 35064 25276 35128 25280
rect 35144 25336 35208 25340
rect 35144 25280 35148 25336
rect 35148 25280 35204 25336
rect 35204 25280 35208 25336
rect 35144 25276 35208 25280
rect 35224 25336 35288 25340
rect 35224 25280 35228 25336
rect 35228 25280 35284 25336
rect 35284 25280 35288 25336
rect 35224 25276 35288 25280
rect 19624 24670 19688 24674
rect 19624 24614 19628 24670
rect 19628 24614 19684 24670
rect 19684 24614 19688 24670
rect 19624 24610 19688 24614
rect 19704 24670 19768 24674
rect 19704 24614 19708 24670
rect 19708 24614 19764 24670
rect 19764 24614 19768 24670
rect 19704 24610 19768 24614
rect 19784 24670 19848 24674
rect 19784 24614 19788 24670
rect 19788 24614 19844 24670
rect 19844 24614 19848 24670
rect 19784 24610 19848 24614
rect 19864 24670 19928 24674
rect 19864 24614 19868 24670
rect 19868 24614 19924 24670
rect 19924 24614 19928 24670
rect 19864 24610 19928 24614
rect 50344 24670 50408 24674
rect 50344 24614 50348 24670
rect 50348 24614 50404 24670
rect 50404 24614 50408 24670
rect 50344 24610 50408 24614
rect 50424 24670 50488 24674
rect 50424 24614 50428 24670
rect 50428 24614 50484 24670
rect 50484 24614 50488 24670
rect 50424 24610 50488 24614
rect 50504 24670 50568 24674
rect 50504 24614 50508 24670
rect 50508 24614 50564 24670
rect 50564 24614 50568 24670
rect 50504 24610 50568 24614
rect 50584 24670 50648 24674
rect 50584 24614 50588 24670
rect 50588 24614 50644 24670
rect 50644 24614 50648 24670
rect 50584 24610 50648 24614
rect 4264 24004 4328 24008
rect 4264 23948 4268 24004
rect 4268 23948 4324 24004
rect 4324 23948 4328 24004
rect 4264 23944 4328 23948
rect 4344 24004 4408 24008
rect 4344 23948 4348 24004
rect 4348 23948 4404 24004
rect 4404 23948 4408 24004
rect 4344 23944 4408 23948
rect 4424 24004 4488 24008
rect 4424 23948 4428 24004
rect 4428 23948 4484 24004
rect 4484 23948 4488 24004
rect 4424 23944 4488 23948
rect 4504 24004 4568 24008
rect 4504 23948 4508 24004
rect 4508 23948 4564 24004
rect 4564 23948 4568 24004
rect 4504 23944 4568 23948
rect 34984 24004 35048 24008
rect 34984 23948 34988 24004
rect 34988 23948 35044 24004
rect 35044 23948 35048 24004
rect 34984 23944 35048 23948
rect 35064 24004 35128 24008
rect 35064 23948 35068 24004
rect 35068 23948 35124 24004
rect 35124 23948 35128 24004
rect 35064 23944 35128 23948
rect 35144 24004 35208 24008
rect 35144 23948 35148 24004
rect 35148 23948 35204 24004
rect 35204 23948 35208 24004
rect 35144 23944 35208 23948
rect 35224 24004 35288 24008
rect 35224 23948 35228 24004
rect 35228 23948 35284 24004
rect 35284 23948 35288 24004
rect 35224 23944 35288 23948
rect 19624 23338 19688 23342
rect 19624 23282 19628 23338
rect 19628 23282 19684 23338
rect 19684 23282 19688 23338
rect 19624 23278 19688 23282
rect 19704 23338 19768 23342
rect 19704 23282 19708 23338
rect 19708 23282 19764 23338
rect 19764 23282 19768 23338
rect 19704 23278 19768 23282
rect 19784 23338 19848 23342
rect 19784 23282 19788 23338
rect 19788 23282 19844 23338
rect 19844 23282 19848 23338
rect 19784 23278 19848 23282
rect 19864 23338 19928 23342
rect 19864 23282 19868 23338
rect 19868 23282 19924 23338
rect 19924 23282 19928 23338
rect 19864 23278 19928 23282
rect 50344 23338 50408 23342
rect 50344 23282 50348 23338
rect 50348 23282 50404 23338
rect 50404 23282 50408 23338
rect 50344 23278 50408 23282
rect 50424 23338 50488 23342
rect 50424 23282 50428 23338
rect 50428 23282 50484 23338
rect 50484 23282 50488 23338
rect 50424 23278 50488 23282
rect 50504 23338 50568 23342
rect 50504 23282 50508 23338
rect 50508 23282 50564 23338
rect 50564 23282 50568 23338
rect 50504 23278 50568 23282
rect 50584 23338 50648 23342
rect 50584 23282 50588 23338
rect 50588 23282 50644 23338
rect 50644 23282 50648 23338
rect 50584 23278 50648 23282
rect 4264 22672 4328 22676
rect 4264 22616 4268 22672
rect 4268 22616 4324 22672
rect 4324 22616 4328 22672
rect 4264 22612 4328 22616
rect 4344 22672 4408 22676
rect 4344 22616 4348 22672
rect 4348 22616 4404 22672
rect 4404 22616 4408 22672
rect 4344 22612 4408 22616
rect 4424 22672 4488 22676
rect 4424 22616 4428 22672
rect 4428 22616 4484 22672
rect 4484 22616 4488 22672
rect 4424 22612 4488 22616
rect 4504 22672 4568 22676
rect 4504 22616 4508 22672
rect 4508 22616 4564 22672
rect 4564 22616 4568 22672
rect 4504 22612 4568 22616
rect 34984 22672 35048 22676
rect 34984 22616 34988 22672
rect 34988 22616 35044 22672
rect 35044 22616 35048 22672
rect 34984 22612 35048 22616
rect 35064 22672 35128 22676
rect 35064 22616 35068 22672
rect 35068 22616 35124 22672
rect 35124 22616 35128 22672
rect 35064 22612 35128 22616
rect 35144 22672 35208 22676
rect 35144 22616 35148 22672
rect 35148 22616 35204 22672
rect 35204 22616 35208 22672
rect 35144 22612 35208 22616
rect 35224 22672 35288 22676
rect 35224 22616 35228 22672
rect 35228 22616 35284 22672
rect 35284 22616 35288 22672
rect 35224 22612 35288 22616
rect 19624 22006 19688 22010
rect 19624 21950 19628 22006
rect 19628 21950 19684 22006
rect 19684 21950 19688 22006
rect 19624 21946 19688 21950
rect 19704 22006 19768 22010
rect 19704 21950 19708 22006
rect 19708 21950 19764 22006
rect 19764 21950 19768 22006
rect 19704 21946 19768 21950
rect 19784 22006 19848 22010
rect 19784 21950 19788 22006
rect 19788 21950 19844 22006
rect 19844 21950 19848 22006
rect 19784 21946 19848 21950
rect 19864 22006 19928 22010
rect 19864 21950 19868 22006
rect 19868 21950 19924 22006
rect 19924 21950 19928 22006
rect 19864 21946 19928 21950
rect 50344 22006 50408 22010
rect 50344 21950 50348 22006
rect 50348 21950 50404 22006
rect 50404 21950 50408 22006
rect 50344 21946 50408 21950
rect 50424 22006 50488 22010
rect 50424 21950 50428 22006
rect 50428 21950 50484 22006
rect 50484 21950 50488 22006
rect 50424 21946 50488 21950
rect 50504 22006 50568 22010
rect 50504 21950 50508 22006
rect 50508 21950 50564 22006
rect 50564 21950 50568 22006
rect 50504 21946 50568 21950
rect 50584 22006 50648 22010
rect 50584 21950 50588 22006
rect 50588 21950 50644 22006
rect 50644 21950 50648 22006
rect 50584 21946 50648 21950
rect 4264 21340 4328 21344
rect 4264 21284 4268 21340
rect 4268 21284 4324 21340
rect 4324 21284 4328 21340
rect 4264 21280 4328 21284
rect 4344 21340 4408 21344
rect 4344 21284 4348 21340
rect 4348 21284 4404 21340
rect 4404 21284 4408 21340
rect 4344 21280 4408 21284
rect 4424 21340 4488 21344
rect 4424 21284 4428 21340
rect 4428 21284 4484 21340
rect 4484 21284 4488 21340
rect 4424 21280 4488 21284
rect 4504 21340 4568 21344
rect 4504 21284 4508 21340
rect 4508 21284 4564 21340
rect 4564 21284 4568 21340
rect 4504 21280 4568 21284
rect 34984 21340 35048 21344
rect 34984 21284 34988 21340
rect 34988 21284 35044 21340
rect 35044 21284 35048 21340
rect 34984 21280 35048 21284
rect 35064 21340 35128 21344
rect 35064 21284 35068 21340
rect 35068 21284 35124 21340
rect 35124 21284 35128 21340
rect 35064 21280 35128 21284
rect 35144 21340 35208 21344
rect 35144 21284 35148 21340
rect 35148 21284 35204 21340
rect 35204 21284 35208 21340
rect 35144 21280 35208 21284
rect 35224 21340 35288 21344
rect 35224 21284 35228 21340
rect 35228 21284 35284 21340
rect 35284 21284 35288 21340
rect 35224 21280 35288 21284
rect 19624 20674 19688 20678
rect 19624 20618 19628 20674
rect 19628 20618 19684 20674
rect 19684 20618 19688 20674
rect 19624 20614 19688 20618
rect 19704 20674 19768 20678
rect 19704 20618 19708 20674
rect 19708 20618 19764 20674
rect 19764 20618 19768 20674
rect 19704 20614 19768 20618
rect 19784 20674 19848 20678
rect 19784 20618 19788 20674
rect 19788 20618 19844 20674
rect 19844 20618 19848 20674
rect 19784 20614 19848 20618
rect 19864 20674 19928 20678
rect 19864 20618 19868 20674
rect 19868 20618 19924 20674
rect 19924 20618 19928 20674
rect 19864 20614 19928 20618
rect 50344 20674 50408 20678
rect 50344 20618 50348 20674
rect 50348 20618 50404 20674
rect 50404 20618 50408 20674
rect 50344 20614 50408 20618
rect 50424 20674 50488 20678
rect 50424 20618 50428 20674
rect 50428 20618 50484 20674
rect 50484 20618 50488 20674
rect 50424 20614 50488 20618
rect 50504 20674 50568 20678
rect 50504 20618 50508 20674
rect 50508 20618 50564 20674
rect 50564 20618 50568 20674
rect 50504 20614 50568 20618
rect 50584 20674 50648 20678
rect 50584 20618 50588 20674
rect 50588 20618 50644 20674
rect 50644 20618 50648 20674
rect 50584 20614 50648 20618
rect 4264 20008 4328 20012
rect 4264 19952 4268 20008
rect 4268 19952 4324 20008
rect 4324 19952 4328 20008
rect 4264 19948 4328 19952
rect 4344 20008 4408 20012
rect 4344 19952 4348 20008
rect 4348 19952 4404 20008
rect 4404 19952 4408 20008
rect 4344 19948 4408 19952
rect 4424 20008 4488 20012
rect 4424 19952 4428 20008
rect 4428 19952 4484 20008
rect 4484 19952 4488 20008
rect 4424 19948 4488 19952
rect 4504 20008 4568 20012
rect 4504 19952 4508 20008
rect 4508 19952 4564 20008
rect 4564 19952 4568 20008
rect 4504 19948 4568 19952
rect 34984 20008 35048 20012
rect 34984 19952 34988 20008
rect 34988 19952 35044 20008
rect 35044 19952 35048 20008
rect 34984 19948 35048 19952
rect 35064 20008 35128 20012
rect 35064 19952 35068 20008
rect 35068 19952 35124 20008
rect 35124 19952 35128 20008
rect 35064 19948 35128 19952
rect 35144 20008 35208 20012
rect 35144 19952 35148 20008
rect 35148 19952 35204 20008
rect 35204 19952 35208 20008
rect 35144 19948 35208 19952
rect 35224 20008 35288 20012
rect 35224 19952 35228 20008
rect 35228 19952 35284 20008
rect 35284 19952 35288 20008
rect 35224 19948 35288 19952
rect 19624 19342 19688 19346
rect 19624 19286 19628 19342
rect 19628 19286 19684 19342
rect 19684 19286 19688 19342
rect 19624 19282 19688 19286
rect 19704 19342 19768 19346
rect 19704 19286 19708 19342
rect 19708 19286 19764 19342
rect 19764 19286 19768 19342
rect 19704 19282 19768 19286
rect 19784 19342 19848 19346
rect 19784 19286 19788 19342
rect 19788 19286 19844 19342
rect 19844 19286 19848 19342
rect 19784 19282 19848 19286
rect 19864 19342 19928 19346
rect 19864 19286 19868 19342
rect 19868 19286 19924 19342
rect 19924 19286 19928 19342
rect 19864 19282 19928 19286
rect 50344 19342 50408 19346
rect 50344 19286 50348 19342
rect 50348 19286 50404 19342
rect 50404 19286 50408 19342
rect 50344 19282 50408 19286
rect 50424 19342 50488 19346
rect 50424 19286 50428 19342
rect 50428 19286 50484 19342
rect 50484 19286 50488 19342
rect 50424 19282 50488 19286
rect 50504 19342 50568 19346
rect 50504 19286 50508 19342
rect 50508 19286 50564 19342
rect 50564 19286 50568 19342
rect 50504 19282 50568 19286
rect 50584 19342 50648 19346
rect 50584 19286 50588 19342
rect 50588 19286 50644 19342
rect 50644 19286 50648 19342
rect 50584 19282 50648 19286
rect 4264 18676 4328 18680
rect 4264 18620 4268 18676
rect 4268 18620 4324 18676
rect 4324 18620 4328 18676
rect 4264 18616 4328 18620
rect 4344 18676 4408 18680
rect 4344 18620 4348 18676
rect 4348 18620 4404 18676
rect 4404 18620 4408 18676
rect 4344 18616 4408 18620
rect 4424 18676 4488 18680
rect 4424 18620 4428 18676
rect 4428 18620 4484 18676
rect 4484 18620 4488 18676
rect 4424 18616 4488 18620
rect 4504 18676 4568 18680
rect 4504 18620 4508 18676
rect 4508 18620 4564 18676
rect 4564 18620 4568 18676
rect 4504 18616 4568 18620
rect 34984 18676 35048 18680
rect 34984 18620 34988 18676
rect 34988 18620 35044 18676
rect 35044 18620 35048 18676
rect 34984 18616 35048 18620
rect 35064 18676 35128 18680
rect 35064 18620 35068 18676
rect 35068 18620 35124 18676
rect 35124 18620 35128 18676
rect 35064 18616 35128 18620
rect 35144 18676 35208 18680
rect 35144 18620 35148 18676
rect 35148 18620 35204 18676
rect 35204 18620 35208 18676
rect 35144 18616 35208 18620
rect 35224 18676 35288 18680
rect 35224 18620 35228 18676
rect 35228 18620 35284 18676
rect 35284 18620 35288 18676
rect 35224 18616 35288 18620
rect 19624 18010 19688 18014
rect 19624 17954 19628 18010
rect 19628 17954 19684 18010
rect 19684 17954 19688 18010
rect 19624 17950 19688 17954
rect 19704 18010 19768 18014
rect 19704 17954 19708 18010
rect 19708 17954 19764 18010
rect 19764 17954 19768 18010
rect 19704 17950 19768 17954
rect 19784 18010 19848 18014
rect 19784 17954 19788 18010
rect 19788 17954 19844 18010
rect 19844 17954 19848 18010
rect 19784 17950 19848 17954
rect 19864 18010 19928 18014
rect 19864 17954 19868 18010
rect 19868 17954 19924 18010
rect 19924 17954 19928 18010
rect 19864 17950 19928 17954
rect 50344 18010 50408 18014
rect 50344 17954 50348 18010
rect 50348 17954 50404 18010
rect 50404 17954 50408 18010
rect 50344 17950 50408 17954
rect 50424 18010 50488 18014
rect 50424 17954 50428 18010
rect 50428 17954 50484 18010
rect 50484 17954 50488 18010
rect 50424 17950 50488 17954
rect 50504 18010 50568 18014
rect 50504 17954 50508 18010
rect 50508 17954 50564 18010
rect 50564 17954 50568 18010
rect 50504 17950 50568 17954
rect 50584 18010 50648 18014
rect 50584 17954 50588 18010
rect 50588 17954 50644 18010
rect 50644 17954 50648 18010
rect 50584 17950 50648 17954
rect 4264 17344 4328 17348
rect 4264 17288 4268 17344
rect 4268 17288 4324 17344
rect 4324 17288 4328 17344
rect 4264 17284 4328 17288
rect 4344 17344 4408 17348
rect 4344 17288 4348 17344
rect 4348 17288 4404 17344
rect 4404 17288 4408 17344
rect 4344 17284 4408 17288
rect 4424 17344 4488 17348
rect 4424 17288 4428 17344
rect 4428 17288 4484 17344
rect 4484 17288 4488 17344
rect 4424 17284 4488 17288
rect 4504 17344 4568 17348
rect 4504 17288 4508 17344
rect 4508 17288 4564 17344
rect 4564 17288 4568 17344
rect 4504 17284 4568 17288
rect 34984 17344 35048 17348
rect 34984 17288 34988 17344
rect 34988 17288 35044 17344
rect 35044 17288 35048 17344
rect 34984 17284 35048 17288
rect 35064 17344 35128 17348
rect 35064 17288 35068 17344
rect 35068 17288 35124 17344
rect 35124 17288 35128 17344
rect 35064 17284 35128 17288
rect 35144 17344 35208 17348
rect 35144 17288 35148 17344
rect 35148 17288 35204 17344
rect 35204 17288 35208 17344
rect 35144 17284 35208 17288
rect 35224 17344 35288 17348
rect 35224 17288 35228 17344
rect 35228 17288 35284 17344
rect 35284 17288 35288 17344
rect 35224 17284 35288 17288
rect 19624 16678 19688 16682
rect 19624 16622 19628 16678
rect 19628 16622 19684 16678
rect 19684 16622 19688 16678
rect 19624 16618 19688 16622
rect 19704 16678 19768 16682
rect 19704 16622 19708 16678
rect 19708 16622 19764 16678
rect 19764 16622 19768 16678
rect 19704 16618 19768 16622
rect 19784 16678 19848 16682
rect 19784 16622 19788 16678
rect 19788 16622 19844 16678
rect 19844 16622 19848 16678
rect 19784 16618 19848 16622
rect 19864 16678 19928 16682
rect 19864 16622 19868 16678
rect 19868 16622 19924 16678
rect 19924 16622 19928 16678
rect 19864 16618 19928 16622
rect 50344 16678 50408 16682
rect 50344 16622 50348 16678
rect 50348 16622 50404 16678
rect 50404 16622 50408 16678
rect 50344 16618 50408 16622
rect 50424 16678 50488 16682
rect 50424 16622 50428 16678
rect 50428 16622 50484 16678
rect 50484 16622 50488 16678
rect 50424 16618 50488 16622
rect 50504 16678 50568 16682
rect 50504 16622 50508 16678
rect 50508 16622 50564 16678
rect 50564 16622 50568 16678
rect 50504 16618 50568 16622
rect 50584 16678 50648 16682
rect 50584 16622 50588 16678
rect 50588 16622 50644 16678
rect 50644 16622 50648 16678
rect 50584 16618 50648 16622
rect 4264 16012 4328 16016
rect 4264 15956 4268 16012
rect 4268 15956 4324 16012
rect 4324 15956 4328 16012
rect 4264 15952 4328 15956
rect 4344 16012 4408 16016
rect 4344 15956 4348 16012
rect 4348 15956 4404 16012
rect 4404 15956 4408 16012
rect 4344 15952 4408 15956
rect 4424 16012 4488 16016
rect 4424 15956 4428 16012
rect 4428 15956 4484 16012
rect 4484 15956 4488 16012
rect 4424 15952 4488 15956
rect 4504 16012 4568 16016
rect 4504 15956 4508 16012
rect 4508 15956 4564 16012
rect 4564 15956 4568 16012
rect 4504 15952 4568 15956
rect 34984 16012 35048 16016
rect 34984 15956 34988 16012
rect 34988 15956 35044 16012
rect 35044 15956 35048 16012
rect 34984 15952 35048 15956
rect 35064 16012 35128 16016
rect 35064 15956 35068 16012
rect 35068 15956 35124 16012
rect 35124 15956 35128 16012
rect 35064 15952 35128 15956
rect 35144 16012 35208 16016
rect 35144 15956 35148 16012
rect 35148 15956 35204 16012
rect 35204 15956 35208 16012
rect 35144 15952 35208 15956
rect 35224 16012 35288 16016
rect 35224 15956 35228 16012
rect 35228 15956 35284 16012
rect 35284 15956 35288 16012
rect 35224 15952 35288 15956
rect 19624 15346 19688 15350
rect 19624 15290 19628 15346
rect 19628 15290 19684 15346
rect 19684 15290 19688 15346
rect 19624 15286 19688 15290
rect 19704 15346 19768 15350
rect 19704 15290 19708 15346
rect 19708 15290 19764 15346
rect 19764 15290 19768 15346
rect 19704 15286 19768 15290
rect 19784 15346 19848 15350
rect 19784 15290 19788 15346
rect 19788 15290 19844 15346
rect 19844 15290 19848 15346
rect 19784 15286 19848 15290
rect 19864 15346 19928 15350
rect 19864 15290 19868 15346
rect 19868 15290 19924 15346
rect 19924 15290 19928 15346
rect 19864 15286 19928 15290
rect 50344 15346 50408 15350
rect 50344 15290 50348 15346
rect 50348 15290 50404 15346
rect 50404 15290 50408 15346
rect 50344 15286 50408 15290
rect 50424 15346 50488 15350
rect 50424 15290 50428 15346
rect 50428 15290 50484 15346
rect 50484 15290 50488 15346
rect 50424 15286 50488 15290
rect 50504 15346 50568 15350
rect 50504 15290 50508 15346
rect 50508 15290 50564 15346
rect 50564 15290 50568 15346
rect 50504 15286 50568 15290
rect 50584 15346 50648 15350
rect 50584 15290 50588 15346
rect 50588 15290 50644 15346
rect 50644 15290 50648 15346
rect 50584 15286 50648 15290
rect 4264 14680 4328 14684
rect 4264 14624 4268 14680
rect 4268 14624 4324 14680
rect 4324 14624 4328 14680
rect 4264 14620 4328 14624
rect 4344 14680 4408 14684
rect 4344 14624 4348 14680
rect 4348 14624 4404 14680
rect 4404 14624 4408 14680
rect 4344 14620 4408 14624
rect 4424 14680 4488 14684
rect 4424 14624 4428 14680
rect 4428 14624 4484 14680
rect 4484 14624 4488 14680
rect 4424 14620 4488 14624
rect 4504 14680 4568 14684
rect 4504 14624 4508 14680
rect 4508 14624 4564 14680
rect 4564 14624 4568 14680
rect 4504 14620 4568 14624
rect 34984 14680 35048 14684
rect 34984 14624 34988 14680
rect 34988 14624 35044 14680
rect 35044 14624 35048 14680
rect 34984 14620 35048 14624
rect 35064 14680 35128 14684
rect 35064 14624 35068 14680
rect 35068 14624 35124 14680
rect 35124 14624 35128 14680
rect 35064 14620 35128 14624
rect 35144 14680 35208 14684
rect 35144 14624 35148 14680
rect 35148 14624 35204 14680
rect 35204 14624 35208 14680
rect 35144 14620 35208 14624
rect 35224 14680 35288 14684
rect 35224 14624 35228 14680
rect 35228 14624 35284 14680
rect 35284 14624 35288 14680
rect 35224 14620 35288 14624
rect 19624 14014 19688 14018
rect 19624 13958 19628 14014
rect 19628 13958 19684 14014
rect 19684 13958 19688 14014
rect 19624 13954 19688 13958
rect 19704 14014 19768 14018
rect 19704 13958 19708 14014
rect 19708 13958 19764 14014
rect 19764 13958 19768 14014
rect 19704 13954 19768 13958
rect 19784 14014 19848 14018
rect 19784 13958 19788 14014
rect 19788 13958 19844 14014
rect 19844 13958 19848 14014
rect 19784 13954 19848 13958
rect 19864 14014 19928 14018
rect 19864 13958 19868 14014
rect 19868 13958 19924 14014
rect 19924 13958 19928 14014
rect 19864 13954 19928 13958
rect 50344 14014 50408 14018
rect 50344 13958 50348 14014
rect 50348 13958 50404 14014
rect 50404 13958 50408 14014
rect 50344 13954 50408 13958
rect 50424 14014 50488 14018
rect 50424 13958 50428 14014
rect 50428 13958 50484 14014
rect 50484 13958 50488 14014
rect 50424 13954 50488 13958
rect 50504 14014 50568 14018
rect 50504 13958 50508 14014
rect 50508 13958 50564 14014
rect 50564 13958 50568 14014
rect 50504 13954 50568 13958
rect 50584 14014 50648 14018
rect 50584 13958 50588 14014
rect 50588 13958 50644 14014
rect 50644 13958 50648 14014
rect 50584 13954 50648 13958
rect 4264 13348 4328 13352
rect 4264 13292 4268 13348
rect 4268 13292 4324 13348
rect 4324 13292 4328 13348
rect 4264 13288 4328 13292
rect 4344 13348 4408 13352
rect 4344 13292 4348 13348
rect 4348 13292 4404 13348
rect 4404 13292 4408 13348
rect 4344 13288 4408 13292
rect 4424 13348 4488 13352
rect 4424 13292 4428 13348
rect 4428 13292 4484 13348
rect 4484 13292 4488 13348
rect 4424 13288 4488 13292
rect 4504 13348 4568 13352
rect 4504 13292 4508 13348
rect 4508 13292 4564 13348
rect 4564 13292 4568 13348
rect 4504 13288 4568 13292
rect 34984 13348 35048 13352
rect 34984 13292 34988 13348
rect 34988 13292 35044 13348
rect 35044 13292 35048 13348
rect 34984 13288 35048 13292
rect 35064 13348 35128 13352
rect 35064 13292 35068 13348
rect 35068 13292 35124 13348
rect 35124 13292 35128 13348
rect 35064 13288 35128 13292
rect 35144 13348 35208 13352
rect 35144 13292 35148 13348
rect 35148 13292 35204 13348
rect 35204 13292 35208 13348
rect 35144 13288 35208 13292
rect 35224 13348 35288 13352
rect 35224 13292 35228 13348
rect 35228 13292 35284 13348
rect 35284 13292 35288 13348
rect 35224 13288 35288 13292
rect 19624 12682 19688 12686
rect 19624 12626 19628 12682
rect 19628 12626 19684 12682
rect 19684 12626 19688 12682
rect 19624 12622 19688 12626
rect 19704 12682 19768 12686
rect 19704 12626 19708 12682
rect 19708 12626 19764 12682
rect 19764 12626 19768 12682
rect 19704 12622 19768 12626
rect 19784 12682 19848 12686
rect 19784 12626 19788 12682
rect 19788 12626 19844 12682
rect 19844 12626 19848 12682
rect 19784 12622 19848 12626
rect 19864 12682 19928 12686
rect 19864 12626 19868 12682
rect 19868 12626 19924 12682
rect 19924 12626 19928 12682
rect 19864 12622 19928 12626
rect 50344 12682 50408 12686
rect 50344 12626 50348 12682
rect 50348 12626 50404 12682
rect 50404 12626 50408 12682
rect 50344 12622 50408 12626
rect 50424 12682 50488 12686
rect 50424 12626 50428 12682
rect 50428 12626 50484 12682
rect 50484 12626 50488 12682
rect 50424 12622 50488 12626
rect 50504 12682 50568 12686
rect 50504 12626 50508 12682
rect 50508 12626 50564 12682
rect 50564 12626 50568 12682
rect 50504 12622 50568 12626
rect 50584 12682 50648 12686
rect 50584 12626 50588 12682
rect 50588 12626 50644 12682
rect 50644 12626 50648 12682
rect 50584 12622 50648 12626
rect 4264 12016 4328 12020
rect 4264 11960 4268 12016
rect 4268 11960 4324 12016
rect 4324 11960 4328 12016
rect 4264 11956 4328 11960
rect 4344 12016 4408 12020
rect 4344 11960 4348 12016
rect 4348 11960 4404 12016
rect 4404 11960 4408 12016
rect 4344 11956 4408 11960
rect 4424 12016 4488 12020
rect 4424 11960 4428 12016
rect 4428 11960 4484 12016
rect 4484 11960 4488 12016
rect 4424 11956 4488 11960
rect 4504 12016 4568 12020
rect 4504 11960 4508 12016
rect 4508 11960 4564 12016
rect 4564 11960 4568 12016
rect 4504 11956 4568 11960
rect 34984 12016 35048 12020
rect 34984 11960 34988 12016
rect 34988 11960 35044 12016
rect 35044 11960 35048 12016
rect 34984 11956 35048 11960
rect 35064 12016 35128 12020
rect 35064 11960 35068 12016
rect 35068 11960 35124 12016
rect 35124 11960 35128 12016
rect 35064 11956 35128 11960
rect 35144 12016 35208 12020
rect 35144 11960 35148 12016
rect 35148 11960 35204 12016
rect 35204 11960 35208 12016
rect 35144 11956 35208 11960
rect 35224 12016 35288 12020
rect 35224 11960 35228 12016
rect 35228 11960 35284 12016
rect 35284 11960 35288 12016
rect 35224 11956 35288 11960
rect 19624 11350 19688 11354
rect 19624 11294 19628 11350
rect 19628 11294 19684 11350
rect 19684 11294 19688 11350
rect 19624 11290 19688 11294
rect 19704 11350 19768 11354
rect 19704 11294 19708 11350
rect 19708 11294 19764 11350
rect 19764 11294 19768 11350
rect 19704 11290 19768 11294
rect 19784 11350 19848 11354
rect 19784 11294 19788 11350
rect 19788 11294 19844 11350
rect 19844 11294 19848 11350
rect 19784 11290 19848 11294
rect 19864 11350 19928 11354
rect 19864 11294 19868 11350
rect 19868 11294 19924 11350
rect 19924 11294 19928 11350
rect 19864 11290 19928 11294
rect 50344 11350 50408 11354
rect 50344 11294 50348 11350
rect 50348 11294 50404 11350
rect 50404 11294 50408 11350
rect 50344 11290 50408 11294
rect 50424 11350 50488 11354
rect 50424 11294 50428 11350
rect 50428 11294 50484 11350
rect 50484 11294 50488 11350
rect 50424 11290 50488 11294
rect 50504 11350 50568 11354
rect 50504 11294 50508 11350
rect 50508 11294 50564 11350
rect 50564 11294 50568 11350
rect 50504 11290 50568 11294
rect 50584 11350 50648 11354
rect 50584 11294 50588 11350
rect 50588 11294 50644 11350
rect 50644 11294 50648 11350
rect 50584 11290 50648 11294
rect 4264 10684 4328 10688
rect 4264 10628 4268 10684
rect 4268 10628 4324 10684
rect 4324 10628 4328 10684
rect 4264 10624 4328 10628
rect 4344 10684 4408 10688
rect 4344 10628 4348 10684
rect 4348 10628 4404 10684
rect 4404 10628 4408 10684
rect 4344 10624 4408 10628
rect 4424 10684 4488 10688
rect 4424 10628 4428 10684
rect 4428 10628 4484 10684
rect 4484 10628 4488 10684
rect 4424 10624 4488 10628
rect 4504 10684 4568 10688
rect 4504 10628 4508 10684
rect 4508 10628 4564 10684
rect 4564 10628 4568 10684
rect 4504 10624 4568 10628
rect 34984 10684 35048 10688
rect 34984 10628 34988 10684
rect 34988 10628 35044 10684
rect 35044 10628 35048 10684
rect 34984 10624 35048 10628
rect 35064 10684 35128 10688
rect 35064 10628 35068 10684
rect 35068 10628 35124 10684
rect 35124 10628 35128 10684
rect 35064 10624 35128 10628
rect 35144 10684 35208 10688
rect 35144 10628 35148 10684
rect 35148 10628 35204 10684
rect 35204 10628 35208 10684
rect 35144 10624 35208 10628
rect 35224 10684 35288 10688
rect 35224 10628 35228 10684
rect 35228 10628 35284 10684
rect 35284 10628 35288 10684
rect 35224 10624 35288 10628
rect 19624 10018 19688 10022
rect 19624 9962 19628 10018
rect 19628 9962 19684 10018
rect 19684 9962 19688 10018
rect 19624 9958 19688 9962
rect 19704 10018 19768 10022
rect 19704 9962 19708 10018
rect 19708 9962 19764 10018
rect 19764 9962 19768 10018
rect 19704 9958 19768 9962
rect 19784 10018 19848 10022
rect 19784 9962 19788 10018
rect 19788 9962 19844 10018
rect 19844 9962 19848 10018
rect 19784 9958 19848 9962
rect 19864 10018 19928 10022
rect 19864 9962 19868 10018
rect 19868 9962 19924 10018
rect 19924 9962 19928 10018
rect 19864 9958 19928 9962
rect 50344 10018 50408 10022
rect 50344 9962 50348 10018
rect 50348 9962 50404 10018
rect 50404 9962 50408 10018
rect 50344 9958 50408 9962
rect 50424 10018 50488 10022
rect 50424 9962 50428 10018
rect 50428 9962 50484 10018
rect 50484 9962 50488 10018
rect 50424 9958 50488 9962
rect 50504 10018 50568 10022
rect 50504 9962 50508 10018
rect 50508 9962 50564 10018
rect 50564 9962 50568 10018
rect 50504 9958 50568 9962
rect 50584 10018 50648 10022
rect 50584 9962 50588 10018
rect 50588 9962 50644 10018
rect 50644 9962 50648 10018
rect 50584 9958 50648 9962
rect 4264 9352 4328 9356
rect 4264 9296 4268 9352
rect 4268 9296 4324 9352
rect 4324 9296 4328 9352
rect 4264 9292 4328 9296
rect 4344 9352 4408 9356
rect 4344 9296 4348 9352
rect 4348 9296 4404 9352
rect 4404 9296 4408 9352
rect 4344 9292 4408 9296
rect 4424 9352 4488 9356
rect 4424 9296 4428 9352
rect 4428 9296 4484 9352
rect 4484 9296 4488 9352
rect 4424 9292 4488 9296
rect 4504 9352 4568 9356
rect 4504 9296 4508 9352
rect 4508 9296 4564 9352
rect 4564 9296 4568 9352
rect 4504 9292 4568 9296
rect 34984 9352 35048 9356
rect 34984 9296 34988 9352
rect 34988 9296 35044 9352
rect 35044 9296 35048 9352
rect 34984 9292 35048 9296
rect 35064 9352 35128 9356
rect 35064 9296 35068 9352
rect 35068 9296 35124 9352
rect 35124 9296 35128 9352
rect 35064 9292 35128 9296
rect 35144 9352 35208 9356
rect 35144 9296 35148 9352
rect 35148 9296 35204 9352
rect 35204 9296 35208 9352
rect 35144 9292 35208 9296
rect 35224 9352 35288 9356
rect 35224 9296 35228 9352
rect 35228 9296 35284 9352
rect 35284 9296 35288 9352
rect 35224 9292 35288 9296
rect 19624 8686 19688 8690
rect 19624 8630 19628 8686
rect 19628 8630 19684 8686
rect 19684 8630 19688 8686
rect 19624 8626 19688 8630
rect 19704 8686 19768 8690
rect 19704 8630 19708 8686
rect 19708 8630 19764 8686
rect 19764 8630 19768 8686
rect 19704 8626 19768 8630
rect 19784 8686 19848 8690
rect 19784 8630 19788 8686
rect 19788 8630 19844 8686
rect 19844 8630 19848 8686
rect 19784 8626 19848 8630
rect 19864 8686 19928 8690
rect 19864 8630 19868 8686
rect 19868 8630 19924 8686
rect 19924 8630 19928 8686
rect 19864 8626 19928 8630
rect 50344 8686 50408 8690
rect 50344 8630 50348 8686
rect 50348 8630 50404 8686
rect 50404 8630 50408 8686
rect 50344 8626 50408 8630
rect 50424 8686 50488 8690
rect 50424 8630 50428 8686
rect 50428 8630 50484 8686
rect 50484 8630 50488 8686
rect 50424 8626 50488 8630
rect 50504 8686 50568 8690
rect 50504 8630 50508 8686
rect 50508 8630 50564 8686
rect 50564 8630 50568 8686
rect 50504 8626 50568 8630
rect 50584 8686 50648 8690
rect 50584 8630 50588 8686
rect 50588 8630 50644 8686
rect 50644 8630 50648 8686
rect 50584 8626 50648 8630
rect 4264 8020 4328 8024
rect 4264 7964 4268 8020
rect 4268 7964 4324 8020
rect 4324 7964 4328 8020
rect 4264 7960 4328 7964
rect 4344 8020 4408 8024
rect 4344 7964 4348 8020
rect 4348 7964 4404 8020
rect 4404 7964 4408 8020
rect 4344 7960 4408 7964
rect 4424 8020 4488 8024
rect 4424 7964 4428 8020
rect 4428 7964 4484 8020
rect 4484 7964 4488 8020
rect 4424 7960 4488 7964
rect 4504 8020 4568 8024
rect 4504 7964 4508 8020
rect 4508 7964 4564 8020
rect 4564 7964 4568 8020
rect 4504 7960 4568 7964
rect 34984 8020 35048 8024
rect 34984 7964 34988 8020
rect 34988 7964 35044 8020
rect 35044 7964 35048 8020
rect 34984 7960 35048 7964
rect 35064 8020 35128 8024
rect 35064 7964 35068 8020
rect 35068 7964 35124 8020
rect 35124 7964 35128 8020
rect 35064 7960 35128 7964
rect 35144 8020 35208 8024
rect 35144 7964 35148 8020
rect 35148 7964 35204 8020
rect 35204 7964 35208 8020
rect 35144 7960 35208 7964
rect 35224 8020 35288 8024
rect 35224 7964 35228 8020
rect 35228 7964 35284 8020
rect 35284 7964 35288 8020
rect 35224 7960 35288 7964
rect 19624 7354 19688 7358
rect 19624 7298 19628 7354
rect 19628 7298 19684 7354
rect 19684 7298 19688 7354
rect 19624 7294 19688 7298
rect 19704 7354 19768 7358
rect 19704 7298 19708 7354
rect 19708 7298 19764 7354
rect 19764 7298 19768 7354
rect 19704 7294 19768 7298
rect 19784 7354 19848 7358
rect 19784 7298 19788 7354
rect 19788 7298 19844 7354
rect 19844 7298 19848 7354
rect 19784 7294 19848 7298
rect 19864 7354 19928 7358
rect 19864 7298 19868 7354
rect 19868 7298 19924 7354
rect 19924 7298 19928 7354
rect 19864 7294 19928 7298
rect 50344 7354 50408 7358
rect 50344 7298 50348 7354
rect 50348 7298 50404 7354
rect 50404 7298 50408 7354
rect 50344 7294 50408 7298
rect 50424 7354 50488 7358
rect 50424 7298 50428 7354
rect 50428 7298 50484 7354
rect 50484 7298 50488 7354
rect 50424 7294 50488 7298
rect 50504 7354 50568 7358
rect 50504 7298 50508 7354
rect 50508 7298 50564 7354
rect 50564 7298 50568 7354
rect 50504 7294 50568 7298
rect 50584 7354 50648 7358
rect 50584 7298 50588 7354
rect 50588 7298 50644 7354
rect 50644 7298 50648 7354
rect 50584 7294 50648 7298
rect 4264 6688 4328 6692
rect 4264 6632 4268 6688
rect 4268 6632 4324 6688
rect 4324 6632 4328 6688
rect 4264 6628 4328 6632
rect 4344 6688 4408 6692
rect 4344 6632 4348 6688
rect 4348 6632 4404 6688
rect 4404 6632 4408 6688
rect 4344 6628 4408 6632
rect 4424 6688 4488 6692
rect 4424 6632 4428 6688
rect 4428 6632 4484 6688
rect 4484 6632 4488 6688
rect 4424 6628 4488 6632
rect 4504 6688 4568 6692
rect 4504 6632 4508 6688
rect 4508 6632 4564 6688
rect 4564 6632 4568 6688
rect 4504 6628 4568 6632
rect 34984 6688 35048 6692
rect 34984 6632 34988 6688
rect 34988 6632 35044 6688
rect 35044 6632 35048 6688
rect 34984 6628 35048 6632
rect 35064 6688 35128 6692
rect 35064 6632 35068 6688
rect 35068 6632 35124 6688
rect 35124 6632 35128 6688
rect 35064 6628 35128 6632
rect 35144 6688 35208 6692
rect 35144 6632 35148 6688
rect 35148 6632 35204 6688
rect 35204 6632 35208 6688
rect 35144 6628 35208 6632
rect 35224 6688 35288 6692
rect 35224 6632 35228 6688
rect 35228 6632 35284 6688
rect 35284 6632 35288 6688
rect 35224 6628 35288 6632
rect 19624 6022 19688 6026
rect 19624 5966 19628 6022
rect 19628 5966 19684 6022
rect 19684 5966 19688 6022
rect 19624 5962 19688 5966
rect 19704 6022 19768 6026
rect 19704 5966 19708 6022
rect 19708 5966 19764 6022
rect 19764 5966 19768 6022
rect 19704 5962 19768 5966
rect 19784 6022 19848 6026
rect 19784 5966 19788 6022
rect 19788 5966 19844 6022
rect 19844 5966 19848 6022
rect 19784 5962 19848 5966
rect 19864 6022 19928 6026
rect 19864 5966 19868 6022
rect 19868 5966 19924 6022
rect 19924 5966 19928 6022
rect 19864 5962 19928 5966
rect 50344 6022 50408 6026
rect 50344 5966 50348 6022
rect 50348 5966 50404 6022
rect 50404 5966 50408 6022
rect 50344 5962 50408 5966
rect 50424 6022 50488 6026
rect 50424 5966 50428 6022
rect 50428 5966 50484 6022
rect 50484 5966 50488 6022
rect 50424 5962 50488 5966
rect 50504 6022 50568 6026
rect 50504 5966 50508 6022
rect 50508 5966 50564 6022
rect 50564 5966 50568 6022
rect 50504 5962 50568 5966
rect 50584 6022 50648 6026
rect 50584 5966 50588 6022
rect 50588 5966 50644 6022
rect 50644 5966 50648 6022
rect 50584 5962 50648 5966
rect 4264 5356 4328 5360
rect 4264 5300 4268 5356
rect 4268 5300 4324 5356
rect 4324 5300 4328 5356
rect 4264 5296 4328 5300
rect 4344 5356 4408 5360
rect 4344 5300 4348 5356
rect 4348 5300 4404 5356
rect 4404 5300 4408 5356
rect 4344 5296 4408 5300
rect 4424 5356 4488 5360
rect 4424 5300 4428 5356
rect 4428 5300 4484 5356
rect 4484 5300 4488 5356
rect 4424 5296 4488 5300
rect 4504 5356 4568 5360
rect 4504 5300 4508 5356
rect 4508 5300 4564 5356
rect 4564 5300 4568 5356
rect 4504 5296 4568 5300
rect 34984 5356 35048 5360
rect 34984 5300 34988 5356
rect 34988 5300 35044 5356
rect 35044 5300 35048 5356
rect 34984 5296 35048 5300
rect 35064 5356 35128 5360
rect 35064 5300 35068 5356
rect 35068 5300 35124 5356
rect 35124 5300 35128 5356
rect 35064 5296 35128 5300
rect 35144 5356 35208 5360
rect 35144 5300 35148 5356
rect 35148 5300 35204 5356
rect 35204 5300 35208 5356
rect 35144 5296 35208 5300
rect 35224 5356 35288 5360
rect 35224 5300 35228 5356
rect 35228 5300 35284 5356
rect 35284 5300 35288 5356
rect 35224 5296 35288 5300
rect 19624 4690 19688 4694
rect 19624 4634 19628 4690
rect 19628 4634 19684 4690
rect 19684 4634 19688 4690
rect 19624 4630 19688 4634
rect 19704 4690 19768 4694
rect 19704 4634 19708 4690
rect 19708 4634 19764 4690
rect 19764 4634 19768 4690
rect 19704 4630 19768 4634
rect 19784 4690 19848 4694
rect 19784 4634 19788 4690
rect 19788 4634 19844 4690
rect 19844 4634 19848 4690
rect 19784 4630 19848 4634
rect 19864 4690 19928 4694
rect 19864 4634 19868 4690
rect 19868 4634 19924 4690
rect 19924 4634 19928 4690
rect 19864 4630 19928 4634
rect 50344 4690 50408 4694
rect 50344 4634 50348 4690
rect 50348 4634 50404 4690
rect 50404 4634 50408 4690
rect 50344 4630 50408 4634
rect 50424 4690 50488 4694
rect 50424 4634 50428 4690
rect 50428 4634 50484 4690
rect 50484 4634 50488 4690
rect 50424 4630 50488 4634
rect 50504 4690 50568 4694
rect 50504 4634 50508 4690
rect 50508 4634 50564 4690
rect 50564 4634 50568 4690
rect 50504 4630 50568 4634
rect 50584 4690 50648 4694
rect 50584 4634 50588 4690
rect 50588 4634 50644 4690
rect 50644 4634 50648 4690
rect 50584 4630 50648 4634
rect 4264 4024 4328 4028
rect 4264 3968 4268 4024
rect 4268 3968 4324 4024
rect 4324 3968 4328 4024
rect 4264 3964 4328 3968
rect 4344 4024 4408 4028
rect 4344 3968 4348 4024
rect 4348 3968 4404 4024
rect 4404 3968 4408 4024
rect 4344 3964 4408 3968
rect 4424 4024 4488 4028
rect 4424 3968 4428 4024
rect 4428 3968 4484 4024
rect 4484 3968 4488 4024
rect 4424 3964 4488 3968
rect 4504 4024 4568 4028
rect 4504 3968 4508 4024
rect 4508 3968 4564 4024
rect 4564 3968 4568 4024
rect 4504 3964 4568 3968
rect 34984 4024 35048 4028
rect 34984 3968 34988 4024
rect 34988 3968 35044 4024
rect 35044 3968 35048 4024
rect 34984 3964 35048 3968
rect 35064 4024 35128 4028
rect 35064 3968 35068 4024
rect 35068 3968 35124 4024
rect 35124 3968 35128 4024
rect 35064 3964 35128 3968
rect 35144 4024 35208 4028
rect 35144 3968 35148 4024
rect 35148 3968 35204 4024
rect 35204 3968 35208 4024
rect 35144 3964 35208 3968
rect 35224 4024 35288 4028
rect 35224 3968 35228 4024
rect 35228 3968 35284 4024
rect 35284 3968 35288 4024
rect 35224 3964 35288 3968
rect 19624 3358 19688 3362
rect 19624 3302 19628 3358
rect 19628 3302 19684 3358
rect 19684 3302 19688 3358
rect 19624 3298 19688 3302
rect 19704 3358 19768 3362
rect 19704 3302 19708 3358
rect 19708 3302 19764 3358
rect 19764 3302 19768 3358
rect 19704 3298 19768 3302
rect 19784 3358 19848 3362
rect 19784 3302 19788 3358
rect 19788 3302 19844 3358
rect 19844 3302 19848 3358
rect 19784 3298 19848 3302
rect 19864 3358 19928 3362
rect 19864 3302 19868 3358
rect 19868 3302 19924 3358
rect 19924 3302 19928 3358
rect 19864 3298 19928 3302
rect 50344 3358 50408 3362
rect 50344 3302 50348 3358
rect 50348 3302 50404 3358
rect 50404 3302 50408 3358
rect 50344 3298 50408 3302
rect 50424 3358 50488 3362
rect 50424 3302 50428 3358
rect 50428 3302 50484 3358
rect 50484 3302 50488 3358
rect 50424 3298 50488 3302
rect 50504 3358 50568 3362
rect 50504 3302 50508 3358
rect 50508 3302 50564 3358
rect 50564 3302 50568 3358
rect 50504 3298 50568 3302
rect 50584 3358 50648 3362
rect 50584 3302 50588 3358
rect 50588 3302 50644 3358
rect 50644 3302 50648 3358
rect 50584 3298 50648 3302
rect 4264 2692 4328 2696
rect 4264 2636 4268 2692
rect 4268 2636 4324 2692
rect 4324 2636 4328 2692
rect 4264 2632 4328 2636
rect 4344 2692 4408 2696
rect 4344 2636 4348 2692
rect 4348 2636 4404 2692
rect 4404 2636 4408 2692
rect 4344 2632 4408 2636
rect 4424 2692 4488 2696
rect 4424 2636 4428 2692
rect 4428 2636 4484 2692
rect 4484 2636 4488 2692
rect 4424 2632 4488 2636
rect 4504 2692 4568 2696
rect 4504 2636 4508 2692
rect 4508 2636 4564 2692
rect 4564 2636 4568 2692
rect 4504 2632 4568 2636
rect 34984 2692 35048 2696
rect 34984 2636 34988 2692
rect 34988 2636 35044 2692
rect 35044 2636 35048 2692
rect 34984 2632 35048 2636
rect 35064 2692 35128 2696
rect 35064 2636 35068 2692
rect 35068 2636 35124 2692
rect 35124 2636 35128 2692
rect 35064 2632 35128 2636
rect 35144 2692 35208 2696
rect 35144 2636 35148 2692
rect 35148 2636 35204 2692
rect 35204 2636 35208 2692
rect 35144 2632 35208 2636
rect 35224 2692 35288 2696
rect 35224 2636 35228 2692
rect 35228 2636 35284 2692
rect 35284 2636 35288 2692
rect 35224 2632 35288 2636
<< metal4 >>
rect 4256 57308 4576 57324
rect 4256 57244 4264 57308
rect 4328 57244 4344 57308
rect 4408 57244 4424 57308
rect 4488 57244 4504 57308
rect 4568 57244 4576 57308
rect 4256 55976 4576 57244
rect 4256 55912 4264 55976
rect 4328 55912 4344 55976
rect 4408 55912 4424 55976
rect 4488 55912 4504 55976
rect 4568 55912 4576 55976
rect 4256 54644 4576 55912
rect 4256 54580 4264 54644
rect 4328 54580 4344 54644
rect 4408 54580 4424 54644
rect 4488 54580 4504 54644
rect 4568 54580 4576 54644
rect 4256 53312 4576 54580
rect 4256 53248 4264 53312
rect 4328 53248 4344 53312
rect 4408 53248 4424 53312
rect 4488 53248 4504 53312
rect 4568 53248 4576 53312
rect 4256 51980 4576 53248
rect 4256 51916 4264 51980
rect 4328 51916 4344 51980
rect 4408 51916 4424 51980
rect 4488 51916 4504 51980
rect 4568 51916 4576 51980
rect 4256 50648 4576 51916
rect 4256 50584 4264 50648
rect 4328 50584 4344 50648
rect 4408 50584 4424 50648
rect 4488 50584 4504 50648
rect 4568 50584 4576 50648
rect 4256 49316 4576 50584
rect 4256 49252 4264 49316
rect 4328 49252 4344 49316
rect 4408 49252 4424 49316
rect 4488 49252 4504 49316
rect 4568 49252 4576 49316
rect 4256 47984 4576 49252
rect 4256 47920 4264 47984
rect 4328 47920 4344 47984
rect 4408 47920 4424 47984
rect 4488 47920 4504 47984
rect 4568 47920 4576 47984
rect 4256 46652 4576 47920
rect 4256 46588 4264 46652
rect 4328 46588 4344 46652
rect 4408 46588 4424 46652
rect 4488 46588 4504 46652
rect 4568 46588 4576 46652
rect 4256 45320 4576 46588
rect 4256 45256 4264 45320
rect 4328 45256 4344 45320
rect 4408 45256 4424 45320
rect 4488 45256 4504 45320
rect 4568 45256 4576 45320
rect 4256 43988 4576 45256
rect 4256 43924 4264 43988
rect 4328 43924 4344 43988
rect 4408 43924 4424 43988
rect 4488 43924 4504 43988
rect 4568 43924 4576 43988
rect 4256 42656 4576 43924
rect 4256 42592 4264 42656
rect 4328 42592 4344 42656
rect 4408 42592 4424 42656
rect 4488 42592 4504 42656
rect 4568 42592 4576 42656
rect 4256 41324 4576 42592
rect 4256 41260 4264 41324
rect 4328 41260 4344 41324
rect 4408 41260 4424 41324
rect 4488 41260 4504 41324
rect 4568 41260 4576 41324
rect 4256 39992 4576 41260
rect 4256 39928 4264 39992
rect 4328 39928 4344 39992
rect 4408 39928 4424 39992
rect 4488 39928 4504 39992
rect 4568 39928 4576 39992
rect 4256 38660 4576 39928
rect 4256 38596 4264 38660
rect 4328 38596 4344 38660
rect 4408 38596 4424 38660
rect 4488 38596 4504 38660
rect 4568 38596 4576 38660
rect 4256 37328 4576 38596
rect 4256 37264 4264 37328
rect 4328 37264 4344 37328
rect 4408 37264 4424 37328
rect 4488 37264 4504 37328
rect 4568 37264 4576 37328
rect 4256 35996 4576 37264
rect 4256 35932 4264 35996
rect 4328 35932 4344 35996
rect 4408 35932 4424 35996
rect 4488 35932 4504 35996
rect 4568 35932 4576 35996
rect 4256 34664 4576 35932
rect 4256 34600 4264 34664
rect 4328 34600 4344 34664
rect 4408 34600 4424 34664
rect 4488 34600 4504 34664
rect 4568 34600 4576 34664
rect 4256 33332 4576 34600
rect 4256 33268 4264 33332
rect 4328 33268 4344 33332
rect 4408 33268 4424 33332
rect 4488 33268 4504 33332
rect 4568 33268 4576 33332
rect 4256 32000 4576 33268
rect 4256 31936 4264 32000
rect 4328 31936 4344 32000
rect 4408 31936 4424 32000
rect 4488 31936 4504 32000
rect 4568 31936 4576 32000
rect 4256 30668 4576 31936
rect 4256 30604 4264 30668
rect 4328 30604 4344 30668
rect 4408 30604 4424 30668
rect 4488 30604 4504 30668
rect 4568 30604 4576 30668
rect 4256 29336 4576 30604
rect 4256 29272 4264 29336
rect 4328 29272 4344 29336
rect 4408 29272 4424 29336
rect 4488 29272 4504 29336
rect 4568 29272 4576 29336
rect 4256 28004 4576 29272
rect 4256 27940 4264 28004
rect 4328 27940 4344 28004
rect 4408 27940 4424 28004
rect 4488 27940 4504 28004
rect 4568 27940 4576 28004
rect 4256 26672 4576 27940
rect 4256 26608 4264 26672
rect 4328 26608 4344 26672
rect 4408 26608 4424 26672
rect 4488 26608 4504 26672
rect 4568 26608 4576 26672
rect 4256 25340 4576 26608
rect 4256 25276 4264 25340
rect 4328 25276 4344 25340
rect 4408 25276 4424 25340
rect 4488 25276 4504 25340
rect 4568 25276 4576 25340
rect 4256 24008 4576 25276
rect 4256 23944 4264 24008
rect 4328 23944 4344 24008
rect 4408 23944 4424 24008
rect 4488 23944 4504 24008
rect 4568 23944 4576 24008
rect 4256 22676 4576 23944
rect 4256 22612 4264 22676
rect 4328 22612 4344 22676
rect 4408 22612 4424 22676
rect 4488 22612 4504 22676
rect 4568 22612 4576 22676
rect 4256 21344 4576 22612
rect 4256 21280 4264 21344
rect 4328 21280 4344 21344
rect 4408 21280 4424 21344
rect 4488 21280 4504 21344
rect 4568 21280 4576 21344
rect 4256 20012 4576 21280
rect 4256 19948 4264 20012
rect 4328 19948 4344 20012
rect 4408 19948 4424 20012
rect 4488 19948 4504 20012
rect 4568 19948 4576 20012
rect 4256 18680 4576 19948
rect 4256 18616 4264 18680
rect 4328 18616 4344 18680
rect 4408 18616 4424 18680
rect 4488 18616 4504 18680
rect 4568 18616 4576 18680
rect 4256 17348 4576 18616
rect 4256 17284 4264 17348
rect 4328 17284 4344 17348
rect 4408 17284 4424 17348
rect 4488 17284 4504 17348
rect 4568 17284 4576 17348
rect 4256 16016 4576 17284
rect 4256 15952 4264 16016
rect 4328 15952 4344 16016
rect 4408 15952 4424 16016
rect 4488 15952 4504 16016
rect 4568 15952 4576 16016
rect 4256 14684 4576 15952
rect 4256 14620 4264 14684
rect 4328 14620 4344 14684
rect 4408 14620 4424 14684
rect 4488 14620 4504 14684
rect 4568 14620 4576 14684
rect 4256 13352 4576 14620
rect 4256 13288 4264 13352
rect 4328 13288 4344 13352
rect 4408 13288 4424 13352
rect 4488 13288 4504 13352
rect 4568 13288 4576 13352
rect 4256 12020 4576 13288
rect 4256 11956 4264 12020
rect 4328 11956 4344 12020
rect 4408 11956 4424 12020
rect 4488 11956 4504 12020
rect 4568 11956 4576 12020
rect 4256 10688 4576 11956
rect 4256 10624 4264 10688
rect 4328 10624 4344 10688
rect 4408 10624 4424 10688
rect 4488 10624 4504 10688
rect 4568 10624 4576 10688
rect 4256 9356 4576 10624
rect 4256 9292 4264 9356
rect 4328 9292 4344 9356
rect 4408 9292 4424 9356
rect 4488 9292 4504 9356
rect 4568 9292 4576 9356
rect 4256 8024 4576 9292
rect 4256 7960 4264 8024
rect 4328 7960 4344 8024
rect 4408 7960 4424 8024
rect 4488 7960 4504 8024
rect 4568 7960 4576 8024
rect 4256 6692 4576 7960
rect 4256 6628 4264 6692
rect 4328 6628 4344 6692
rect 4408 6628 4424 6692
rect 4488 6628 4504 6692
rect 4568 6628 4576 6692
rect 4256 5360 4576 6628
rect 4256 5296 4264 5360
rect 4328 5296 4344 5360
rect 4408 5296 4424 5360
rect 4488 5296 4504 5360
rect 4568 5296 4576 5360
rect 4256 4028 4576 5296
rect 4256 3964 4264 4028
rect 4328 3964 4344 4028
rect 4408 3964 4424 4028
rect 4488 3964 4504 4028
rect 4568 3964 4576 4028
rect 4256 2696 4576 3964
rect 4256 2632 4264 2696
rect 4328 2632 4344 2696
rect 4408 2632 4424 2696
rect 4488 2632 4504 2696
rect 4568 2632 4576 2696
rect 4916 2664 5236 57276
rect 5576 2664 5896 57276
rect 6236 2664 6556 57276
rect 19616 56642 19936 57324
rect 34976 57308 35296 57324
rect 19616 56578 19624 56642
rect 19688 56578 19704 56642
rect 19768 56578 19784 56642
rect 19848 56578 19864 56642
rect 19928 56578 19936 56642
rect 19616 55310 19936 56578
rect 19616 55246 19624 55310
rect 19688 55246 19704 55310
rect 19768 55246 19784 55310
rect 19848 55246 19864 55310
rect 19928 55246 19936 55310
rect 19616 53978 19936 55246
rect 19616 53914 19624 53978
rect 19688 53914 19704 53978
rect 19768 53914 19784 53978
rect 19848 53914 19864 53978
rect 19928 53914 19936 53978
rect 19616 52646 19936 53914
rect 19616 52582 19624 52646
rect 19688 52582 19704 52646
rect 19768 52582 19784 52646
rect 19848 52582 19864 52646
rect 19928 52582 19936 52646
rect 19616 51314 19936 52582
rect 19616 51250 19624 51314
rect 19688 51250 19704 51314
rect 19768 51250 19784 51314
rect 19848 51250 19864 51314
rect 19928 51250 19936 51314
rect 19616 49982 19936 51250
rect 19616 49918 19624 49982
rect 19688 49918 19704 49982
rect 19768 49918 19784 49982
rect 19848 49918 19864 49982
rect 19928 49918 19936 49982
rect 19616 48650 19936 49918
rect 19616 48586 19624 48650
rect 19688 48586 19704 48650
rect 19768 48586 19784 48650
rect 19848 48586 19864 48650
rect 19928 48586 19936 48650
rect 19616 47318 19936 48586
rect 19616 47254 19624 47318
rect 19688 47254 19704 47318
rect 19768 47254 19784 47318
rect 19848 47254 19864 47318
rect 19928 47254 19936 47318
rect 19616 45986 19936 47254
rect 19616 45922 19624 45986
rect 19688 45922 19704 45986
rect 19768 45922 19784 45986
rect 19848 45922 19864 45986
rect 19928 45922 19936 45986
rect 19616 44654 19936 45922
rect 19616 44590 19624 44654
rect 19688 44590 19704 44654
rect 19768 44590 19784 44654
rect 19848 44590 19864 44654
rect 19928 44590 19936 44654
rect 19616 43322 19936 44590
rect 19616 43258 19624 43322
rect 19688 43258 19704 43322
rect 19768 43258 19784 43322
rect 19848 43258 19864 43322
rect 19928 43258 19936 43322
rect 19616 41990 19936 43258
rect 19616 41926 19624 41990
rect 19688 41926 19704 41990
rect 19768 41926 19784 41990
rect 19848 41926 19864 41990
rect 19928 41926 19936 41990
rect 19616 40658 19936 41926
rect 19616 40594 19624 40658
rect 19688 40594 19704 40658
rect 19768 40594 19784 40658
rect 19848 40594 19864 40658
rect 19928 40594 19936 40658
rect 19616 39326 19936 40594
rect 19616 39262 19624 39326
rect 19688 39262 19704 39326
rect 19768 39262 19784 39326
rect 19848 39262 19864 39326
rect 19928 39262 19936 39326
rect 19616 37994 19936 39262
rect 19616 37930 19624 37994
rect 19688 37930 19704 37994
rect 19768 37930 19784 37994
rect 19848 37930 19864 37994
rect 19928 37930 19936 37994
rect 19616 36662 19936 37930
rect 19616 36598 19624 36662
rect 19688 36598 19704 36662
rect 19768 36598 19784 36662
rect 19848 36598 19864 36662
rect 19928 36598 19936 36662
rect 19616 35330 19936 36598
rect 19616 35266 19624 35330
rect 19688 35266 19704 35330
rect 19768 35266 19784 35330
rect 19848 35266 19864 35330
rect 19928 35266 19936 35330
rect 19616 33998 19936 35266
rect 19616 33934 19624 33998
rect 19688 33934 19704 33998
rect 19768 33934 19784 33998
rect 19848 33934 19864 33998
rect 19928 33934 19936 33998
rect 19616 32666 19936 33934
rect 19616 32602 19624 32666
rect 19688 32602 19704 32666
rect 19768 32602 19784 32666
rect 19848 32602 19864 32666
rect 19928 32602 19936 32666
rect 19616 31334 19936 32602
rect 19616 31270 19624 31334
rect 19688 31270 19704 31334
rect 19768 31270 19784 31334
rect 19848 31270 19864 31334
rect 19928 31270 19936 31334
rect 19616 30002 19936 31270
rect 19616 29938 19624 30002
rect 19688 29938 19704 30002
rect 19768 29938 19784 30002
rect 19848 29938 19864 30002
rect 19928 29938 19936 30002
rect 19616 28670 19936 29938
rect 19616 28606 19624 28670
rect 19688 28606 19704 28670
rect 19768 28606 19784 28670
rect 19848 28606 19864 28670
rect 19928 28606 19936 28670
rect 19616 27338 19936 28606
rect 19616 27274 19624 27338
rect 19688 27274 19704 27338
rect 19768 27274 19784 27338
rect 19848 27274 19864 27338
rect 19928 27274 19936 27338
rect 19616 26006 19936 27274
rect 19616 25942 19624 26006
rect 19688 25942 19704 26006
rect 19768 25942 19784 26006
rect 19848 25942 19864 26006
rect 19928 25942 19936 26006
rect 19616 24674 19936 25942
rect 19616 24610 19624 24674
rect 19688 24610 19704 24674
rect 19768 24610 19784 24674
rect 19848 24610 19864 24674
rect 19928 24610 19936 24674
rect 19616 23342 19936 24610
rect 19616 23278 19624 23342
rect 19688 23278 19704 23342
rect 19768 23278 19784 23342
rect 19848 23278 19864 23342
rect 19928 23278 19936 23342
rect 19616 22010 19936 23278
rect 19616 21946 19624 22010
rect 19688 21946 19704 22010
rect 19768 21946 19784 22010
rect 19848 21946 19864 22010
rect 19928 21946 19936 22010
rect 19616 20678 19936 21946
rect 19616 20614 19624 20678
rect 19688 20614 19704 20678
rect 19768 20614 19784 20678
rect 19848 20614 19864 20678
rect 19928 20614 19936 20678
rect 19616 19346 19936 20614
rect 19616 19282 19624 19346
rect 19688 19282 19704 19346
rect 19768 19282 19784 19346
rect 19848 19282 19864 19346
rect 19928 19282 19936 19346
rect 19616 18014 19936 19282
rect 19616 17950 19624 18014
rect 19688 17950 19704 18014
rect 19768 17950 19784 18014
rect 19848 17950 19864 18014
rect 19928 17950 19936 18014
rect 19616 16682 19936 17950
rect 19616 16618 19624 16682
rect 19688 16618 19704 16682
rect 19768 16618 19784 16682
rect 19848 16618 19864 16682
rect 19928 16618 19936 16682
rect 19616 15350 19936 16618
rect 19616 15286 19624 15350
rect 19688 15286 19704 15350
rect 19768 15286 19784 15350
rect 19848 15286 19864 15350
rect 19928 15286 19936 15350
rect 19616 14018 19936 15286
rect 19616 13954 19624 14018
rect 19688 13954 19704 14018
rect 19768 13954 19784 14018
rect 19848 13954 19864 14018
rect 19928 13954 19936 14018
rect 19616 12686 19936 13954
rect 19616 12622 19624 12686
rect 19688 12622 19704 12686
rect 19768 12622 19784 12686
rect 19848 12622 19864 12686
rect 19928 12622 19936 12686
rect 19616 11354 19936 12622
rect 19616 11290 19624 11354
rect 19688 11290 19704 11354
rect 19768 11290 19784 11354
rect 19848 11290 19864 11354
rect 19928 11290 19936 11354
rect 19616 10022 19936 11290
rect 19616 9958 19624 10022
rect 19688 9958 19704 10022
rect 19768 9958 19784 10022
rect 19848 9958 19864 10022
rect 19928 9958 19936 10022
rect 19616 8690 19936 9958
rect 19616 8626 19624 8690
rect 19688 8626 19704 8690
rect 19768 8626 19784 8690
rect 19848 8626 19864 8690
rect 19928 8626 19936 8690
rect 19616 7358 19936 8626
rect 19616 7294 19624 7358
rect 19688 7294 19704 7358
rect 19768 7294 19784 7358
rect 19848 7294 19864 7358
rect 19928 7294 19936 7358
rect 19616 6026 19936 7294
rect 19616 5962 19624 6026
rect 19688 5962 19704 6026
rect 19768 5962 19784 6026
rect 19848 5962 19864 6026
rect 19928 5962 19936 6026
rect 19616 4694 19936 5962
rect 19616 4630 19624 4694
rect 19688 4630 19704 4694
rect 19768 4630 19784 4694
rect 19848 4630 19864 4694
rect 19928 4630 19936 4694
rect 19616 3362 19936 4630
rect 19616 3298 19624 3362
rect 19688 3298 19704 3362
rect 19768 3298 19784 3362
rect 19848 3298 19864 3362
rect 19928 3298 19936 3362
rect 4256 2616 4576 2632
rect 19616 2616 19936 3298
rect 20276 2664 20596 57276
rect 20936 2664 21256 57276
rect 21596 2664 21916 57276
rect 34976 57244 34984 57308
rect 35048 57244 35064 57308
rect 35128 57244 35144 57308
rect 35208 57244 35224 57308
rect 35288 57244 35296 57308
rect 34976 55976 35296 57244
rect 34976 55912 34984 55976
rect 35048 55912 35064 55976
rect 35128 55912 35144 55976
rect 35208 55912 35224 55976
rect 35288 55912 35296 55976
rect 34976 54644 35296 55912
rect 34976 54580 34984 54644
rect 35048 54580 35064 54644
rect 35128 54580 35144 54644
rect 35208 54580 35224 54644
rect 35288 54580 35296 54644
rect 34976 53312 35296 54580
rect 34976 53248 34984 53312
rect 35048 53248 35064 53312
rect 35128 53248 35144 53312
rect 35208 53248 35224 53312
rect 35288 53248 35296 53312
rect 34976 51980 35296 53248
rect 34976 51916 34984 51980
rect 35048 51916 35064 51980
rect 35128 51916 35144 51980
rect 35208 51916 35224 51980
rect 35288 51916 35296 51980
rect 34976 50648 35296 51916
rect 34976 50584 34984 50648
rect 35048 50584 35064 50648
rect 35128 50584 35144 50648
rect 35208 50584 35224 50648
rect 35288 50584 35296 50648
rect 34976 49316 35296 50584
rect 34976 49252 34984 49316
rect 35048 49252 35064 49316
rect 35128 49252 35144 49316
rect 35208 49252 35224 49316
rect 35288 49252 35296 49316
rect 34976 47984 35296 49252
rect 34976 47920 34984 47984
rect 35048 47920 35064 47984
rect 35128 47920 35144 47984
rect 35208 47920 35224 47984
rect 35288 47920 35296 47984
rect 34976 46652 35296 47920
rect 34976 46588 34984 46652
rect 35048 46588 35064 46652
rect 35128 46588 35144 46652
rect 35208 46588 35224 46652
rect 35288 46588 35296 46652
rect 34976 45320 35296 46588
rect 34976 45256 34984 45320
rect 35048 45256 35064 45320
rect 35128 45256 35144 45320
rect 35208 45256 35224 45320
rect 35288 45256 35296 45320
rect 34976 43988 35296 45256
rect 34976 43924 34984 43988
rect 35048 43924 35064 43988
rect 35128 43924 35144 43988
rect 35208 43924 35224 43988
rect 35288 43924 35296 43988
rect 34976 42656 35296 43924
rect 34976 42592 34984 42656
rect 35048 42592 35064 42656
rect 35128 42592 35144 42656
rect 35208 42592 35224 42656
rect 35288 42592 35296 42656
rect 34976 41324 35296 42592
rect 34976 41260 34984 41324
rect 35048 41260 35064 41324
rect 35128 41260 35144 41324
rect 35208 41260 35224 41324
rect 35288 41260 35296 41324
rect 34976 39992 35296 41260
rect 34976 39928 34984 39992
rect 35048 39928 35064 39992
rect 35128 39928 35144 39992
rect 35208 39928 35224 39992
rect 35288 39928 35296 39992
rect 34976 38660 35296 39928
rect 34976 38596 34984 38660
rect 35048 38596 35064 38660
rect 35128 38596 35144 38660
rect 35208 38596 35224 38660
rect 35288 38596 35296 38660
rect 34976 37328 35296 38596
rect 34976 37264 34984 37328
rect 35048 37264 35064 37328
rect 35128 37264 35144 37328
rect 35208 37264 35224 37328
rect 35288 37264 35296 37328
rect 34976 35996 35296 37264
rect 34976 35932 34984 35996
rect 35048 35932 35064 35996
rect 35128 35932 35144 35996
rect 35208 35932 35224 35996
rect 35288 35932 35296 35996
rect 34976 34664 35296 35932
rect 34976 34600 34984 34664
rect 35048 34600 35064 34664
rect 35128 34600 35144 34664
rect 35208 34600 35224 34664
rect 35288 34600 35296 34664
rect 34976 33332 35296 34600
rect 34976 33268 34984 33332
rect 35048 33268 35064 33332
rect 35128 33268 35144 33332
rect 35208 33268 35224 33332
rect 35288 33268 35296 33332
rect 34976 32000 35296 33268
rect 34976 31936 34984 32000
rect 35048 31936 35064 32000
rect 35128 31936 35144 32000
rect 35208 31936 35224 32000
rect 35288 31936 35296 32000
rect 34976 30668 35296 31936
rect 34976 30604 34984 30668
rect 35048 30604 35064 30668
rect 35128 30604 35144 30668
rect 35208 30604 35224 30668
rect 35288 30604 35296 30668
rect 34976 29336 35296 30604
rect 34976 29272 34984 29336
rect 35048 29272 35064 29336
rect 35128 29272 35144 29336
rect 35208 29272 35224 29336
rect 35288 29272 35296 29336
rect 34976 28004 35296 29272
rect 34976 27940 34984 28004
rect 35048 27940 35064 28004
rect 35128 27940 35144 28004
rect 35208 27940 35224 28004
rect 35288 27940 35296 28004
rect 34976 26672 35296 27940
rect 34976 26608 34984 26672
rect 35048 26608 35064 26672
rect 35128 26608 35144 26672
rect 35208 26608 35224 26672
rect 35288 26608 35296 26672
rect 34976 25340 35296 26608
rect 34976 25276 34984 25340
rect 35048 25276 35064 25340
rect 35128 25276 35144 25340
rect 35208 25276 35224 25340
rect 35288 25276 35296 25340
rect 34976 24008 35296 25276
rect 34976 23944 34984 24008
rect 35048 23944 35064 24008
rect 35128 23944 35144 24008
rect 35208 23944 35224 24008
rect 35288 23944 35296 24008
rect 34976 22676 35296 23944
rect 34976 22612 34984 22676
rect 35048 22612 35064 22676
rect 35128 22612 35144 22676
rect 35208 22612 35224 22676
rect 35288 22612 35296 22676
rect 34976 21344 35296 22612
rect 34976 21280 34984 21344
rect 35048 21280 35064 21344
rect 35128 21280 35144 21344
rect 35208 21280 35224 21344
rect 35288 21280 35296 21344
rect 34976 20012 35296 21280
rect 34976 19948 34984 20012
rect 35048 19948 35064 20012
rect 35128 19948 35144 20012
rect 35208 19948 35224 20012
rect 35288 19948 35296 20012
rect 34976 18680 35296 19948
rect 34976 18616 34984 18680
rect 35048 18616 35064 18680
rect 35128 18616 35144 18680
rect 35208 18616 35224 18680
rect 35288 18616 35296 18680
rect 34976 17348 35296 18616
rect 34976 17284 34984 17348
rect 35048 17284 35064 17348
rect 35128 17284 35144 17348
rect 35208 17284 35224 17348
rect 35288 17284 35296 17348
rect 34976 16016 35296 17284
rect 34976 15952 34984 16016
rect 35048 15952 35064 16016
rect 35128 15952 35144 16016
rect 35208 15952 35224 16016
rect 35288 15952 35296 16016
rect 34976 14684 35296 15952
rect 34976 14620 34984 14684
rect 35048 14620 35064 14684
rect 35128 14620 35144 14684
rect 35208 14620 35224 14684
rect 35288 14620 35296 14684
rect 34976 13352 35296 14620
rect 34976 13288 34984 13352
rect 35048 13288 35064 13352
rect 35128 13288 35144 13352
rect 35208 13288 35224 13352
rect 35288 13288 35296 13352
rect 34976 12020 35296 13288
rect 34976 11956 34984 12020
rect 35048 11956 35064 12020
rect 35128 11956 35144 12020
rect 35208 11956 35224 12020
rect 35288 11956 35296 12020
rect 34976 10688 35296 11956
rect 34976 10624 34984 10688
rect 35048 10624 35064 10688
rect 35128 10624 35144 10688
rect 35208 10624 35224 10688
rect 35288 10624 35296 10688
rect 34976 9356 35296 10624
rect 34976 9292 34984 9356
rect 35048 9292 35064 9356
rect 35128 9292 35144 9356
rect 35208 9292 35224 9356
rect 35288 9292 35296 9356
rect 34976 8024 35296 9292
rect 34976 7960 34984 8024
rect 35048 7960 35064 8024
rect 35128 7960 35144 8024
rect 35208 7960 35224 8024
rect 35288 7960 35296 8024
rect 34976 6692 35296 7960
rect 34976 6628 34984 6692
rect 35048 6628 35064 6692
rect 35128 6628 35144 6692
rect 35208 6628 35224 6692
rect 35288 6628 35296 6692
rect 34976 5360 35296 6628
rect 34976 5296 34984 5360
rect 35048 5296 35064 5360
rect 35128 5296 35144 5360
rect 35208 5296 35224 5360
rect 35288 5296 35296 5360
rect 34976 4028 35296 5296
rect 34976 3964 34984 4028
rect 35048 3964 35064 4028
rect 35128 3964 35144 4028
rect 35208 3964 35224 4028
rect 35288 3964 35296 4028
rect 34976 2696 35296 3964
rect 34976 2632 34984 2696
rect 35048 2632 35064 2696
rect 35128 2632 35144 2696
rect 35208 2632 35224 2696
rect 35288 2632 35296 2696
rect 35636 2664 35956 57276
rect 36296 2664 36616 57276
rect 36956 2664 37276 57276
rect 50336 56642 50656 57324
rect 50336 56578 50344 56642
rect 50408 56578 50424 56642
rect 50488 56578 50504 56642
rect 50568 56578 50584 56642
rect 50648 56578 50656 56642
rect 50336 55310 50656 56578
rect 50336 55246 50344 55310
rect 50408 55246 50424 55310
rect 50488 55246 50504 55310
rect 50568 55246 50584 55310
rect 50648 55246 50656 55310
rect 50336 53978 50656 55246
rect 50336 53914 50344 53978
rect 50408 53914 50424 53978
rect 50488 53914 50504 53978
rect 50568 53914 50584 53978
rect 50648 53914 50656 53978
rect 50336 52646 50656 53914
rect 50336 52582 50344 52646
rect 50408 52582 50424 52646
rect 50488 52582 50504 52646
rect 50568 52582 50584 52646
rect 50648 52582 50656 52646
rect 50336 51314 50656 52582
rect 50336 51250 50344 51314
rect 50408 51250 50424 51314
rect 50488 51250 50504 51314
rect 50568 51250 50584 51314
rect 50648 51250 50656 51314
rect 50336 49982 50656 51250
rect 50336 49918 50344 49982
rect 50408 49918 50424 49982
rect 50488 49918 50504 49982
rect 50568 49918 50584 49982
rect 50648 49918 50656 49982
rect 50336 48650 50656 49918
rect 50336 48586 50344 48650
rect 50408 48586 50424 48650
rect 50488 48586 50504 48650
rect 50568 48586 50584 48650
rect 50648 48586 50656 48650
rect 50336 47318 50656 48586
rect 50336 47254 50344 47318
rect 50408 47254 50424 47318
rect 50488 47254 50504 47318
rect 50568 47254 50584 47318
rect 50648 47254 50656 47318
rect 50336 45986 50656 47254
rect 50336 45922 50344 45986
rect 50408 45922 50424 45986
rect 50488 45922 50504 45986
rect 50568 45922 50584 45986
rect 50648 45922 50656 45986
rect 50336 44654 50656 45922
rect 50336 44590 50344 44654
rect 50408 44590 50424 44654
rect 50488 44590 50504 44654
rect 50568 44590 50584 44654
rect 50648 44590 50656 44654
rect 50336 43322 50656 44590
rect 50336 43258 50344 43322
rect 50408 43258 50424 43322
rect 50488 43258 50504 43322
rect 50568 43258 50584 43322
rect 50648 43258 50656 43322
rect 50336 41990 50656 43258
rect 50336 41926 50344 41990
rect 50408 41926 50424 41990
rect 50488 41926 50504 41990
rect 50568 41926 50584 41990
rect 50648 41926 50656 41990
rect 50336 40658 50656 41926
rect 50336 40594 50344 40658
rect 50408 40594 50424 40658
rect 50488 40594 50504 40658
rect 50568 40594 50584 40658
rect 50648 40594 50656 40658
rect 50336 39326 50656 40594
rect 50336 39262 50344 39326
rect 50408 39262 50424 39326
rect 50488 39262 50504 39326
rect 50568 39262 50584 39326
rect 50648 39262 50656 39326
rect 50336 37994 50656 39262
rect 50336 37930 50344 37994
rect 50408 37930 50424 37994
rect 50488 37930 50504 37994
rect 50568 37930 50584 37994
rect 50648 37930 50656 37994
rect 50336 36662 50656 37930
rect 50336 36598 50344 36662
rect 50408 36598 50424 36662
rect 50488 36598 50504 36662
rect 50568 36598 50584 36662
rect 50648 36598 50656 36662
rect 50336 35330 50656 36598
rect 50336 35266 50344 35330
rect 50408 35266 50424 35330
rect 50488 35266 50504 35330
rect 50568 35266 50584 35330
rect 50648 35266 50656 35330
rect 50336 33998 50656 35266
rect 50336 33934 50344 33998
rect 50408 33934 50424 33998
rect 50488 33934 50504 33998
rect 50568 33934 50584 33998
rect 50648 33934 50656 33998
rect 50336 32666 50656 33934
rect 50336 32602 50344 32666
rect 50408 32602 50424 32666
rect 50488 32602 50504 32666
rect 50568 32602 50584 32666
rect 50648 32602 50656 32666
rect 50336 31334 50656 32602
rect 50336 31270 50344 31334
rect 50408 31270 50424 31334
rect 50488 31270 50504 31334
rect 50568 31270 50584 31334
rect 50648 31270 50656 31334
rect 50336 30002 50656 31270
rect 50336 29938 50344 30002
rect 50408 29938 50424 30002
rect 50488 29938 50504 30002
rect 50568 29938 50584 30002
rect 50648 29938 50656 30002
rect 50336 28670 50656 29938
rect 50336 28606 50344 28670
rect 50408 28606 50424 28670
rect 50488 28606 50504 28670
rect 50568 28606 50584 28670
rect 50648 28606 50656 28670
rect 50336 27338 50656 28606
rect 50336 27274 50344 27338
rect 50408 27274 50424 27338
rect 50488 27274 50504 27338
rect 50568 27274 50584 27338
rect 50648 27274 50656 27338
rect 50336 26006 50656 27274
rect 50336 25942 50344 26006
rect 50408 25942 50424 26006
rect 50488 25942 50504 26006
rect 50568 25942 50584 26006
rect 50648 25942 50656 26006
rect 50336 24674 50656 25942
rect 50336 24610 50344 24674
rect 50408 24610 50424 24674
rect 50488 24610 50504 24674
rect 50568 24610 50584 24674
rect 50648 24610 50656 24674
rect 50336 23342 50656 24610
rect 50336 23278 50344 23342
rect 50408 23278 50424 23342
rect 50488 23278 50504 23342
rect 50568 23278 50584 23342
rect 50648 23278 50656 23342
rect 50336 22010 50656 23278
rect 50336 21946 50344 22010
rect 50408 21946 50424 22010
rect 50488 21946 50504 22010
rect 50568 21946 50584 22010
rect 50648 21946 50656 22010
rect 50336 20678 50656 21946
rect 50336 20614 50344 20678
rect 50408 20614 50424 20678
rect 50488 20614 50504 20678
rect 50568 20614 50584 20678
rect 50648 20614 50656 20678
rect 50336 19346 50656 20614
rect 50336 19282 50344 19346
rect 50408 19282 50424 19346
rect 50488 19282 50504 19346
rect 50568 19282 50584 19346
rect 50648 19282 50656 19346
rect 50336 18014 50656 19282
rect 50336 17950 50344 18014
rect 50408 17950 50424 18014
rect 50488 17950 50504 18014
rect 50568 17950 50584 18014
rect 50648 17950 50656 18014
rect 50336 16682 50656 17950
rect 50336 16618 50344 16682
rect 50408 16618 50424 16682
rect 50488 16618 50504 16682
rect 50568 16618 50584 16682
rect 50648 16618 50656 16682
rect 50336 15350 50656 16618
rect 50336 15286 50344 15350
rect 50408 15286 50424 15350
rect 50488 15286 50504 15350
rect 50568 15286 50584 15350
rect 50648 15286 50656 15350
rect 50336 14018 50656 15286
rect 50336 13954 50344 14018
rect 50408 13954 50424 14018
rect 50488 13954 50504 14018
rect 50568 13954 50584 14018
rect 50648 13954 50656 14018
rect 50336 12686 50656 13954
rect 50336 12622 50344 12686
rect 50408 12622 50424 12686
rect 50488 12622 50504 12686
rect 50568 12622 50584 12686
rect 50648 12622 50656 12686
rect 50336 11354 50656 12622
rect 50336 11290 50344 11354
rect 50408 11290 50424 11354
rect 50488 11290 50504 11354
rect 50568 11290 50584 11354
rect 50648 11290 50656 11354
rect 50336 10022 50656 11290
rect 50336 9958 50344 10022
rect 50408 9958 50424 10022
rect 50488 9958 50504 10022
rect 50568 9958 50584 10022
rect 50648 9958 50656 10022
rect 50336 8690 50656 9958
rect 50336 8626 50344 8690
rect 50408 8626 50424 8690
rect 50488 8626 50504 8690
rect 50568 8626 50584 8690
rect 50648 8626 50656 8690
rect 50336 7358 50656 8626
rect 50336 7294 50344 7358
rect 50408 7294 50424 7358
rect 50488 7294 50504 7358
rect 50568 7294 50584 7358
rect 50648 7294 50656 7358
rect 50336 6026 50656 7294
rect 50336 5962 50344 6026
rect 50408 5962 50424 6026
rect 50488 5962 50504 6026
rect 50568 5962 50584 6026
rect 50648 5962 50656 6026
rect 50336 4694 50656 5962
rect 50336 4630 50344 4694
rect 50408 4630 50424 4694
rect 50488 4630 50504 4694
rect 50568 4630 50584 4694
rect 50648 4630 50656 4694
rect 50336 3362 50656 4630
rect 50336 3298 50344 3362
rect 50408 3298 50424 3362
rect 50488 3298 50504 3362
rect 50568 3298 50584 3362
rect 50648 3298 50656 3362
rect 34976 2616 35296 2632
rect 50336 2616 50656 3298
rect 50996 2664 51316 57276
rect 51656 2664 51976 57276
rect 52316 2664 52636 57276
use sky130_fd_sc_ls__decap_4  FILLER_1_8 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1920 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_8
timestamp 1621261055
transform 1 0 1920 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input296 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input295
timestamp 1621261055
transform 1 0 1536 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_2
timestamp 1621261055
transform 1 0 1152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_0
timestamp 1621261055
transform 1 0 1152 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_16
timestamp 1621261055
transform 1 0 2688 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_16
timestamp 1621261055
transform 1 0 2688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input319
timestamp 1621261055
transform 1 0 2304 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input297
timestamp 1621261055
transform 1 0 2304 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_24
timestamp 1621261055
transform 1 0 3456 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_24
timestamp 1621261055
transform 1 0 3456 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input323
timestamp 1621261055
transform 1 0 3072 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input322
timestamp 1621261055
transform 1 0 3072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_32
timestamp 1621261055
transform 1 0 4224 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3936 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input324
timestamp 1621261055
transform 1 0 3840 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_164 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 3840 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 4704 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input325
timestamp 1621261055
transform 1 0 4608 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_40
timestamp 1621261055
transform 1 0 4992 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input298
timestamp 1621261055
transform 1 0 4896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_44
timestamp 1621261055
transform 1 0 5376 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_43
timestamp 1621261055
transform 1 0 5280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input300
timestamp 1621261055
transform 1 0 5568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input299
timestamp 1621261055
transform 1 0 5664 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_50
timestamp 1621261055
transform 1 0 5952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_51
timestamp 1621261055
transform 1 0 6048 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_56
timestamp 1621261055
transform 1 0 6528 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 6336 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_57
timestamp 1621261055
transform 1 0 6624 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_55
timestamp 1621261055
transform 1 0 6432 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_185
timestamp 1621261055
transform 1 0 6432 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_165
timestamp 1621261055
transform 1 0 6528 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input302
timestamp 1621261055
transform 1 0 6912 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input301
timestamp 1621261055
transform 1 0 7008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_64
timestamp 1621261055
transform 1 0 7296 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_65
timestamp 1621261055
transform 1 0 7392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input304
timestamp 1621261055
transform 1 0 7680 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input303
timestamp 1621261055
transform 1 0 7776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_72
timestamp 1621261055
transform 1 0 8064 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_73
timestamp 1621261055
transform 1 0 8160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_80
timestamp 1621261055
transform 1 0 8832 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_80
timestamp 1621261055
transform 1 0 8832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input306
timestamp 1621261055
transform 1 0 8448 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 8544 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_85
timestamp 1621261055
transform 1 0 9312 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input309
timestamp 1621261055
transform 1 0 9216 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_166
timestamp 1621261055
transform 1 0 9216 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_88
timestamp 1621261055
transform 1 0 9600 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input307
timestamp 1621261055
transform 1 0 9696 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_93
timestamp 1621261055
transform 1 0 10080 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input311
timestamp 1621261055
transform 1 0 9984 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_96
timestamp 1621261055
transform 1 0 10368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input310
timestamp 1621261055
transform 1 0 10464 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_104
timestamp 1621261055
transform 1 0 11136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_101
timestamp 1621261055
transform 1 0 10848 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input313
timestamp 1621261055
transform 1 0 10752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_1_111
timestamp 1621261055
transform 1 0 11808 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_108
timestamp 1621261055
transform 1 0 11520 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_113
timestamp 1621261055
transform 1 0 12000 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_0_111
timestamp 1621261055
transform 1 0 11808 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_109
timestamp 1621261055
transform 1 0 11616 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_186
timestamp 1621261055
transform 1 0 11712 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_167
timestamp 1621261055
transform 1 0 11904 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_1_121
timestamp 1621261055
transform 1 0 12768 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_119
timestamp 1621261055
transform 1 0 12576 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_121
timestamp 1621261055
transform 1 0 12768 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input167
timestamp 1621261055
transform 1 0 12864 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input39
timestamp 1621261055
transform 1 0 12960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_126
timestamp 1621261055
transform 1 0 13248 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_127
timestamp 1621261055
transform 1 0 13344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input89
timestamp 1621261055
transform 1 0 13632 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input78
timestamp 1621261055
transform 1 0 13728 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_134
timestamp 1621261055
transform 1 0 14016 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_135
timestamp 1621261055
transform 1 0 14112 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_141
timestamp 1621261055
transform 1 0 14688 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_139
timestamp 1621261055
transform 1 0 14496 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input100
timestamp 1621261055
transform 1 0 14400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_168
timestamp 1621261055
transform 1 0 14592 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_142
timestamp 1621261055
transform 1 0 14784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input122 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 15168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input111
timestamp 1621261055
transform 1 0 15072 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_150
timestamp 1621261055
transform 1 0 15552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_149
timestamp 1621261055
transform 1 0 15456 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_156
timestamp 1621261055
transform 1 0 16128 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input133
timestamp 1621261055
transform 1 0 15936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _066_
timestamp 1621261055
transform 1 0 15840 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_158
timestamp 1621261055
transform 1 0 16320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input50
timestamp 1621261055
transform 1 0 16512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_164
timestamp 1621261055
transform 1 0 16896 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_162
timestamp 1621261055
transform 1 0 16704 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_164
timestamp 1621261055
transform 1 0 16896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_187
timestamp 1621261055
transform 1 0 16992 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_166
timestamp 1621261055
transform 1 0 17088 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_169
timestamp 1621261055
transform 1 0 17376 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_169
timestamp 1621261055
transform 1 0 17280 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_174
timestamp 1621261055
transform 1 0 17856 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input70
timestamp 1621261055
transform 1 0 17472 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input61
timestamp 1621261055
transform 1 0 17760 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_177
timestamp 1621261055
transform 1 0 18144 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input72
timestamp 1621261055
transform 1 0 18240 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_182
timestamp 1621261055
transform 1 0 18624 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input71
timestamp 1621261055
transform 1 0 18528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_185
timestamp 1621261055
transform 1 0 18912 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_22 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform -1 0 19296 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input73
timestamp 1621261055
transform 1 0 19008 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _009_
timestamp 1621261055
transform -1 0 19584 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_190
timestamp 1621261055
transform 1 0 19392 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_192
timestamp 1621261055
transform 1 0 19584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_198
timestamp 1621261055
transform 1 0 20160 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_197
timestamp 1621261055
transform 1 0 20064 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input75
timestamp 1621261055
transform 1 0 19776 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_170
timestamp 1621261055
transform 1 0 19968 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_206
timestamp 1621261055
transform 1 0 20928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_205
timestamp 1621261055
transform 1 0 20832 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  input77 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 20544 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input74
timestamp 1621261055
transform 1 0 20448 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_214
timestamp 1621261055
transform 1 0 21696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_213
timestamp 1621261055
transform 1 0 21600 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input80
timestamp 1621261055
transform 1 0 21312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input76
timestamp 1621261055
transform 1 0 21216 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_221
timestamp 1621261055
transform 1 0 22368 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_218
timestamp 1621261055
transform 1 0 22080 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_0_223
timestamp 1621261055
transform 1 0 22560 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_221
timestamp 1621261055
transform 1 0 22368 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_188
timestamp 1621261055
transform 1 0 22272 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_171
timestamp 1621261055
transform 1 0 22656 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_229
timestamp 1621261055
transform 1 0 23136 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_225
timestamp 1621261055
transform 1 0 22752 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input84
timestamp 1621261055
transform 1 0 22752 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input82
timestamp 1621261055
transform 1 0 23136 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_237
timestamp 1621261055
transform 1 0 23904 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_233
timestamp 1621261055
transform 1 0 23520 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input86
timestamp 1621261055
transform 1 0 23520 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input85
timestamp 1621261055
transform 1 0 23904 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_245
timestamp 1621261055
transform 1 0 24672 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_241
timestamp 1621261055
transform 1 0 24288 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input88
timestamp 1621261055
transform 1 0 24288 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_253
timestamp 1621261055
transform 1 0 25440 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_253
timestamp 1621261055
transform 1 0 25440 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_251
timestamp 1621261055
transform 1 0 25248 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_249
timestamp 1621261055
transform 1 0 25056 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input92
timestamp 1621261055
transform 1 0 25824 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input91
timestamp 1621261055
transform 1 0 25056 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input90
timestamp 1621261055
transform 1 0 25824 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_172
timestamp 1621261055
transform 1 0 25344 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_261
timestamp 1621261055
transform 1 0 26208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_261
timestamp 1621261055
transform 1 0 26208 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_269
timestamp 1621261055
transform 1 0 26976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_269
timestamp 1621261055
transform 1 0 26976 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input95
timestamp 1621261055
transform 1 0 26592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input93
timestamp 1621261055
transform 1 0 26592 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_276
timestamp 1621261055
transform 1 0 27648 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_273
timestamp 1621261055
transform 1 0 27360 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_0_281
timestamp 1621261055
transform 1 0 28128 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_279
timestamp 1621261055
transform 1 0 27936 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_277
timestamp 1621261055
transform 1 0 27744 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input99
timestamp 1621261055
transform 1 0 28032 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_189
timestamp 1621261055
transform 1 0 27552 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_173
timestamp 1621261055
transform 1 0 28032 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_284
timestamp 1621261055
transform 1 0 28416 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_289
timestamp 1621261055
transform 1 0 28896 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input102
timestamp 1621261055
transform 1 0 28800 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input98
timestamp 1621261055
transform 1 0 28512 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_292
timestamp 1621261055
transform 1 0 29184 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_297
timestamp 1621261055
transform 1 0 29664 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input104
timestamp 1621261055
transform 1 0 29568 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input101
timestamp 1621261055
transform 1 0 29280 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_300
timestamp 1621261055
transform 1 0 29952 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_305
timestamp 1621261055
transform 1 0 30432 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input106
timestamp 1621261055
transform 1 0 30336 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_308
timestamp 1621261055
transform 1 0 30720 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_309
timestamp 1621261055
transform 1 0 30816 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_307
timestamp 1621261055
transform 1 0 30624 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_174
timestamp 1621261055
transform 1 0 30720 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_316
timestamp 1621261055
transform 1 0 31488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input108
timestamp 1621261055
transform 1 0 31104 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input107
timestamp 1621261055
transform 1 0 31200 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_317
timestamp 1621261055
transform 1 0 31584 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input112
timestamp 1621261055
transform 1 0 31872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input109
timestamp 1621261055
transform 1 0 31968 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_324
timestamp 1621261055
transform 1 0 32256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_325
timestamp 1621261055
transform 1 0 32352 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_328
timestamp 1621261055
transform 1 0 32640 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_190
timestamp 1621261055
transform 1 0 32832 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _197_
timestamp 1621261055
transform 1 0 32736 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_331
timestamp 1621261055
transform 1 0 32928 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_337
timestamp 1621261055
transform 1 0 33504 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_332
timestamp 1621261055
transform 1 0 33024 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input115
timestamp 1621261055
transform 1 0 33312 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_175
timestamp 1621261055
transform 1 0 33408 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_347
timestamp 1621261055
transform 1 0 34464 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_339
timestamp 1621261055
transform 1 0 33696 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_345
timestamp 1621261055
transform 1 0 34272 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input118
timestamp 1621261055
transform 1 0 34080 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input114
timestamp 1621261055
transform 1 0 33888 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_355
timestamp 1621261055
transform 1 0 35232 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_353
timestamp 1621261055
transform 1 0 35040 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input120
timestamp 1621261055
transform 1 0 34848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input117
timestamp 1621261055
transform 1 0 34656 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_363
timestamp 1621261055
transform 1 0 36000 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_363
timestamp 1621261055
transform 1 0 36000 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_361
timestamp 1621261055
transform 1 0 35808 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input123
timestamp 1621261055
transform 1 0 35616 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_371
timestamp 1621261055
transform 1 0 36768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_365
timestamp 1621261055
transform 1 0 36192 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input125
timestamp 1621261055
transform 1 0 36384 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input124
timestamp 1621261055
transform 1 0 36576 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_176
timestamp 1621261055
transform 1 0 36096 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_379
timestamp 1621261055
transform 1 0 37536 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_373
timestamp 1621261055
transform 1 0 36960 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input127
timestamp 1621261055
transform 1 0 37152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input126
timestamp 1621261055
transform 1 0 37344 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_386
timestamp 1621261055
transform 1 0 38208 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_383
timestamp 1621261055
transform 1 0 37920 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_389
timestamp 1621261055
transform 1 0 38496 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_0_381
timestamp 1621261055
transform 1 0 37728 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_191
timestamp 1621261055
transform 1 0 38112 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_394
timestamp 1621261055
transform 1 0 38976 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_393
timestamp 1621261055
transform 1 0 38880 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_391
timestamp 1621261055
transform 1 0 38688 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input131
timestamp 1621261055
transform 1 0 38592 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_177
timestamp 1621261055
transform 1 0 38784 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input134
timestamp 1621261055
transform 1 0 39360 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input130
timestamp 1621261055
transform 1 0 39264 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_402
timestamp 1621261055
transform 1 0 39744 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_401
timestamp 1621261055
transform 1 0 39648 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input132
timestamp 1621261055
transform 1 0 40032 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_410
timestamp 1621261055
transform 1 0 40512 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_409
timestamp 1621261055
transform 1 0 40416 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input136
timestamp 1621261055
transform 1 0 40128 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_83
timestamp 1621261055
transform 1 0 40608 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input138
timestamp 1621261055
transform 1 0 40896 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _058_
timestamp 1621261055
transform 1 0 40800 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_418
timestamp 1621261055
transform 1 0 41280 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_416
timestamp 1621261055
transform 1 0 41088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_178
timestamp 1621261055
transform 1 0 41472 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_421
timestamp 1621261055
transform 1 0 41568 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input140
timestamp 1621261055
transform 1 0 41664 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_426
timestamp 1621261055
transform 1 0 42048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_429
timestamp 1621261055
transform 1 0 42336 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input139
timestamp 1621261055
transform 1 0 41952 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input142
timestamp 1621261055
transform 1 0 42432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input141
timestamp 1621261055
transform 1 0 42720 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_438
timestamp 1621261055
transform 1 0 43200 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_434
timestamp 1621261055
transform 1 0 42816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_437
timestamp 1621261055
transform 1 0 43104 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_441
timestamp 1621261055
transform 1 0 43488 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_61
timestamp 1621261055
transform -1 0 43488 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_192
timestamp 1621261055
transform 1 0 43392 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _050_
timestamp 1621261055
transform -1 0 43776 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_0_444
timestamp 1621261055
transform 1 0 43776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input146
timestamp 1621261055
transform 1 0 43872 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_179
timestamp 1621261055
transform 1 0 44160 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_449
timestamp 1621261055
transform 1 0 44256 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_449
timestamp 1621261055
transform 1 0 44256 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input149
timestamp 1621261055
transform 1 0 44640 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input147
timestamp 1621261055
transform 1 0 44640 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_457
timestamp 1621261055
transform 1 0 45024 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_457
timestamp 1621261055
transform 1 0 45024 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input151
timestamp 1621261055
transform 1 0 45408 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input150
timestamp 1621261055
transform 1 0 45408 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_465
timestamp 1621261055
transform 1 0 45792 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_465
timestamp 1621261055
transform 1 0 45792 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input153
timestamp 1621261055
transform 1 0 46176 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_473
timestamp 1621261055
transform 1 0 46560 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_477
timestamp 1621261055
transform 1 0 46944 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_475
timestamp 1621261055
transform 1 0 46752 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_473
timestamp 1621261055
transform 1 0 46560 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input156
timestamp 1621261055
transform 1 0 46944 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_180
timestamp 1621261055
transform 1 0 46848 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_481
timestamp 1621261055
transform 1 0 47328 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_485
timestamp 1621261055
transform 1 0 47712 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input159
timestamp 1621261055
transform 1 0 47712 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input154
timestamp 1621261055
transform 1 0 47328 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_493
timestamp 1621261055
transform 1 0 48480 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_1_489
timestamp 1621261055
transform 1 0 48096 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_493
timestamp 1621261055
transform 1 0 48480 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input157
timestamp 1621261055
transform 1 0 48096 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_193
timestamp 1621261055
transform 1 0 48672 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_496
timestamp 1621261055
transform 1 0 48768 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_503
timestamp 1621261055
transform 1 0 49440 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_501
timestamp 1621261055
transform 1 0 49248 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input162
timestamp 1621261055
transform 1 0 49152 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_512
timestamp 1621261055
transform 1 0 50304 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_504
timestamp 1621261055
transform 1 0 49536 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_505
timestamp 1621261055
transform 1 0 49632 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input40
timestamp 1621261055
transform 1 0 50016 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_181
timestamp 1621261055
transform 1 0 49536 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_517
timestamp 1621261055
transform 1 0 50784 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_521
timestamp 1621261055
transform 1 0 51168 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_513
timestamp 1621261055
transform 1 0 50400 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input43
timestamp 1621261055
transform 1 0 51168 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input42
timestamp 1621261055
transform 1 0 50400 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input41
timestamp 1621261055
transform 1 0 50784 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_525
timestamp 1621261055
transform 1 0 51552 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_528
timestamp 1621261055
transform 1 0 51840 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _129_
timestamp 1621261055
transform 1 0 51552 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_533
timestamp 1621261055
transform 1 0 52320 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_533
timestamp 1621261055
transform 1 0 52320 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input44
timestamp 1621261055
transform 1 0 51936 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_182
timestamp 1621261055
transform 1 0 52224 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_1_541
timestamp 1621261055
transform 1 0 53088 0 1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_0_541
timestamp 1621261055
transform 1 0 53088 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input47
timestamp 1621261055
transform 1 0 53472 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input46
timestamp 1621261055
transform 1 0 52704 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input45
timestamp 1621261055
transform 1 0 52704 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_551
timestamp 1621261055
transform 1 0 54048 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_1_549
timestamp 1621261055
transform 1 0 53856 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_0_549
timestamp 1621261055
transform 1 0 53856 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_194
timestamp 1621261055
transform 1 0 53952 0 1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _189_
timestamp 1621261055
transform 1 0 54240 0 -1 3330
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_1_559
timestamp 1621261055
transform 1 0 54816 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_561
timestamp 1621261055
transform 1 0 55008 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_556
timestamp 1621261055
transform 1 0 54528 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input51
timestamp 1621261055
transform 1 0 54432 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_183
timestamp 1621261055
transform 1 0 54912 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_1_567
timestamp 1621261055
transform 1 0 55584 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_0_569
timestamp 1621261055
transform 1 0 55776 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input54
timestamp 1621261055
transform 1 0 55200 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input52
timestamp 1621261055
transform 1 0 55392 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_575
timestamp 1621261055
transform 1 0 56352 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_577
timestamp 1621261055
transform 1 0 56544 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input56
timestamp 1621261055
transform 1 0 55968 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input55
timestamp 1621261055
transform 1 0 56160 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_583
timestamp 1621261055
transform 1 0 57120 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_0_587
timestamp 1621261055
transform 1 0 57504 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_0_585
timestamp 1621261055
transform 1 0 57312 0 -1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input59
timestamp 1621261055
transform 1 0 57504 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input58
timestamp 1621261055
transform 1 0 56736 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_1_591
timestamp 1621261055
transform 1 0 57888 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_0_589
timestamp 1621261055
transform 1 0 57696 0 -1 3330
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_184
timestamp 1621261055
transform 1 0 57600 0 -1 3330
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_1
timestamp 1621261055
transform -1 0 58848 0 -1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_3
timestamp 1621261055
transform -1 0 58848 0 1 3330
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_1_595
timestamp 1621261055
transform 1 0 58272 0 1 3330
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input308
timestamp 1621261055
transform 1 0 1536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_4
timestamp 1621261055
transform 1 0 1152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_8
timestamp 1621261055
transform 1 0 1920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input330
timestamp 1621261055
transform 1 0 2304 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_16
timestamp 1621261055
transform 1 0 2688 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_24
timestamp 1621261055
transform 1 0 3456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input341
timestamp 1621261055
transform 1 0 3072 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_195
timestamp 1621261055
transform 1 0 3840 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_29
timestamp 1621261055
transform 1 0 3936 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input326
timestamp 1621261055
transform 1 0 4320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input305
timestamp 1621261055
transform 1 0 7392 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input328
timestamp 1621261055
transform 1 0 5088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input331
timestamp 1621261055
transform 1 0 5856 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input333
timestamp 1621261055
transform 1 0 6624 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_37
timestamp 1621261055
transform 1 0 4704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_45
timestamp 1621261055
transform 1 0 5472 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_53
timestamp 1621261055
transform 1 0 6240 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_61
timestamp 1621261055
transform 1 0 7008 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_196
timestamp 1621261055
transform 1 0 9120 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input312
timestamp 1621261055
transform 1 0 9600 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input314
timestamp 1621261055
transform 1 0 10368 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input335
timestamp 1621261055
transform 1 0 8160 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_69
timestamp 1621261055
transform 1 0 7776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_77
timestamp 1621261055
transform 1 0 8544 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_81
timestamp 1621261055
transform 1 0 8928 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_84
timestamp 1621261055
transform 1 0 9216 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_92
timestamp 1621261055
transform 1 0 9984 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input206
timestamp 1621261055
transform 1 0 13536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input315
timestamp 1621261055
transform 1 0 11136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input316
timestamp 1621261055
transform 1 0 11904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input317
timestamp 1621261055
transform 1 0 12672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_100
timestamp 1621261055
transform 1 0 10752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_108
timestamp 1621261055
transform 1 0 11520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_116
timestamp 1621261055
transform 1 0 12288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_124
timestamp 1621261055
transform 1 0 13056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_128
timestamp 1621261055
transform 1 0 13440 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_139
timestamp 1621261055
transform 1 0 14496 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_2_137
timestamp 1621261055
transform 1 0 14304 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_133
timestamp 1621261055
transform 1 0 13920 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_197
timestamp 1621261055
transform 1 0 14400 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_147
timestamp 1621261055
transform 1 0 15264 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__buf_1  input144
timestamp 1621261055
transform 1 0 15456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_153
timestamp 1621261055
transform 1 0 15840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input155
timestamp 1621261055
transform 1 0 16224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_161
timestamp 1621261055
transform 1 0 16608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__buf_1  input166
timestamp 1621261055
transform 1 0 16992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_198
timestamp 1621261055
transform 1 0 19680 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input178
timestamp 1621261055
transform 1 0 17760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input198
timestamp 1621261055
transform 1 0 18528 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_169
timestamp 1621261055
transform 1 0 17376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_177
timestamp 1621261055
transform 1 0 18144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_185
timestamp 1621261055
transform 1 0 18912 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_194
timestamp 1621261055
transform 1 0 19776 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_198
timestamp 1621261055
transform 1 0 20160 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__buf_1  input79
timestamp 1621261055
transform 1 0 20256 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input81
timestamp 1621261055
transform 1 0 21024 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input83
timestamp 1621261055
transform 1 0 21792 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input87
timestamp 1621261055
transform 1 0 23232 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_203
timestamp 1621261055
transform 1 0 20640 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_211
timestamp 1621261055
transform 1 0 21408 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_219
timestamp 1621261055
transform 1 0 22176 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_227
timestamp 1621261055
transform 1 0 22944 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_229
timestamp 1621261055
transform 1 0 23136 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_199
timestamp 1621261055
transform 1 0 24960 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input94
timestamp 1621261055
transform 1 0 25440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input96
timestamp 1621261055
transform 1 0 26208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input211
timestamp 1621261055
transform 1 0 24000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_234
timestamp 1621261055
transform 1 0 23616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_242
timestamp 1621261055
transform 1 0 24384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_246
timestamp 1621261055
transform 1 0 24768 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_249
timestamp 1621261055
transform 1 0 25056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_257
timestamp 1621261055
transform 1 0 25824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input97
timestamp 1621261055
transform 1 0 26976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input103
timestamp 1621261055
transform 1 0 28320 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input105
timestamp 1621261055
transform 1 0 29088 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_265
timestamp 1621261055
transform 1 0 26592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_273
timestamp 1621261055
transform 1 0 27360 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_281
timestamp 1621261055
transform 1 0 28128 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_287
timestamp 1621261055
transform 1 0 28704 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_295
timestamp 1621261055
transform 1 0 29472 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_304
timestamp 1621261055
transform 1 0 30336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_200
timestamp 1621261055
transform 1 0 30240 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_308
timestamp 1621261055
transform 1 0 30720 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input110
timestamp 1621261055
transform 1 0 30912 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_314
timestamp 1621261055
transform 1 0 31296 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input113
timestamp 1621261055
transform 1 0 31680 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_322
timestamp 1621261055
transform 1 0 32064 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_328
timestamp 1621261055
transform 1 0 32640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_326
timestamp 1621261055
transform 1 0 32448 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input116
timestamp 1621261055
transform 1 0 32736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_201
timestamp 1621261055
transform 1 0 35520 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input119
timestamp 1621261055
transform 1 0 33888 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input121
timestamp 1621261055
transform 1 0 34656 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input247
timestamp 1621261055
transform 1 0 36000 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_333
timestamp 1621261055
transform 1 0 33120 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_345
timestamp 1621261055
transform 1 0 34272 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_353
timestamp 1621261055
transform 1 0 35040 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_357
timestamp 1621261055
transform 1 0 35424 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_359
timestamp 1621261055
transform 1 0 35616 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _195_
timestamp 1621261055
transform -1 0 38592 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input128
timestamp 1621261055
transform 1 0 36768 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input129
timestamp 1621261055
transform 1 0 37536 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input135
timestamp 1621261055
transform 1 0 38976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_231
timestamp 1621261055
transform -1 0 38304 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_367
timestamp 1621261055
transform 1 0 36384 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_375
timestamp 1621261055
transform 1 0 37152 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_383
timestamp 1621261055
transform 1 0 37920 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_390
timestamp 1621261055
transform 1 0 38592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_398
timestamp 1621261055
transform 1 0 39360 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input137
timestamp 1621261055
transform 1 0 39744 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_412
timestamp 1621261055
transform 1 0 40704 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_410
timestamp 1621261055
transform 1 0 40512 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_406
timestamp 1621261055
transform 1 0 40128 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_202
timestamp 1621261055
transform 1 0 40800 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_422
timestamp 1621261055
transform 1 0 41664 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_2_414
timestamp 1621261055
transform 1 0 40896 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_2_429
timestamp 1621261055
transform 1 0 42336 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_2_424
timestamp 1621261055
transform 1 0 41856 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input143
timestamp 1621261055
transform 1 0 41952 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input145
timestamp 1621261055
transform 1 0 42720 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input148
timestamp 1621261055
transform 1 0 43488 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input152
timestamp 1621261055
transform 1 0 44928 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_437
timestamp 1621261055
transform 1 0 43104 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_445
timestamp 1621261055
transform 1 0 43872 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_453
timestamp 1621261055
transform 1 0 44640 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_455
timestamp 1621261055
transform 1 0 44832 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_2_460
timestamp 1621261055
transform 1 0 45312 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_203
timestamp 1621261055
transform 1 0 46080 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input158
timestamp 1621261055
transform 1 0 46752 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input160
timestamp 1621261055
transform 1 0 47520 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input161
timestamp 1621261055
transform 1 0 48288 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_469
timestamp 1621261055
transform 1 0 46176 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_473
timestamp 1621261055
transform 1 0 46560 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_479
timestamp 1621261055
transform 1 0 47136 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_487
timestamp 1621261055
transform 1 0 47904 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_495
timestamp 1621261055
transform 1 0 48672 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_204
timestamp 1621261055
transform 1 0 51360 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input163
timestamp 1621261055
transform 1 0 49056 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input164
timestamp 1621261055
transform 1 0 49824 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input168
timestamp 1621261055
transform 1 0 50592 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input171
timestamp 1621261055
transform 1 0 51840 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_503
timestamp 1621261055
transform 1 0 49440 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_511
timestamp 1621261055
transform 1 0 50208 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_519
timestamp 1621261055
transform 1 0 50976 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_524
timestamp 1621261055
transform 1 0 51456 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _014_
timestamp 1621261055
transform -1 0 55200 0 -1 4662
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input48
timestamp 1621261055
transform 1 0 52608 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input49
timestamp 1621261055
transform 1 0 53376 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input53
timestamp 1621261055
transform 1 0 54144 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_29
timestamp 1621261055
transform -1 0 54912 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_2_532
timestamp 1621261055
transform 1 0 52224 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_540
timestamp 1621261055
transform 1 0 52992 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_548
timestamp 1621261055
transform 1 0 53760 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_556
timestamp 1621261055
transform 1 0 54528 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_205
timestamp 1621261055
transform 1 0 56640 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input57
timestamp 1621261055
transform 1 0 55584 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input60
timestamp 1621261055
transform 1 0 57120 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_563
timestamp 1621261055
transform 1 0 55200 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_2_571
timestamp 1621261055
transform 1 0 55968 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_575
timestamp 1621261055
transform 1 0 56352 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_2_577
timestamp 1621261055
transform 1 0 56544 0 -1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_2_579
timestamp 1621261055
transform 1 0 56736 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_2_587
timestamp 1621261055
transform 1 0 57504 0 -1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_5
timestamp 1621261055
transform -1 0 58848 0 -1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_2_595
timestamp 1621261055
transform 1 0 58272 0 -1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input329
timestamp 1621261055
transform 1 0 1536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_6
timestamp 1621261055
transform 1 0 1152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_8
timestamp 1621261055
transform 1 0 1920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input352
timestamp 1621261055
transform 1 0 2304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_16
timestamp 1621261055
transform 1 0 2688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_24
timestamp 1621261055
transform 1 0 3456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input355
timestamp 1621261055
transform 1 0 3072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_28
timestamp 1621261055
transform 1 0 3840 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_30
timestamp 1621261055
transform 1 0 4032 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input327
timestamp 1621261055
transform 1 0 4128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_35
timestamp 1621261055
transform 1 0 4512 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_3_48
timestamp 1621261055
transform 1 0 5760 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_43
timestamp 1621261055
transform 1 0 5280 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input332
timestamp 1621261055
transform 1 0 5376 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_56
timestamp 1621261055
transform 1 0 6528 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_54
timestamp 1621261055
transform 1 0 6336 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_52
timestamp 1621261055
transform 1 0 6144 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_206
timestamp 1621261055
transform 1 0 6432 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_64
timestamp 1621261055
transform 1 0 7296 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_71
timestamp 1621261055
transform 1 0 7488 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input334
timestamp 1621261055
transform 1 0 6912 0 1 4662
box -38 -49 422 715
use AND2X1  AND2X1
timestamp 1623617396
transform 1 0 7680 0 1 4662
box 0 -48 1152 714
use sky130_fd_sc_ls__clkbuf_1  input339
timestamp 1621261055
transform 1 0 9216 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input340
timestamp 1621261055
transform 1 0 9984 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_80
timestamp 1621261055
transform 1 0 8832 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_88
timestamp 1621261055
transform 1 0 9600 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_96
timestamp 1621261055
transform 1 0 10368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input343
timestamp 1621261055
transform 1 0 10752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_108
timestamp 1621261055
transform 1 0 11520 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_104
timestamp 1621261055
transform 1 0 11136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_111
timestamp 1621261055
transform 1 0 11808 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_207
timestamp 1621261055
transform 1 0 11712 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input318
timestamp 1621261055
transform 1 0 12192 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_119
timestamp 1621261055
transform 1 0 12576 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input320
timestamp 1621261055
transform 1 0 12960 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_127
timestamp 1621261055
transform 1 0 13344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_131
timestamp 1621261055
transform 1 0 13728 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_208
timestamp 1621261055
transform 1 0 16992 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input217
timestamp 1621261055
transform 1 0 13920 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input228
timestamp 1621261055
transform 1 0 14688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input239
timestamp 1621261055
transform 1 0 15456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input261
timestamp 1621261055
transform 1 0 16224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_137
timestamp 1621261055
transform 1 0 14304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_145
timestamp 1621261055
transform 1 0 15072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_153
timestamp 1621261055
transform 1 0 15840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_161
timestamp 1621261055
transform 1 0 16608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input189
timestamp 1621261055
transform 1 0 17472 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input199
timestamp 1621261055
transform 1 0 18240 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input200
timestamp 1621261055
transform 1 0 19008 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input202
timestamp 1621261055
transform 1 0 19776 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_166
timestamp 1621261055
transform 1 0 17088 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_174
timestamp 1621261055
transform 1 0 17856 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_182
timestamp 1621261055
transform 1 0 18624 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_190
timestamp 1621261055
transform 1 0 19392 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_198
timestamp 1621261055
transform 1 0 20160 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_209
timestamp 1621261055
transform 1 0 22272 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input203
timestamp 1621261055
transform 1 0 20544 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input205
timestamp 1621261055
transform 1 0 21312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input209
timestamp 1621261055
transform 1 0 22752 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_206
timestamp 1621261055
transform 1 0 20928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_214
timestamp 1621261055
transform 1 0 21696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_218
timestamp 1621261055
transform 1 0 22080 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_221
timestamp 1621261055
transform 1 0 22368 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_229
timestamp 1621261055
transform 1 0 23136 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input212
timestamp 1621261055
transform 1 0 23520 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input214
timestamp 1621261055
transform 1 0 24288 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input216
timestamp 1621261055
transform 1 0 25056 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input218
timestamp 1621261055
transform 1 0 25824 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_237
timestamp 1621261055
transform 1 0 23904 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_245
timestamp 1621261055
transform 1 0 24672 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_253
timestamp 1621261055
transform 1 0 25440 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_261
timestamp 1621261055
transform 1 0 26208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input220
timestamp 1621261055
transform 1 0 26592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_273
timestamp 1621261055
transform 1 0 27360 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_269
timestamp 1621261055
transform 1 0 26976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_276
timestamp 1621261055
transform 1 0 27648 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_210
timestamp 1621261055
transform 1 0 27552 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input224
timestamp 1621261055
transform 1 0 28032 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_284
timestamp 1621261055
transform 1 0 28416 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input227
timestamp 1621261055
transform 1 0 28800 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_292
timestamp 1621261055
transform 1 0 29184 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input230
timestamp 1621261055
transform 1 0 29568 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_211
timestamp 1621261055
transform 1 0 32832 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input232
timestamp 1621261055
transform 1 0 30336 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input233
timestamp 1621261055
transform 1 0 31104 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input236
timestamp 1621261055
transform 1 0 31872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_300
timestamp 1621261055
transform 1 0 29952 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_308
timestamp 1621261055
transform 1 0 30720 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_316
timestamp 1621261055
transform 1 0 31488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_324
timestamp 1621261055
transform 1 0 32256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_328
timestamp 1621261055
transform 1 0 32640 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input241
timestamp 1621261055
transform 1 0 33312 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input243
timestamp 1621261055
transform 1 0 34080 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input245
timestamp 1621261055
transform 1 0 34848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input248
timestamp 1621261055
transform 1 0 35616 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_331
timestamp 1621261055
transform 1 0 32928 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_339
timestamp 1621261055
transform 1 0 33696 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_347
timestamp 1621261055
transform 1 0 34464 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_355
timestamp 1621261055
transform 1 0 35232 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_363
timestamp 1621261055
transform 1 0 36000 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_212
timestamp 1621261055
transform 1 0 38112 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input249
timestamp 1621261055
transform 1 0 36384 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input252
timestamp 1621261055
transform 1 0 37152 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input256
timestamp 1621261055
transform 1 0 38592 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_371
timestamp 1621261055
transform 1 0 36768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_379
timestamp 1621261055
transform 1 0 37536 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_383
timestamp 1621261055
transform 1 0 37920 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_386
timestamp 1621261055
transform 1 0 38208 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_394
timestamp 1621261055
transform 1 0 38976 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input258
timestamp 1621261055
transform 1 0 39360 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input260
timestamp 1621261055
transform 1 0 40128 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input264
timestamp 1621261055
transform 1 0 40896 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input265
timestamp 1621261055
transform 1 0 41664 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_402
timestamp 1621261055
transform 1 0 39744 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_410
timestamp 1621261055
transform 1 0 40512 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_418
timestamp 1621261055
transform 1 0 41280 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_426
timestamp 1621261055
transform 1 0 42048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input268
timestamp 1621261055
transform 1 0 42432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_438
timestamp 1621261055
transform 1 0 43200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_434
timestamp 1621261055
transform 1 0 42816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_441
timestamp 1621261055
transform 1 0 43488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_213
timestamp 1621261055
transform 1 0 43392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input273
timestamp 1621261055
transform 1 0 43872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_449
timestamp 1621261055
transform 1 0 44256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input275
timestamp 1621261055
transform 1 0 44640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_457
timestamp 1621261055
transform 1 0 45024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input277
timestamp 1621261055
transform 1 0 45408 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_214
timestamp 1621261055
transform 1 0 48672 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input279
timestamp 1621261055
transform 1 0 46176 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input280
timestamp 1621261055
transform 1 0 46944 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input284
timestamp 1621261055
transform 1 0 47712 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_465
timestamp 1621261055
transform 1 0 45792 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_473
timestamp 1621261055
transform 1 0 46560 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_481
timestamp 1621261055
transform 1 0 47328 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_489
timestamp 1621261055
transform 1 0 48096 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_493
timestamp 1621261055
transform 1 0 48480 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_496
timestamp 1621261055
transform 1 0 48768 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_500
timestamp 1621261055
transform 1 0 49152 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input165
timestamp 1621261055
transform 1 0 49344 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_506
timestamp 1621261055
transform 1 0 49728 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_510
timestamp 1621261055
transform 1 0 50112 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input169
timestamp 1621261055
transform 1 0 50304 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_516
timestamp 1621261055
transform 1 0 50688 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input170
timestamp 1621261055
transform 1 0 51072 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_524
timestamp 1621261055
transform 1 0 51456 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input172
timestamp 1621261055
transform 1 0 51840 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_215
timestamp 1621261055
transform 1 0 53952 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input173
timestamp 1621261055
transform 1 0 52608 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input177
timestamp 1621261055
transform 1 0 54432 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_532
timestamp 1621261055
transform 1 0 52224 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_540
timestamp 1621261055
transform 1 0 52992 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_548
timestamp 1621261055
transform 1 0 53760 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_3_551
timestamp 1621261055
transform 1 0 54048 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_559
timestamp 1621261055
transform 1 0 54816 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input62
timestamp 1621261055
transform 1 0 57024 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input64
timestamp 1621261055
transform 1 0 56256 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input68
timestamp 1621261055
transform 1 0 55488 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_563
timestamp 1621261055
transform 1 0 55200 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_3_565
timestamp 1621261055
transform 1 0 55392 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_3_570
timestamp 1621261055
transform 1 0 55872 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_3_578
timestamp 1621261055
transform 1 0 56640 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_3_586
timestamp 1621261055
transform 1 0 57408 0 1 4662
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_3_594
timestamp 1621261055
transform 1 0 58176 0 1 4662
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_7
timestamp 1621261055
transform -1 0 58848 0 1 4662
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_3_596
timestamp 1621261055
transform 1 0 58368 0 1 4662
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_4_8
timestamp 1621261055
transform 1 0 1920 0 -1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input362
timestamp 1621261055
transform 1 0 1536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_8
timestamp 1621261055
transform 1 0 1152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_16
timestamp 1621261055
transform 1 0 2688 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input356
timestamp 1621261055
transform 1 0 2784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_25
timestamp 1621261055
transform 1 0 3552 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_21
timestamp 1621261055
transform 1 0 3168 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_29
timestamp 1621261055
transform 1 0 3936 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_27
timestamp 1621261055
transform 1 0 3744 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input358
timestamp 1621261055
transform 1 0 4320 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_216
timestamp 1621261055
transform 1 0 3840 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input336
timestamp 1621261055
transform 1 0 6816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input360
timestamp 1621261055
transform 1 0 5088 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output574
timestamp 1621261055
transform 1 0 5856 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_37
timestamp 1621261055
transform 1 0 4704 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_45
timestamp 1621261055
transform 1 0 5472 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_53
timestamp 1621261055
transform 1 0 6240 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_57
timestamp 1621261055
transform 1 0 6624 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_63
timestamp 1621261055
transform 1 0 7200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_217
timestamp 1621261055
transform 1 0 9120 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input337
timestamp 1621261055
transform 1 0 7584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input338
timestamp 1621261055
transform 1 0 8352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input342
timestamp 1621261055
transform 1 0 9600 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input345
timestamp 1621261055
transform 1 0 10368 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_71
timestamp 1621261055
transform 1 0 7968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_79
timestamp 1621261055
transform 1 0 8736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_84
timestamp 1621261055
transform 1 0 9216 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_92
timestamp 1621261055
transform 1 0 9984 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _071_
timestamp 1621261055
transform 1 0 11904 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input321
timestamp 1621261055
transform 1 0 12576 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input347
timestamp 1621261055
transform 1 0 11136 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input351
timestamp 1621261055
transform 1 0 13344 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_100
timestamp 1621261055
transform 1 0 10752 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_108
timestamp 1621261055
transform 1 0 11520 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_115
timestamp 1621261055
transform 1 0 12192 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_123
timestamp 1621261055
transform 1 0 12960 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_131
timestamp 1621261055
transform 1 0 13728 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_135
timestamp 1621261055
transform 1 0 14112 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_139
timestamp 1621261055
transform 1 0 14496 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_137
timestamp 1621261055
transform 1 0 14304 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_218
timestamp 1621261055
transform 1 0 14400 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_4_143
timestamp 1621261055
transform 1 0 14880 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input250
timestamp 1621261055
transform 1 0 14976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_148
timestamp 1621261055
transform 1 0 15360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_156
timestamp 1621261055
transform 1 0 16128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input272
timestamp 1621261055
transform 1 0 15744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input283
timestamp 1621261055
transform 1 0 16512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_164
timestamp 1621261055
transform 1 0 16896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input294
timestamp 1621261055
transform 1 0 17280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_172
timestamp 1621261055
transform 1 0 17664 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_51
timestamp 1621261055
transform 1 0 17856 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_179
timestamp 1621261055
transform 1 0 18336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _048_
timestamp 1621261055
transform 1 0 18048 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_1  input201
timestamp 1621261055
transform 1 0 18720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_187
timestamp 1621261055
transform 1 0 19104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_191
timestamp 1621261055
transform 1 0 19488 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_219
timestamp 1621261055
transform 1 0 19680 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_194
timestamp 1621261055
transform 1 0 19776 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input204
timestamp 1621261055
transform 1 0 20160 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input207
timestamp 1621261055
transform 1 0 20928 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input208
timestamp 1621261055
transform 1 0 21696 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input210
timestamp 1621261055
transform 1 0 22464 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input213
timestamp 1621261055
transform 1 0 23232 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_202
timestamp 1621261055
transform 1 0 20544 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_210
timestamp 1621261055
transform 1 0 21312 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_218
timestamp 1621261055
transform 1 0 22080 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_226
timestamp 1621261055
transform 1 0 22848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_220
timestamp 1621261055
transform 1 0 24960 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input215
timestamp 1621261055
transform 1 0 24000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input219
timestamp 1621261055
transform 1 0 25440 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input221
timestamp 1621261055
transform 1 0 26208 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_234
timestamp 1621261055
transform 1 0 23616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_242
timestamp 1621261055
transform 1 0 24384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_246
timestamp 1621261055
transform 1 0 24768 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_249
timestamp 1621261055
transform 1 0 25056 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_257
timestamp 1621261055
transform 1 0 25824 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input223
timestamp 1621261055
transform 1 0 26976 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input226
timestamp 1621261055
transform 1 0 27744 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input229
timestamp 1621261055
transform 1 0 28512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input231
timestamp 1621261055
transform 1 0 29280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_265
timestamp 1621261055
transform 1 0 26592 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_273
timestamp 1621261055
transform 1 0 27360 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_281
timestamp 1621261055
transform 1 0 28128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_289
timestamp 1621261055
transform 1 0 28896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_297
timestamp 1621261055
transform 1 0 29664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_221
timestamp 1621261055
transform 1 0 30240 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input235
timestamp 1621261055
transform 1 0 30720 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input237
timestamp 1621261055
transform 1 0 31488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input240
timestamp 1621261055
transform 1 0 32256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_301
timestamp 1621261055
transform 1 0 30048 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_304
timestamp 1621261055
transform 1 0 30336 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_312
timestamp 1621261055
transform 1 0 31104 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_320
timestamp 1621261055
transform 1 0 31872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_328
timestamp 1621261055
transform 1 0 32640 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input242
timestamp 1621261055
transform 1 0 33024 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_336
timestamp 1621261055
transform 1 0 33408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_344
timestamp 1621261055
transform 1 0 34176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input244
timestamp 1621261055
transform 1 0 33792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input246
timestamp 1621261055
transform 1 0 34560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_352
timestamp 1621261055
transform 1 0 34944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_356
timestamp 1621261055
transform 1 0 35328 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_222
timestamp 1621261055
transform 1 0 35520 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_359
timestamp 1621261055
transform 1 0 35616 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input251
timestamp 1621261055
transform 1 0 36000 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input253
timestamp 1621261055
transform 1 0 36768 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input255
timestamp 1621261055
transform 1 0 37536 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input257
timestamp 1621261055
transform 1 0 38304 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input259
timestamp 1621261055
transform 1 0 39072 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_367
timestamp 1621261055
transform 1 0 36384 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_375
timestamp 1621261055
transform 1 0 37152 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_383
timestamp 1621261055
transform 1 0 37920 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_391
timestamp 1621261055
transform 1 0 38688 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_223
timestamp 1621261055
transform 1 0 40800 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input263
timestamp 1621261055
transform 1 0 39840 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input267
timestamp 1621261055
transform 1 0 41280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input269
timestamp 1621261055
transform 1 0 42048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_399
timestamp 1621261055
transform 1 0 39456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_407
timestamp 1621261055
transform 1 0 40224 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_411
timestamp 1621261055
transform 1 0 40608 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_414
timestamp 1621261055
transform 1 0 40896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_422
timestamp 1621261055
transform 1 0 41664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input271
timestamp 1621261055
transform 1 0 42816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input274
timestamp 1621261055
transform 1 0 43584 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input276
timestamp 1621261055
transform 1 0 44352 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input278
timestamp 1621261055
transform 1 0 45120 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_430
timestamp 1621261055
transform 1 0 42432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_438
timestamp 1621261055
transform 1 0 43200 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_446
timestamp 1621261055
transform 1 0 43968 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_454
timestamp 1621261055
transform 1 0 44736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_462
timestamp 1621261055
transform 1 0 45504 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_224
timestamp 1621261055
transform 1 0 46080 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input282
timestamp 1621261055
transform 1 0 46560 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input285
timestamp 1621261055
transform 1 0 47328 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input287
timestamp 1621261055
transform 1 0 48096 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_466
timestamp 1621261055
transform 1 0 45888 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_469
timestamp 1621261055
transform 1 0 46176 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_477
timestamp 1621261055
transform 1 0 46944 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_485
timestamp 1621261055
transform 1 0 47712 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_493
timestamp 1621261055
transform 1 0 48480 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input289
timestamp 1621261055
transform 1 0 48864 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_501
timestamp 1621261055
transform 1 0 49248 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_509
timestamp 1621261055
transform 1 0 50016 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input290
timestamp 1621261055
transform 1 0 49632 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input292
timestamp 1621261055
transform 1 0 50400 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_517
timestamp 1621261055
transform 1 0 50784 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_521
timestamp 1621261055
transform 1 0 51168 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_225
timestamp 1621261055
transform 1 0 51360 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_528
timestamp 1621261055
transform 1 0 51840 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_524
timestamp 1621261055
transform 1 0 51456 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input174
timestamp 1621261055
transform 1 0 52128 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input175
timestamp 1621261055
transform 1 0 52896 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input176
timestamp 1621261055
transform 1 0 53664 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input179
timestamp 1621261055
transform 1 0 54432 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_530
timestamp 1621261055
transform 1 0 52032 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_4_535
timestamp 1621261055
transform 1 0 52512 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_543
timestamp 1621261055
transform 1 0 53280 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_551
timestamp 1621261055
transform 1 0 54048 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_559
timestamp 1621261055
transform 1 0 54816 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _104_
timestamp 1621261055
transform 1 0 55200 0 -1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_4_566
timestamp 1621261055
transform 1 0 55488 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input69
timestamp 1621261055
transform 1 0 55872 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_574
timestamp 1621261055
transform 1 0 56256 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_4_579
timestamp 1621261055
transform 1 0 56736 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_226
timestamp 1621261055
transform 1 0 56640 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_4_585
timestamp 1621261055
transform 1 0 57312 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_583
timestamp 1621261055
transform 1 0 57120 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input63
timestamp 1621261055
transform 1 0 57408 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_4_594
timestamp 1621261055
transform 1 0 58176 0 -1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_4_590
timestamp 1621261055
transform 1 0 57792 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_9
timestamp 1621261055
transform -1 0 58848 0 -1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_4_596
timestamp 1621261055
transform 1 0 58368 0 -1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input363
timestamp 1621261055
transform 1 0 1536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_10
timestamp 1621261055
transform 1 0 1152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_8
timestamp 1621261055
transform 1 0 1920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input364
timestamp 1621261055
transform 1 0 2304 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_16
timestamp 1621261055
transform 1 0 2688 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_20
timestamp 1621261055
transform 1 0 3072 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input357
timestamp 1621261055
transform 1 0 3168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_25
timestamp 1621261055
transform 1 0 3552 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_33
timestamp 1621261055
transform 1 0 4320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input359
timestamp 1621261055
transform 1 0 3936 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input361
timestamp 1621261055
transform 1 0 4704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_41
timestamp 1621261055
transform 1 0 5088 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_230
timestamp 1621261055
transform 1 0 5280 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output575
timestamp 1621261055
transform 1 0 5472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_49
timestamp 1621261055
transform 1 0 5856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_56
timestamp 1621261055
transform 1 0 6528 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_53
timestamp 1621261055
transform 1 0 6240 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_227
timestamp 1621261055
transform 1 0 6432 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_232
timestamp 1621261055
transform 1 0 6720 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output577
timestamp 1621261055
transform 1 0 6912 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_64
timestamp 1621261055
transform 1 0 7296 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_87
timestamp 1621261055
transform 1 0 7488 0 1 5994
box -38 -49 230 715
use AND2X2  AND2X2
timestamp 1623617396
transform 1 0 7680 0 1 5994
box 0 -48 1152 714
use sky130_fd_sc_ls__clkbuf_1  input344
timestamp 1621261055
transform 1 0 9408 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input346
timestamp 1621261055
transform 1 0 10176 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_80
timestamp 1621261055
transform 1 0 8832 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_84
timestamp 1621261055
transform 1 0 9216 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_90
timestamp 1621261055
transform 1 0 9792 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_98
timestamp 1621261055
transform 1 0 10560 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input348
timestamp 1621261055
transform 1 0 10944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_106
timestamp 1621261055
transform 1 0 11328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_111
timestamp 1621261055
transform 1 0 11808 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_228
timestamp 1621261055
transform 1 0 11712 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input350
timestamp 1621261055
transform 1 0 12192 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_119
timestamp 1621261055
transform 1 0 12576 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input353
timestamp 1621261055
transform 1 0 12960 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_127
timestamp 1621261055
transform 1 0 13344 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_98
timestamp 1621261055
transform 1 0 13536 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output444
timestamp 1621261055
transform 1 0 13728 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_229
timestamp 1621261055
transform 1 0 16992 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output494
timestamp 1621261055
transform 1 0 14496 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output505
timestamp 1621261055
transform 1 0 15264 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output527
timestamp 1621261055
transform 1 0 16032 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_135
timestamp 1621261055
transform 1 0 14112 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_143
timestamp 1621261055
transform 1 0 14880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_151
timestamp 1621261055
transform 1 0 15648 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_159
timestamp 1621261055
transform 1 0 16416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_163
timestamp 1621261055
transform 1 0 16800 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_166
timestamp 1621261055
transform 1 0 17088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_174
timestamp 1621261055
transform 1 0 17856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output455
timestamp 1621261055
transform 1 0 17472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output475
timestamp 1621261055
transform 1 0 18240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_182
timestamp 1621261055
transform 1 0 18624 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_144
timestamp 1621261055
transform 1 0 18816 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output477
timestamp 1621261055
transform 1 0 19008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_190
timestamp 1621261055
transform 1 0 19392 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_198
timestamp 1621261055
transform 1 0 20160 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output479
timestamp 1621261055
transform 1 0 19776 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_146
timestamp 1621261055
transform 1 0 20352 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output480
timestamp 1621261055
transform 1 0 20544 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_206
timestamp 1621261055
transform 1 0 20928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output482
timestamp 1621261055
transform 1 0 21312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_214
timestamp 1621261055
transform 1 0 21696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_221
timestamp 1621261055
transform 1 0 22368 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_218
timestamp 1621261055
transform 1 0 22080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_230
timestamp 1621261055
transform 1 0 22272 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_150
timestamp 1621261055
transform 1 0 22560 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output487
timestamp 1621261055
transform 1 0 22752 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_229
timestamp 1621261055
transform 1 0 23136 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input222
timestamp 1621261055
transform 1 0 25632 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output489
timestamp 1621261055
transform 1 0 23520 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output491
timestamp 1621261055
transform -1 0 24672 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_154
timestamp 1621261055
transform -1 0 24288 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_237
timestamp 1621261055
transform 1 0 23904 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_245
timestamp 1621261055
transform 1 0 24672 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_253
timestamp 1621261055
transform 1 0 25440 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_5_259
timestamp 1621261055
transform 1 0 26016 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_1  input225
timestamp 1621261055
transform 1 0 26784 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_271
timestamp 1621261055
transform 1 0 27168 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_276
timestamp 1621261055
transform 1 0 27648 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_168
timestamp 1621261055
transform 1 0 27840 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_231
timestamp 1621261055
transform 1 0 27552 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output501
timestamp 1621261055
transform 1 0 28032 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_284
timestamp 1621261055
transform 1 0 28416 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output504
timestamp 1621261055
transform 1 0 28800 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_292
timestamp 1621261055
transform 1 0 29184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_296
timestamp 1621261055
transform 1 0 29568 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input234
timestamp 1621261055
transform 1 0 29664 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_301
timestamp 1621261055
transform 1 0 30048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output509
timestamp 1621261055
transform 1 0 30432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_309
timestamp 1621261055
transform 1 0 30816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input238
timestamp 1621261055
transform 1 0 31200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_317
timestamp 1621261055
transform 1 0 31584 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_180
timestamp 1621261055
transform 1 0 31776 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output513
timestamp 1621261055
transform 1 0 31968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_325
timestamp 1621261055
transform 1 0 32352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_329
timestamp 1621261055
transform 1 0 32736 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_232
timestamp 1621261055
transform 1 0 32832 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output518
timestamp 1621261055
transform 1 0 33312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output520
timestamp 1621261055
transform 1 0 34080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output522
timestamp 1621261055
transform 1 0 34848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_331
timestamp 1621261055
transform 1 0 32928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_339
timestamp 1621261055
transform 1 0 33696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_347
timestamp 1621261055
transform 1 0 34464 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_355
timestamp 1621261055
transform 1 0 35232 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_363
timestamp 1621261055
transform 1 0 36000 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_365
timestamp 1621261055
transform 1 0 36192 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input254
timestamp 1621261055
transform 1 0 36288 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_370
timestamp 1621261055
transform 1 0 36672 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output529
timestamp 1621261055
transform 1 0 37056 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_382
timestamp 1621261055
transform 1 0 37824 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_378
timestamp 1621261055
transform 1 0 37440 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_386
timestamp 1621261055
transform 1 0 38208 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_384
timestamp 1621261055
transform 1 0 38016 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_233
timestamp 1621261055
transform 1 0 38112 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_390
timestamp 1621261055
transform 1 0 38592 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_392
timestamp 1621261055
transform 1 0 38784 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input262
timestamp 1621261055
transform 1 0 38880 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input266
timestamp 1621261055
transform 1 0 40320 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input270
timestamp 1621261055
transform 1 0 41856 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output540
timestamp 1621261055
transform 1 0 41088 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_5_397
timestamp 1621261055
transform 1 0 39264 0 1 5994
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_405
timestamp 1621261055
transform 1 0 40032 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_5_407
timestamp 1621261055
transform 1 0 40224 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_412
timestamp 1621261055
transform 1 0 40704 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_420
timestamp 1621261055
transform 1 0 41472 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_428
timestamp 1621261055
transform 1 0 42240 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output544
timestamp 1621261055
transform 1 0 42624 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_436
timestamp 1621261055
transform 1 0 43008 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_441
timestamp 1621261055
transform 1 0 43488 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_234
timestamp 1621261055
transform 1 0 43392 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output548
timestamp 1621261055
transform 1 0 43872 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_449
timestamp 1621261055
transform 1 0 44256 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output552
timestamp 1621261055
transform 1 0 44640 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_457
timestamp 1621261055
transform 1 0 45024 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_5_461
timestamp 1621261055
transform 1 0 45408 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input281
timestamp 1621261055
transform 1 0 45504 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_466
timestamp 1621261055
transform 1 0 45888 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_69
timestamp 1621261055
transform 1 0 46080 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _053_
timestamp 1621261055
transform 1 0 46272 0 1 5994
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_5_473
timestamp 1621261055
transform 1 0 46560 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_481
timestamp 1621261055
transform 1 0 47328 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input286
timestamp 1621261055
transform 1 0 46944 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input288
timestamp 1621261055
transform 1 0 47712 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_489
timestamp 1621261055
transform 1 0 48096 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_493
timestamp 1621261055
transform 1 0 48480 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_235
timestamp 1621261055
transform 1 0 48672 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_5_496
timestamp 1621261055
transform 1 0 48768 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_504
timestamp 1621261055
transform 1 0 49536 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input291
timestamp 1621261055
transform 1 0 49152 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input293
timestamp 1621261055
transform 1 0 49920 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_512
timestamp 1621261055
transform 1 0 50304 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_100
timestamp 1621261055
transform -1 0 50688 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output445
timestamp 1621261055
transform -1 0 51072 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_520
timestamp 1621261055
transform 1 0 51072 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_105
timestamp 1621261055
transform -1 0 51456 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_528
timestamp 1621261055
transform 1 0 51840 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output447
timestamp 1621261055
transform -1 0 51840 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_107
timestamp 1621261055
transform -1 0 52224 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output448
timestamp 1621261055
transform -1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_536
timestamp 1621261055
transform 1 0 52608 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_540
timestamp 1621261055
transform 1 0 52992 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input192
timestamp 1621261055
transform 1 0 53184 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_546
timestamp 1621261055
transform 1 0 53568 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_551
timestamp 1621261055
transform 1 0 54048 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_236
timestamp 1621261055
transform 1 0 53952 0 1 5994
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input180
timestamp 1621261055
transform 1 0 54432 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_559
timestamp 1621261055
transform 1 0 54816 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input65
timestamp 1621261055
transform 1 0 57696 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input67
timestamp 1621261055
transform 1 0 56928 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input181
timestamp 1621261055
transform 1 0 55200 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input183
timestamp 1621261055
transform 1 0 55968 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_567
timestamp 1621261055
transform 1 0 55584 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_575
timestamp 1621261055
transform 1 0 56352 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_5_579
timestamp 1621261055
transform 1 0 56736 0 1 5994
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_5_585
timestamp 1621261055
transform 1 0 57312 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_5_593
timestamp 1621261055
transform 1 0 58080 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_11
timestamp 1621261055
transform -1 0 58848 0 1 5994
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_8
timestamp 1621261055
transform 1 0 1920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input366
timestamp 1621261055
transform 1 0 1536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_12
timestamp 1621261055
transform 1 0 1152 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_12
timestamp 1621261055
transform 1 0 2304 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input365
timestamp 1621261055
transform 1 0 2496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_26
timestamp 1621261055
transform 1 0 3648 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_18
timestamp 1621261055
transform 1 0 2880 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_6_29
timestamp 1621261055
transform 1 0 3936 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output598
timestamp 1621261055
transform 1 0 4320 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_237
timestamp 1621261055
transform 1 0 3840 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output576
timestamp 1621261055
transform 1 0 5856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output578
timestamp 1621261055
transform 1 0 6624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output579
timestamp 1621261055
transform 1 0 7392 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output601
timestamp 1621261055
transform 1 0 5088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_259
timestamp 1621261055
transform 1 0 4896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_37
timestamp 1621261055
transform 1 0 4704 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_45
timestamp 1621261055
transform 1 0 5472 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_53
timestamp 1621261055
transform 1 0 6240 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_61
timestamp 1621261055
transform 1 0 7008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_69
timestamp 1621261055
transform 1 0 7776 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_234
timestamp 1621261055
transform 1 0 7968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output580
timestamp 1621261055
transform 1 0 8160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_79
timestamp 1621261055
transform 1 0 8736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_235
timestamp 1621261055
transform 1 0 8544 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_84
timestamp 1621261055
transform 1 0 9216 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_238
timestamp 1621261055
transform 1 0 9120 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_237
timestamp 1621261055
transform 1 0 9408 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output582
timestamp 1621261055
transform 1 0 9600 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_92
timestamp 1621261055
transform 1 0 9984 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output585
timestamp 1621261055
transform 1 0 10368 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_104
timestamp 1621261055
transform 1 0 11136 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_100
timestamp 1621261055
transform 1 0 10752 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input349
timestamp 1621261055
transform 1 0 11232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_109
timestamp 1621261055
transform 1 0 11616 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_6_124
timestamp 1621261055
transform 1 0 13056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_119
timestamp 1621261055
transform 1 0 12576 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_117
timestamp 1621261055
transform 1 0 12384 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input354
timestamp 1621261055
transform 1 0 12672 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_132
timestamp 1621261055
transform 1 0 13824 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output483
timestamp 1621261055
transform 1 0 13440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_136
timestamp 1621261055
transform 1 0 14208 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_139
timestamp 1621261055
transform 1 0 14496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_239
timestamp 1621261055
transform 1 0 14400 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output516
timestamp 1621261055
transform 1 0 14880 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_147
timestamp 1621261055
transform 1 0 15264 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output538
timestamp 1621261055
transform 1 0 15648 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_155
timestamp 1621261055
transform 1 0 16032 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_37
timestamp 1621261055
transform 1 0 16224 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _042_
timestamp 1621261055
transform 1 0 16416 0 -1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_162
timestamp 1621261055
transform 1 0 16704 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_131
timestamp 1621261055
transform 1 0 16896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output466
timestamp 1621261055
transform 1 0 17088 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_170
timestamp 1621261055
transform 1 0 17472 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output476
timestamp 1621261055
transform 1 0 17856 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_178
timestamp 1621261055
transform 1 0 18240 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output478
timestamp 1621261055
transform 1 0 18624 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_186
timestamp 1621261055
transform 1 0 19008 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_192
timestamp 1621261055
transform 1 0 19584 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_190
timestamp 1621261055
transform 1 0 19392 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_240
timestamp 1621261055
transform 1 0 19680 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_194
timestamp 1621261055
transform 1 0 19776 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output481
timestamp 1621261055
transform 1 0 20160 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_202
timestamp 1621261055
transform 1 0 20544 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_148
timestamp 1621261055
transform 1 0 20736 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output484
timestamp 1621261055
transform 1 0 20928 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_210
timestamp 1621261055
transform 1 0 21312 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output486
timestamp 1621261055
transform 1 0 21696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_218
timestamp 1621261055
transform 1 0 22080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output488
timestamp 1621261055
transform 1 0 22464 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_226
timestamp 1621261055
transform 1 0 22848 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_152
timestamp 1621261055
transform 1 0 23040 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output490
timestamp 1621261055
transform 1 0 23232 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_234
timestamp 1621261055
transform 1 0 23616 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_156
timestamp 1621261055
transform 1 0 23808 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output492
timestamp 1621261055
transform 1 0 24000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_242
timestamp 1621261055
transform 1 0 24384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_249
timestamp 1621261055
transform 1 0 25056 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_246
timestamp 1621261055
transform 1 0 24768 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_241
timestamp 1621261055
transform 1 0 24960 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output496
timestamp 1621261055
transform 1 0 25440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_257
timestamp 1621261055
transform 1 0 25824 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_162
timestamp 1621261055
transform -1 0 26208 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output498
timestamp 1621261055
transform -1 0 26592 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_265
timestamp 1621261055
transform 1 0 26592 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_166
timestamp 1621261055
transform 1 0 26784 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_273
timestamp 1621261055
transform 1 0 27360 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output500
timestamp 1621261055
transform 1 0 26976 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output503
timestamp 1621261055
transform 1 0 27744 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_281
timestamp 1621261055
transform 1 0 28128 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_170
timestamp 1621261055
transform -1 0 28512 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output506
timestamp 1621261055
transform -1 0 28896 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_289
timestamp 1621261055
transform 1 0 28896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_174
timestamp 1621261055
transform -1 0 29280 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_297
timestamp 1621261055
transform 1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output508
timestamp 1621261055
transform -1 0 29664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_301
timestamp 1621261055
transform 1 0 30048 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_304
timestamp 1621261055
transform 1 0 30336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_242
timestamp 1621261055
transform 1 0 30240 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output512
timestamp 1621261055
transform 1 0 30720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_312
timestamp 1621261055
transform 1 0 31104 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_182
timestamp 1621261055
transform 1 0 31296 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output514
timestamp 1621261055
transform 1 0 31488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_320
timestamp 1621261055
transform 1 0 31872 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output517
timestamp 1621261055
transform 1 0 32256 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_328
timestamp 1621261055
transform 1 0 32640 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output519
timestamp 1621261055
transform 1 0 33024 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_336
timestamp 1621261055
transform 1 0 33408 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_184
timestamp 1621261055
transform -1 0 33792 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_344
timestamp 1621261055
transform 1 0 34176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output521
timestamp 1621261055
transform -1 0 34176 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output524
timestamp 1621261055
transform 1 0 34560 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_352
timestamp 1621261055
transform 1 0 34944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_356
timestamp 1621261055
transform 1 0 35328 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_243
timestamp 1621261055
transform 1 0 35520 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_359
timestamp 1621261055
transform 1 0 35616 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output528
timestamp 1621261055
transform 1 0 36000 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_367
timestamp 1621261055
transform 1 0 36384 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output531
timestamp 1621261055
transform 1 0 36768 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_375
timestamp 1621261055
transform 1 0 37152 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_191
timestamp 1621261055
transform 1 0 37344 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output533
timestamp 1621261055
transform 1 0 37536 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_383
timestamp 1621261055
transform 1 0 37920 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output534
timestamp 1621261055
transform 1 0 38304 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_391
timestamp 1621261055
transform 1 0 38688 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_193
timestamp 1621261055
transform -1 0 39072 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output535
timestamp 1621261055
transform -1 0 39456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_399
timestamp 1621261055
transform 1 0 39456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output537
timestamp 1621261055
transform 1 0 39840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_407
timestamp 1621261055
transform 1 0 40224 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_414
timestamp 1621261055
transform 1 0 40896 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_411
timestamp 1621261055
transform 1 0 40608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_244
timestamp 1621261055
transform 1 0 40800 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_199
timestamp 1621261055
transform -1 0 41280 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output542
timestamp 1621261055
transform -1 0 41664 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_424
timestamp 1621261055
transform 1 0 41856 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_200
timestamp 1621261055
transform -1 0 41856 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output545
timestamp 1621261055
transform 1 0 42048 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_430
timestamp 1621261055
transform 1 0 42432 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_438
timestamp 1621261055
transform 1 0 43200 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output547
timestamp 1621261055
transform 1 0 42816 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output551
timestamp 1621261055
transform 1 0 43584 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_446
timestamp 1621261055
transform 1 0 43968 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_207
timestamp 1621261055
transform -1 0 44352 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output553
timestamp 1621261055
transform -1 0 44736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_454
timestamp 1621261055
transform 1 0 44736 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_462
timestamp 1621261055
transform 1 0 45504 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output555
timestamp 1621261055
transform 1 0 45120 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_466
timestamp 1621261055
transform 1 0 45888 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_469
timestamp 1621261055
transform 1 0 46176 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_212
timestamp 1621261055
transform -1 0 46560 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_245
timestamp 1621261055
transform 1 0 46080 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output558
timestamp 1621261055
transform -1 0 46944 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_477
timestamp 1621261055
transform 1 0 46944 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_216
timestamp 1621261055
transform 1 0 47136 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output561
timestamp 1621261055
transform 1 0 47328 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_485
timestamp 1621261055
transform 1 0 47712 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output563
timestamp 1621261055
transform 1 0 48096 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_493
timestamp 1621261055
transform 1 0 48480 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_223
timestamp 1621261055
transform -1 0 48864 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output565
timestamp 1621261055
transform -1 0 49248 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_503
timestamp 1621261055
transform 1 0 49440 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_224
timestamp 1621261055
transform -1 0 49440 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_6_507
timestamp 1621261055
transform 1 0 49824 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_102
timestamp 1621261055
transform -1 0 50112 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_103
timestamp 1621261055
transform -1 0 50688 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output446
timestamp 1621261055
transform -1 0 50496 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_516
timestamp 1621261055
transform 1 0 50688 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_6_522
timestamp 1621261055
transform 1 0 51264 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_520
timestamp 1621261055
transform 1 0 51072 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_246
timestamp 1621261055
transform 1 0 51360 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_6_524
timestamp 1621261055
transform 1 0 51456 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output449
timestamp 1621261055
transform 1 0 51840 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input182
timestamp 1621261055
transform 1 0 54720 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input196
timestamp 1621261055
transform 1 0 53952 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output451
timestamp 1621261055
transform -1 0 52992 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_110
timestamp 1621261055
transform -1 0 52608 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_532
timestamp 1621261055
transform 1 0 52224 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_6_540
timestamp 1621261055
transform 1 0 52992 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_548
timestamp 1621261055
transform 1 0 53760 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_554
timestamp 1621261055
transform 1 0 54336 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_247
timestamp 1621261055
transform 1 0 56640 0 -1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input66
timestamp 1621261055
transform 1 0 57696 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input184
timestamp 1621261055
transform 1 0 55488 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_6_562
timestamp 1621261055
transform 1 0 55104 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_6_570
timestamp 1621261055
transform 1 0 55872 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_6_579
timestamp 1621261055
transform 1 0 56736 0 -1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_6_587
timestamp 1621261055
transform 1 0 57504 0 -1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_6_593
timestamp 1621261055
transform 1 0 58080 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_13
timestamp 1621261055
transform -1 0 58848 0 -1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output572
timestamp 1621261055
transform 1 0 1536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input367
timestamp 1621261055
transform 1 0 1536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_16
timestamp 1621261055
transform 1 0 1152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_14
timestamp 1621261055
transform 1 0 1152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_8
timestamp 1621261055
transform 1 0 1920 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_8
timestamp 1621261055
transform 1 0 1920 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_241
timestamp 1621261055
transform -1 0 2304 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_228
timestamp 1621261055
transform 1 0 2112 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output584
timestamp 1621261055
transform -1 0 2688 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output573
timestamp 1621261055
transform 1 0 2304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_16
timestamp 1621261055
transform 1 0 2688 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_16
timestamp 1621261055
transform 1 0 2688 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_255
timestamp 1621261055
transform 1 0 2880 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_24
timestamp 1621261055
transform 1 0 3456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_24
timestamp 1621261055
transform 1 0 3456 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output599
timestamp 1621261055
transform 1 0 3072 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output595
timestamp 1621261055
transform 1 0 3072 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_257
timestamp 1621261055
transform 1 0 3648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output600
timestamp 1621261055
transform 1 0 3840 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_258
timestamp 1621261055
transform 1 0 3840 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_29
timestamp 1621261055
transform 1 0 3936 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_32
timestamp 1621261055
transform 1 0 4224 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output603
timestamp 1621261055
transform 1 0 4320 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_37
timestamp 1621261055
transform 1 0 4704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_40
timestamp 1621261055
transform 1 0 4992 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output602
timestamp 1621261055
transform 1 0 4608 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _212_
timestamp 1621261055
transform 1 0 5088 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_44
timestamp 1621261055
transform 1 0 5376 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_48
timestamp 1621261055
transform 1 0 5760 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_261
timestamp 1621261055
transform 1 0 5184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output604
timestamp 1621261055
transform 1 0 5376 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_52
timestamp 1621261055
transform 1 0 6144 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_56
timestamp 1621261055
transform 1 0 6528 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_54
timestamp 1621261055
transform 1 0 6336 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_52
timestamp 1621261055
transform 1 0 6144 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_248
timestamp 1621261055
transform 1 0 6432 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_60
timestamp 1621261055
transform 1 0 6912 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_64
timestamp 1621261055
transform 1 0 7296 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_95
timestamp 1621261055
transform 1 0 7488 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_72
timestamp 1621261055
transform 1 0 8064 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output581
timestamp 1621261055
transform 1 0 7680 0 -1 8658
box -38 -49 422 715
use AOI21X1  AOI21X1
timestamp 1623617396
transform 1 0 7680 0 1 7326
box 0 -48 1152 714
use sky130_fd_sc_ls__diode_2  ANTENNA_239
timestamp 1621261055
transform 1 0 9024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_80
timestamp 1621261055
transform 1 0 8832 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_80
timestamp 1621261055
transform 1 0 8832 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_8_82
timestamp 1621261055
transform 1 0 9024 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_259
timestamp 1621261055
transform 1 0 9120 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output583
timestamp 1621261055
transform 1 0 9216 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_243
timestamp 1621261055
transform 1 0 9408 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_84
timestamp 1621261055
transform 1 0 9216 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output587
timestamp 1621261055
transform 1 0 9600 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_88
timestamp 1621261055
transform 1 0 9600 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_92
timestamp 1621261055
transform 1 0 9984 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_96
timestamp 1621261055
transform 1 0 10368 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_247
timestamp 1621261055
transform 1 0 10176 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_245
timestamp 1621261055
transform 1 0 10560 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output589
timestamp 1621261055
transform 1 0 10368 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output586
timestamp 1621261055
transform 1 0 9984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_100
timestamp 1621261055
transform 1 0 10752 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_249
timestamp 1621261055
transform 1 0 10944 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output588
timestamp 1621261055
transform 1 0 10752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_108
timestamp 1621261055
transform 1 0 11520 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_108
timestamp 1621261055
transform 1 0 11520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_104
timestamp 1621261055
transform 1 0 11136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output590
timestamp 1621261055
transform 1 0 11136 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_111
timestamp 1621261055
transform 1 0 11808 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_251
timestamp 1621261055
transform 1 0 12000 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output592
timestamp 1621261055
transform 1 0 11904 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_249
timestamp 1621261055
transform 1 0 11712 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_116
timestamp 1621261055
transform 1 0 12288 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_253
timestamp 1621261055
transform -1 0 12672 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output591
timestamp 1621261055
transform 1 0 12192 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_119
timestamp 1621261055
transform 1 0 12576 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output594
timestamp 1621261055
transform -1 0 13056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output593
timestamp 1621261055
transform 1 0 12960 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_124
timestamp 1621261055
transform 1 0 13056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_127
timestamp 1621261055
transform 1 0 13344 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_132
timestamp 1621261055
transform 1 0 13824 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output597
timestamp 1621261055
transform 1 0 13440 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output596
timestamp 1621261055
transform 1 0 13728 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_139
timestamp 1621261055
transform 1 0 14496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_136
timestamp 1621261055
transform 1 0 14208 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_135
timestamp 1621261055
transform 1 0 14112 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_260
timestamp 1621261055
transform 1 0 14400 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_147
timestamp 1621261055
transform 1 0 15264 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_147
timestamp 1621261055
transform 1 0 15264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_143
timestamp 1621261055
transform 1 0 14880 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_203
timestamp 1621261055
transform 1 0 15456 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_151
timestamp 1621261055
transform 1 0 15648 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_7_155
timestamp 1621261055
transform 1 0 16032 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_214
timestamp 1621261055
transform 1 0 15840 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output560
timestamp 1621261055
transform 1 0 16032 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output549
timestamp 1621261055
transform 1 0 15648 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_159
timestamp 1621261055
transform 1 0 16416 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_163
timestamp 1621261055
transform 1 0 16800 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output571
timestamp 1621261055
transform 1 0 16800 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_250
timestamp 1621261055
transform 1 0 16992 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_167
timestamp 1621261055
transform 1 0 17184 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_166
timestamp 1621261055
transform 1 0 17088 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_175
timestamp 1621261055
transform 1 0 17952 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_182
timestamp 1621261055
transform 1 0 18624 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_174
timestamp 1621261055
transform 1 0 17856 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_191
timestamp 1621261055
transform 1 0 19488 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_183
timestamp 1621261055
transform 1 0 18720 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_190
timestamp 1621261055
transform 1 0 19392 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_194
timestamp 1621261055
transform 1 0 19776 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_198
timestamp 1621261055
transform 1 0 20160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_261
timestamp 1621261055
transform 1 0 19680 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_202
timestamp 1621261055
transform 1 0 20544 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_202
timestamp 1621261055
transform 1 0 20544 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output485
timestamp 1621261055
transform 1 0 20736 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_210
timestamp 1621261055
transform 1 0 21312 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_208
timestamp 1621261055
transform 1 0 21120 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_218
timestamp 1621261055
transform 1 0 22080 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_221
timestamp 1621261055
transform 1 0 22368 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_216
timestamp 1621261055
transform 1 0 21888 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_251
timestamp 1621261055
transform 1 0 22272 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_226
timestamp 1621261055
transform 1 0 22848 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_229
timestamp 1621261055
transform 1 0 23136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_234
timestamp 1621261055
transform 1 0 23616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_239
timestamp 1621261055
transform 1 0 24096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_158
timestamp 1621261055
transform 1 0 23520 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output493
timestamp 1621261055
transform 1 0 23712 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_246
timestamp 1621261055
transform 1 0 24768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_242
timestamp 1621261055
transform 1 0 24384 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_247
timestamp 1621261055
transform 1 0 24864 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output495
timestamp 1621261055
transform 1 0 24480 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_262
timestamp 1621261055
transform 1 0 24960 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_256
timestamp 1621261055
transform 1 0 25728 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_8_249
timestamp 1621261055
transform 1 0 25056 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_255
timestamp 1621261055
transform 1 0 25632 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_164
timestamp 1621261055
transform -1 0 26016 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_160
timestamp 1621261055
transform 1 0 25056 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output497
timestamp 1621261055
transform 1 0 25248 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _171_
timestamp 1621261055
transform 1 0 25440 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_264
timestamp 1621261055
transform 1 0 26496 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_263
timestamp 1621261055
transform 1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output499
timestamp 1621261055
transform -1 0 26400 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_272
timestamp 1621261055
transform 1 0 27264 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_271
timestamp 1621261055
transform 1 0 27168 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output502
timestamp 1621261055
transform 1 0 26784 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_280
timestamp 1621261055
transform 1 0 28032 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_278
timestamp 1621261055
transform 1 0 27840 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_276
timestamp 1621261055
transform 1 0 27648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_172
timestamp 1621261055
transform -1 0 28128 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output507
timestamp 1621261055
transform -1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_252
timestamp 1621261055
transform 1 0 27552 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_288
timestamp 1621261055
transform 1 0 28800 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_289
timestamp 1621261055
transform 1 0 28896 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_285
timestamp 1621261055
transform 1 0 28512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_176
timestamp 1621261055
transform -1 0 29184 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_296
timestamp 1621261055
transform 1 0 29568 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_296
timestamp 1621261055
transform 1 0 29568 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output510
timestamp 1621261055
transform -1 0 29568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_304
timestamp 1621261055
transform 1 0 30336 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_302
timestamp 1621261055
transform 1 0 30144 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_300
timestamp 1621261055
transform 1 0 29952 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_304
timestamp 1621261055
transform 1 0 30336 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_178
timestamp 1621261055
transform 1 0 29760 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output511
timestamp 1621261055
transform 1 0 29952 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_263
timestamp 1621261055
transform 1 0 30240 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_312
timestamp 1621261055
transform 1 0 31104 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_310
timestamp 1621261055
transform 1 0 30912 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_308
timestamp 1621261055
transform 1 0 30720 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output515
timestamp 1621261055
transform 1 0 31008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_320
timestamp 1621261055
transform 1 0 31872 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_322
timestamp 1621261055
transform 1 0 32064 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_315
timestamp 1621261055
transform 1 0 31392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _116_
timestamp 1621261055
transform 1 0 31776 0 1 7326
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_328
timestamp 1621261055
transform 1 0 32640 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_324
timestamp 1621261055
transform 1 0 32256 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_253
timestamp 1621261055
transform 1 0 32832 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _152_
timestamp 1621261055
transform 1 0 32352 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_336
timestamp 1621261055
transform 1 0 33408 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_7_335
timestamp 1621261055
transform 1 0 33312 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_331
timestamp 1621261055
transform 1 0 32928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_186
timestamp 1621261055
transform -1 0 33600 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output523
timestamp 1621261055
transform -1 0 33984 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_344
timestamp 1621261055
transform 1 0 34176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_342
timestamp 1621261055
transform 1 0 33984 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_188
timestamp 1621261055
transform 1 0 34176 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output525
timestamp 1621261055
transform 1 0 34368 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_356
timestamp 1621261055
transform 1 0 35328 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_352
timestamp 1621261055
transform 1 0 34944 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_350
timestamp 1621261055
transform 1 0 34752 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output526
timestamp 1621261055
transform 1 0 35136 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_359
timestamp 1621261055
transform 1 0 35616 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_358
timestamp 1621261055
transform 1 0 35520 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output530
timestamp 1621261055
transform 1 0 35904 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_264
timestamp 1621261055
transform 1 0 35520 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_367
timestamp 1621261055
transform 1 0 36384 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_366
timestamp 1621261055
transform 1 0 36288 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_189
timestamp 1621261055
transform -1 0 36672 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output532
timestamp 1621261055
transform -1 0 37056 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_375
timestamp 1621261055
transform 1 0 37152 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_374
timestamp 1621261055
transform 1 0 37056 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_383
timestamp 1621261055
transform 1 0 37920 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_386
timestamp 1621261055
transform 1 0 38208 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_7_384
timestamp 1621261055
transform 1 0 38016 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_382
timestamp 1621261055
transform 1 0 37824 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_195
timestamp 1621261055
transform -1 0 38592 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_254
timestamp 1621261055
transform 1 0 38112 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_391
timestamp 1621261055
transform 1 0 38688 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_394
timestamp 1621261055
transform 1 0 38976 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_197
timestamp 1621261055
transform -1 0 39360 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output536
timestamp 1621261055
transform -1 0 38976 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_399
timestamp 1621261055
transform 1 0 39456 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_402
timestamp 1621261055
transform 1 0 39744 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output539
timestamp 1621261055
transform -1 0 39744 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_411
timestamp 1621261055
transform 1 0 40608 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_407
timestamp 1621261055
transform 1 0 40224 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_410
timestamp 1621261055
transform 1 0 40512 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output541
timestamp 1621261055
transform 1 0 40128 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_265
timestamp 1621261055
transform 1 0 40800 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_422
timestamp 1621261055
transform 1 0 41664 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_414
timestamp 1621261055
transform 1 0 40896 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_418
timestamp 1621261055
transform 1 0 41280 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_201
timestamp 1621261055
transform -1 0 41664 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output546
timestamp 1621261055
transform -1 0 42048 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output543
timestamp 1621261055
transform 1 0 40896 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_426
timestamp 1621261055
transform 1 0 42048 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_205
timestamp 1621261055
transform 1 0 42240 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_8_430
timestamp 1621261055
transform 1 0 42432 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_434
timestamp 1621261055
transform 1 0 42816 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output550
timestamp 1621261055
transform 1 0 42432 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_446
timestamp 1621261055
transform 1 0 43968 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_8_438
timestamp 1621261055
transform 1 0 43200 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_441
timestamp 1621261055
transform 1 0 43488 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_438
timestamp 1621261055
transform 1 0 43200 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_209
timestamp 1621261055
transform 1 0 43680 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output554
timestamp 1621261055
transform 1 0 43872 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_255
timestamp 1621261055
transform 1 0 43392 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_454
timestamp 1621261055
transform 1 0 44736 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_449
timestamp 1621261055
transform 1 0 44256 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output556
timestamp 1621261055
transform 1 0 44640 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_458
timestamp 1621261055
transform 1 0 45120 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_457
timestamp 1621261055
transform 1 0 45024 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_210
timestamp 1621261055
transform -1 0 45408 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output557
timestamp 1621261055
transform -1 0 45792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _122_
timestamp 1621261055
transform 1 0 45312 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_469
timestamp 1621261055
transform 1 0 46176 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_8_467
timestamp 1621261055
transform 1 0 45984 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_463
timestamp 1621261055
transform 1 0 45600 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_465
timestamp 1621261055
transform 1 0 45792 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output559
timestamp 1621261055
transform 1 0 46176 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_266
timestamp 1621261055
transform 1 0 46080 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_477
timestamp 1621261055
transform 1 0 46944 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_473
timestamp 1621261055
transform 1 0 46560 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_218
timestamp 1621261055
transform -1 0 46944 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output562
timestamp 1621261055
transform -1 0 47328 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_8_487
timestamp 1621261055
transform 1 0 47904 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_485
timestamp 1621261055
transform 1 0 47712 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_481
timestamp 1621261055
transform 1 0 47328 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_220
timestamp 1621261055
transform -1 0 47712 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output566
timestamp 1621261055
transform 1 0 48000 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output564
timestamp 1621261055
transform -1 0 48096 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_492
timestamp 1621261055
transform 1 0 48384 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_7_491
timestamp 1621261055
transform 1 0 48288 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_226
timestamp 1621261055
transform -1 0 48768 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_221
timestamp 1621261055
transform -1 0 48288 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_256
timestamp 1621261055
transform 1 0 48672 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_8_500
timestamp 1621261055
transform 1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_496
timestamp 1621261055
transform 1 0 48768 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output568
timestamp 1621261055
transform -1 0 49152 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output567
timestamp 1621261055
transform 1 0 49152 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_508
timestamp 1621261055
transform 1 0 49920 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_512
timestamp 1621261055
transform 1 0 50304 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_504
timestamp 1621261055
transform 1 0 49536 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output570
timestamp 1621261055
transform 1 0 49536 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output569
timestamp 1621261055
transform 1 0 49920 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _192_
timestamp 1621261055
transform 1 0 50304 0 -1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_8_515
timestamp 1621261055
transform 1 0 50592 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_141
timestamp 1621261055
transform -1 0 50880 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output473
timestamp 1621261055
transform -1 0 51264 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_528
timestamp 1621261055
transform 1 0 51840 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_8_524
timestamp 1621261055
transform 1 0 51456 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_522
timestamp 1621261055
transform 1 0 51264 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_108
timestamp 1621261055
transform -1 0 51648 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output450
timestamp 1621261055
transform -1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_267
timestamp 1621261055
transform 1 0 51360 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_530
timestamp 1621261055
transform 1 0 52032 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_7_530
timestamp 1621261055
transform 1 0 52032 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_138
timestamp 1621261055
transform -1 0 52320 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output472
timestamp 1621261055
transform -1 0 52704 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output452
timestamp 1621261055
transform 1 0 52416 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_545
timestamp 1621261055
transform 1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_538
timestamp 1621261055
transform 1 0 52800 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_139
timestamp 1621261055
transform -1 0 52896 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_112
timestamp 1621261055
transform -1 0 53088 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output454
timestamp 1621261055
transform -1 0 53472 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output453
timestamp 1621261055
transform 1 0 53184 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_8_553
timestamp 1621261055
transform 1 0 54240 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_7_551
timestamp 1621261055
transform 1 0 54048 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_7_546
timestamp 1621261055
transform 1 0 53568 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output456
timestamp 1621261055
transform 1 0 53856 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_257
timestamp 1621261055
transform 1 0 53952 0 1 7326
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_8_561
timestamp 1621261055
transform 1 0 55008 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_7_559
timestamp 1621261055
transform 1 0 54816 0 1 7326
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input194
timestamp 1621261055
transform 1 0 55008 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_566
timestamp 1621261055
transform 1 0 55488 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_565
timestamp 1621261055
transform 1 0 55392 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input197
timestamp 1621261055
transform 1 0 55104 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input185
timestamp 1621261055
transform 1 0 55776 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_8_574
timestamp 1621261055
transform 1 0 56256 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_573
timestamp 1621261055
transform 1 0 56160 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input193
timestamp 1621261055
transform 1 0 55872 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input186
timestamp 1621261055
transform 1 0 56544 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_268
timestamp 1621261055
transform 1 0 56640 0 -1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_8_587
timestamp 1621261055
transform 1 0 57504 0 -1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_8_579
timestamp 1621261055
transform 1 0 56736 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_7_581
timestamp 1621261055
transform 1 0 56928 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input188
timestamp 1621261055
transform 1 0 57120 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input187
timestamp 1621261055
transform 1 0 57312 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_7_589
timestamp 1621261055
transform 1 0 57696 0 1 7326
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_15
timestamp 1621261055
transform -1 0 58848 0 1 7326
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_17
timestamp 1621261055
transform -1 0 58848 0 -1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_8_595
timestamp 1621261055
transform 1 0 58272 0 -1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_18
timestamp 1621261055
transform 1 0 1152 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_4
timestamp 1621261055
transform 1 0 1536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_12
timestamp 1621261055
transform 1 0 2304 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_20
timestamp 1621261055
transform 1 0 3072 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_28
timestamp 1621261055
transform 1 0 3840 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_269
timestamp 1621261055
transform 1 0 6432 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_43
timestamp 1621261055
transform 1 0 7488 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_36
timestamp 1621261055
transform 1 0 4608 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_44
timestamp 1621261055
transform 1 0 5376 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_52
timestamp 1621261055
transform 1 0 6144 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_54
timestamp 1621261055
transform 1 0 6336 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_56
timestamp 1621261055
transform 1 0 6528 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_64
timestamp 1621261055
transform 1 0 7296 0 1 8658
box -38 -49 230 715
use AOI22X1  AOI22X1
timestamp 1623617396
transform 1 0 7680 0 1 8658
box 0 -48 1440 714
use sky130_fd_sc_ls__conb_1  _167_
timestamp 1621261055
transform 1 0 9696 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_118
timestamp 1621261055
transform 1 0 9504 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_9_83
timestamp 1621261055
transform 1 0 9120 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_92
timestamp 1621261055
transform 1 0 9984 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _046_
timestamp 1621261055
transform 1 0 12192 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_270
timestamp 1621261055
transform 1 0 11712 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_45
timestamp 1621261055
transform 1 0 12000 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_100
timestamp 1621261055
transform 1 0 10752 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_108
timestamp 1621261055
transform 1 0 11520 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_111
timestamp 1621261055
transform 1 0 11808 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_118
timestamp 1621261055
transform 1 0 12480 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_126
timestamp 1621261055
transform 1 0 13248 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_271
timestamp 1621261055
transform 1 0 16992 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_134
timestamp 1621261055
transform 1 0 14016 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_142
timestamp 1621261055
transform 1 0 14784 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_150
timestamp 1621261055
transform 1 0 15552 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_158
timestamp 1621261055
transform 1 0 16320 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_162
timestamp 1621261055
transform 1 0 16704 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_164
timestamp 1621261055
transform 1 0 16896 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_166
timestamp 1621261055
transform 1 0 17088 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_174
timestamp 1621261055
transform 1 0 17856 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_182
timestamp 1621261055
transform 1 0 18624 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_190
timestamp 1621261055
transform 1 0 19392 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_198
timestamp 1621261055
transform 1 0 20160 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_272
timestamp 1621261055
transform 1 0 22272 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_206
timestamp 1621261055
transform 1 0 20928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_214
timestamp 1621261055
transform 1 0 21696 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_218
timestamp 1621261055
transform 1 0 22080 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_221
timestamp 1621261055
transform 1 0 22368 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_229
timestamp 1621261055
transform 1 0 23136 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_237
timestamp 1621261055
transform 1 0 23904 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_245
timestamp 1621261055
transform 1 0 24672 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_253
timestamp 1621261055
transform 1 0 25440 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_261
timestamp 1621261055
transform 1 0 26208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_273
timestamp 1621261055
transform 1 0 27552 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_269
timestamp 1621261055
transform 1 0 26976 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_273
timestamp 1621261055
transform 1 0 27360 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_276
timestamp 1621261055
transform 1 0 27648 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_284
timestamp 1621261055
transform 1 0 28416 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_292
timestamp 1621261055
transform 1 0 29184 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_274
timestamp 1621261055
transform 1 0 32832 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_300
timestamp 1621261055
transform 1 0 29952 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_308
timestamp 1621261055
transform 1 0 30720 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_316
timestamp 1621261055
transform 1 0 31488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_324
timestamp 1621261055
transform 1 0 32256 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_328
timestamp 1621261055
transform 1 0 32640 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_331
timestamp 1621261055
transform 1 0 32928 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_339
timestamp 1621261055
transform 1 0 33696 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_347
timestamp 1621261055
transform 1 0 34464 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_355
timestamp 1621261055
transform 1 0 35232 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_363
timestamp 1621261055
transform 1 0 36000 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_275
timestamp 1621261055
transform 1 0 38112 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_371
timestamp 1621261055
transform 1 0 36768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_379
timestamp 1621261055
transform 1 0 37536 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_383
timestamp 1621261055
transform 1 0 37920 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_386
timestamp 1621261055
transform 1 0 38208 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_394
timestamp 1621261055
transform 1 0 38976 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_402
timestamp 1621261055
transform 1 0 39744 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_410
timestamp 1621261055
transform 1 0 40512 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_418
timestamp 1621261055
transform 1 0 41280 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_426
timestamp 1621261055
transform 1 0 42048 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_276
timestamp 1621261055
transform 1 0 43392 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_434
timestamp 1621261055
transform 1 0 42816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_438
timestamp 1621261055
transform 1 0 43200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_441
timestamp 1621261055
transform 1 0 43488 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_449
timestamp 1621261055
transform 1 0 44256 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_457
timestamp 1621261055
transform 1 0 45024 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _142_
timestamp 1621261055
transform 1 0 46080 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_277
timestamp 1621261055
transform 1 0 48672 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_465
timestamp 1621261055
transform 1 0 45792 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_9_467
timestamp 1621261055
transform 1 0 45984 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_9_471
timestamp 1621261055
transform 1 0 46368 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_479
timestamp 1621261055
transform 1 0 47136 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_487
timestamp 1621261055
transform 1 0 47904 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _018_
timestamp 1621261055
transform 1 0 51456 0 1 8658
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_31
timestamp 1621261055
transform 1 0 51264 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_496
timestamp 1621261055
transform 1 0 48768 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_504
timestamp 1621261055
transform 1 0 49536 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_9_512
timestamp 1621261055
transform 1 0 50304 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_520
timestamp 1621261055
transform 1 0 51072 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_9_527
timestamp 1621261055
transform 1 0 51744 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_9_535
timestamp 1621261055
transform 1 0 52512 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_541
timestamp 1621261055
transform 1 0 53088 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_539
timestamp 1621261055
transform 1 0 52896 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output469
timestamp 1621261055
transform 1 0 53184 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_9_546
timestamp 1621261055
transform 1 0 53568 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_551
timestamp 1621261055
transform 1 0 54048 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_278
timestamp 1621261055
transform 1 0 53952 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_113
timestamp 1621261055
transform -1 0 54432 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output457
timestamp 1621261055
transform -1 0 54816 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_9_559
timestamp 1621261055
transform 1 0 54816 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_117
timestamp 1621261055
transform -1 0 55200 0 1 8658
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input190
timestamp 1621261055
transform 1 0 57216 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input195
timestamp 1621261055
transform 1 0 56448 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output459
timestamp 1621261055
transform -1 0 55584 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_567
timestamp 1621261055
transform 1 0 55584 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_9_575
timestamp 1621261055
transform 1 0 56352 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_9_580
timestamp 1621261055
transform 1 0 56832 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_9_588
timestamp 1621261055
transform 1 0 57600 0 1 8658
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_19
timestamp 1621261055
transform -1 0 58848 0 1 8658
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_9_596
timestamp 1621261055
transform 1 0 58368 0 1 8658
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_20
timestamp 1621261055
transform 1 0 1152 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_279
timestamp 1621261055
transform 1 0 3840 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_4
timestamp 1621261055
transform 1 0 1536 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_12
timestamp 1621261055
transform 1 0 2304 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_20
timestamp 1621261055
transform 1 0 3072 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_29
timestamp 1621261055
transform 1 0 3936 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _060_
timestamp 1621261055
transform 1 0 5472 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_10_37
timestamp 1621261055
transform 1 0 4704 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_48
timestamp 1621261055
transform 1 0 5760 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_56
timestamp 1621261055
transform 1 0 6528 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_64
timestamp 1621261055
transform 1 0 7296 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_280
timestamp 1621261055
transform 1 0 9120 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_72
timestamp 1621261055
transform 1 0 8064 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_80
timestamp 1621261055
transform 1 0 8832 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_82
timestamp 1621261055
transform 1 0 9024 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_84
timestamp 1621261055
transform 1 0 9216 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_92
timestamp 1621261055
transform 1 0 9984 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_100
timestamp 1621261055
transform 1 0 10752 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_108
timestamp 1621261055
transform 1 0 11520 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_116
timestamp 1621261055
transform 1 0 12288 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_124
timestamp 1621261055
transform 1 0 13056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_132
timestamp 1621261055
transform 1 0 13824 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_281
timestamp 1621261055
transform 1 0 14400 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_136
timestamp 1621261055
transform 1 0 14208 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_139
timestamp 1621261055
transform 1 0 14496 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_147
timestamp 1621261055
transform 1 0 15264 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_155
timestamp 1621261055
transform 1 0 16032 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_163
timestamp 1621261055
transform 1 0 16800 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_282
timestamp 1621261055
transform 1 0 19680 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_171
timestamp 1621261055
transform 1 0 17568 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_179
timestamp 1621261055
transform 1 0 18336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_187
timestamp 1621261055
transform 1 0 19104 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_191
timestamp 1621261055
transform 1 0 19488 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_194
timestamp 1621261055
transform 1 0 19776 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_202
timestamp 1621261055
transform 1 0 20544 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_210
timestamp 1621261055
transform 1 0 21312 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_218
timestamp 1621261055
transform 1 0 22080 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_226
timestamp 1621261055
transform 1 0 22848 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_283
timestamp 1621261055
transform 1 0 24960 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_234
timestamp 1621261055
transform 1 0 23616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_242
timestamp 1621261055
transform 1 0 24384 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_246
timestamp 1621261055
transform 1 0 24768 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_249
timestamp 1621261055
transform 1 0 25056 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_257
timestamp 1621261055
transform 1 0 25824 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _073_
timestamp 1621261055
transform 1 0 28416 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_10_265
timestamp 1621261055
transform 1 0 26592 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_273
timestamp 1621261055
transform 1 0 27360 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_281
timestamp 1621261055
transform 1 0 28128 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_283
timestamp 1621261055
transform 1 0 28320 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_287
timestamp 1621261055
transform 1 0 28704 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_295
timestamp 1621261055
transform 1 0 29472 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_284
timestamp 1621261055
transform 1 0 30240 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_304
timestamp 1621261055
transform 1 0 30336 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_312
timestamp 1621261055
transform 1 0 31104 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_320
timestamp 1621261055
transform 1 0 31872 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_328
timestamp 1621261055
transform 1 0 32640 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_285
timestamp 1621261055
transform 1 0 35520 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_336
timestamp 1621261055
transform 1 0 33408 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_344
timestamp 1621261055
transform 1 0 34176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_352
timestamp 1621261055
transform 1 0 34944 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_356
timestamp 1621261055
transform 1 0 35328 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_359
timestamp 1621261055
transform 1 0 35616 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _114_
timestamp 1621261055
transform 1 0 36576 0 -1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_367
timestamp 1621261055
transform 1 0 36384 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_372
timestamp 1621261055
transform 1 0 36864 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_380
timestamp 1621261055
transform 1 0 37632 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_388
timestamp 1621261055
transform 1 0 38400 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_396
timestamp 1621261055
transform 1 0 39168 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_286
timestamp 1621261055
transform 1 0 40800 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_404
timestamp 1621261055
transform 1 0 39936 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_10_412
timestamp 1621261055
transform 1 0 40704 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_414
timestamp 1621261055
transform 1 0 40896 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_422
timestamp 1621261055
transform 1 0 41664 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_430
timestamp 1621261055
transform 1 0 42432 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_438
timestamp 1621261055
transform 1 0 43200 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_446
timestamp 1621261055
transform 1 0 43968 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_454
timestamp 1621261055
transform 1 0 44736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_462
timestamp 1621261055
transform 1 0 45504 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_287
timestamp 1621261055
transform 1 0 46080 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_466
timestamp 1621261055
transform 1 0 45888 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_469
timestamp 1621261055
transform 1 0 46176 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_477
timestamp 1621261055
transform 1 0 46944 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_485
timestamp 1621261055
transform 1 0 47712 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_493
timestamp 1621261055
transform 1 0 48480 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_288
timestamp 1621261055
transform 1 0 51360 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_501
timestamp 1621261055
transform 1 0 49248 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_509
timestamp 1621261055
transform 1 0 50016 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_517
timestamp 1621261055
transform 1 0 50784 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_521
timestamp 1621261055
transform 1 0 51168 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_524
timestamp 1621261055
transform 1 0 51456 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output458
timestamp 1621261055
transform -1 0 54624 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output460
timestamp 1621261055
transform -1 0 55392 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_115
timestamp 1621261055
transform -1 0 54240 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_116
timestamp 1621261055
transform -1 0 54816 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_119
timestamp 1621261055
transform -1 0 55008 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_10_532
timestamp 1621261055
transform 1 0 52224 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_10_540
timestamp 1621261055
transform 1 0 52992 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_548
timestamp 1621261055
transform 1 0 53760 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_10_550
timestamp 1621261055
transform 1 0 53952 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_10_565
timestamp 1621261055
transform 1 0 55392 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_121
timestamp 1621261055
transform 1 0 55584 0 -1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output461
timestamp 1621261055
transform 1 0 55776 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_577
timestamp 1621261055
transform 1 0 56544 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_10_573
timestamp 1621261055
transform 1 0 56160 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_289
timestamp 1621261055
transform 1 0 56640 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_10_587
timestamp 1621261055
transform 1 0 57504 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_10_579
timestamp 1621261055
transform 1 0 56736 0 -1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_10_592
timestamp 1621261055
transform 1 0 57984 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input191
timestamp 1621261055
transform 1 0 57600 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_21
timestamp 1621261055
transform -1 0 58848 0 -1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_10_596
timestamp 1621261055
transform 1 0 58368 0 -1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_22
timestamp 1621261055
transform 1 0 1152 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_4
timestamp 1621261055
transform 1 0 1536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_12
timestamp 1621261055
transform 1 0 2304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_20
timestamp 1621261055
transform 1 0 3072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_28
timestamp 1621261055
transform 1 0 3840 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_32
timestamp 1621261055
transform 1 0 4224 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _203_
timestamp 1621261055
transform 1 0 4416 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_290
timestamp 1621261055
transform 1 0 6432 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_47
timestamp 1621261055
transform 1 0 7488 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_37
timestamp 1621261055
transform 1 0 4704 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_45
timestamp 1621261055
transform 1 0 5472 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_53
timestamp 1621261055
transform 1 0 6240 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_56
timestamp 1621261055
transform 1 0 6528 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_64
timestamp 1621261055
transform 1 0 7296 0 1 9990
box -38 -49 230 715
use BUFX2  BUFX2
timestamp 1623617396
transform 1 0 7680 0 1 9990
box 0 -48 864 714
use sky130_fd_sc_ls__decap_8  FILLER_11_77
timestamp 1621261055
transform 1 0 8544 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_85
timestamp 1621261055
transform 1 0 9312 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_93
timestamp 1621261055
transform 1 0 10080 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_291
timestamp 1621261055
transform 1 0 11712 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_101
timestamp 1621261055
transform 1 0 10848 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_11_109
timestamp 1621261055
transform 1 0 11616 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_111
timestamp 1621261055
transform 1 0 11808 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_119
timestamp 1621261055
transform 1 0 12576 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_127
timestamp 1621261055
transform 1 0 13344 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_292
timestamp 1621261055
transform 1 0 16992 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_135
timestamp 1621261055
transform 1 0 14112 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_143
timestamp 1621261055
transform 1 0 14880 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_151
timestamp 1621261055
transform 1 0 15648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_159
timestamp 1621261055
transform 1 0 16416 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_163
timestamp 1621261055
transform 1 0 16800 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_166
timestamp 1621261055
transform 1 0 17088 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_174
timestamp 1621261055
transform 1 0 17856 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_182
timestamp 1621261055
transform 1 0 18624 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_190
timestamp 1621261055
transform 1 0 19392 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_198
timestamp 1621261055
transform 1 0 20160 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_293
timestamp 1621261055
transform 1 0 22272 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_206
timestamp 1621261055
transform 1 0 20928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_214
timestamp 1621261055
transform 1 0 21696 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_218
timestamp 1621261055
transform 1 0 22080 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_221
timestamp 1621261055
transform 1 0 22368 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_229
timestamp 1621261055
transform 1 0 23136 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_237
timestamp 1621261055
transform 1 0 23904 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_245
timestamp 1621261055
transform 1 0 24672 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_253
timestamp 1621261055
transform 1 0 25440 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_261
timestamp 1621261055
transform 1 0 26208 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_294
timestamp 1621261055
transform 1 0 27552 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_269
timestamp 1621261055
transform 1 0 26976 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_273
timestamp 1621261055
transform 1 0 27360 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_276
timestamp 1621261055
transform 1 0 27648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_284
timestamp 1621261055
transform 1 0 28416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_292
timestamp 1621261055
transform 1 0 29184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_295
timestamp 1621261055
transform 1 0 32832 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_300
timestamp 1621261055
transform 1 0 29952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_308
timestamp 1621261055
transform 1 0 30720 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_316
timestamp 1621261055
transform 1 0 31488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_324
timestamp 1621261055
transform 1 0 32256 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_328
timestamp 1621261055
transform 1 0 32640 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_331
timestamp 1621261055
transform 1 0 32928 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_339
timestamp 1621261055
transform 1 0 33696 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_347
timestamp 1621261055
transform 1 0 34464 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_355
timestamp 1621261055
transform 1 0 35232 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_363
timestamp 1621261055
transform 1 0 36000 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _102_
timestamp 1621261055
transform 1 0 38592 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_296
timestamp 1621261055
transform 1 0 38112 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_371
timestamp 1621261055
transform 1 0 36768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_379
timestamp 1621261055
transform 1 0 37536 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_383
timestamp 1621261055
transform 1 0 37920 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_386
timestamp 1621261055
transform 1 0 38208 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_393
timestamp 1621261055
transform 1 0 38880 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_401
timestamp 1621261055
transform 1 0 39648 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_409
timestamp 1621261055
transform 1 0 40416 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_417
timestamp 1621261055
transform 1 0 41184 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_425
timestamp 1621261055
transform 1 0 41952 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_297
timestamp 1621261055
transform 1 0 43392 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_11_433
timestamp 1621261055
transform 1 0 42720 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_437
timestamp 1621261055
transform 1 0 43104 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_439
timestamp 1621261055
transform 1 0 43296 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_441
timestamp 1621261055
transform 1 0 43488 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_449
timestamp 1621261055
transform 1 0 44256 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_457
timestamp 1621261055
transform 1 0 45024 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _083_
timestamp 1621261055
transform 1 0 45888 0 1 9990
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_298
timestamp 1621261055
transform 1 0 48672 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_11_465
timestamp 1621261055
transform 1 0 45792 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_11_469
timestamp 1621261055
transform 1 0 46176 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_477
timestamp 1621261055
transform 1 0 46944 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_485
timestamp 1621261055
transform 1 0 47712 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_493
timestamp 1621261055
transform 1 0 48480 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_496
timestamp 1621261055
transform 1 0 48768 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_504
timestamp 1621261055
transform 1 0 49536 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_512
timestamp 1621261055
transform 1 0 50304 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_520
timestamp 1621261055
transform 1 0 51072 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_11_528
timestamp 1621261055
transform 1 0 51840 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_299
timestamp 1621261055
transform 1 0 53952 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output471
timestamp 1621261055
transform -1 0 55296 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_136
timestamp 1621261055
transform -1 0 54912 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_11_536
timestamp 1621261055
transform 1 0 52608 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_11_544
timestamp 1621261055
transform 1 0 53376 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_548
timestamp 1621261055
transform 1 0 53760 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_11_551
timestamp 1621261055
transform 1 0 54048 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_555
timestamp 1621261055
transform 1 0 54432 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_11_557
timestamp 1621261055
transform 1 0 54624 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_564
timestamp 1621261055
transform 1 0 55296 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_123
timestamp 1621261055
transform -1 0 55680 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output462
timestamp 1621261055
transform -1 0 56064 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_125
timestamp 1621261055
transform -1 0 56448 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_124
timestamp 1621261055
transform -1 0 56256 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output463
timestamp 1621261055
transform -1 0 56832 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_11_580
timestamp 1621261055
transform 1 0 56832 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_126
timestamp 1621261055
transform -1 0 57216 0 1 9990
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output464
timestamp 1621261055
transform -1 0 57600 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_11_588
timestamp 1621261055
transform 1 0 57600 0 1 9990
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_23
timestamp 1621261055
transform -1 0 58848 0 1 9990
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_11_596
timestamp 1621261055
transform 1 0 58368 0 1 9990
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_24
timestamp 1621261055
transform 1 0 1152 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_300
timestamp 1621261055
transform 1 0 3840 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_4
timestamp 1621261055
transform 1 0 1536 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_12
timestamp 1621261055
transform 1 0 2304 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_20
timestamp 1621261055
transform 1 0 3072 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_29
timestamp 1621261055
transform 1 0 3936 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _214_
timestamp 1621261055
transform -1 0 5664 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_25
timestamp 1621261055
transform -1 0 5376 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_12_37
timestamp 1621261055
transform 1 0 4704 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_12_41
timestamp 1621261055
transform 1 0 5088 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_47
timestamp 1621261055
transform 1 0 5664 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_55
timestamp 1621261055
transform 1 0 6432 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_63
timestamp 1621261055
transform 1 0 7200 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_301
timestamp 1621261055
transform 1 0 9120 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_71
timestamp 1621261055
transform 1 0 7968 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_79
timestamp 1621261055
transform 1 0 8736 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_84
timestamp 1621261055
transform 1 0 9216 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_92
timestamp 1621261055
transform 1 0 9984 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_100
timestamp 1621261055
transform 1 0 10752 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_108
timestamp 1621261055
transform 1 0 11520 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_116
timestamp 1621261055
transform 1 0 12288 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_124
timestamp 1621261055
transform 1 0 13056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_132
timestamp 1621261055
transform 1 0 13824 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_302
timestamp 1621261055
transform 1 0 14400 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_136
timestamp 1621261055
transform 1 0 14208 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_139
timestamp 1621261055
transform 1 0 14496 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_147
timestamp 1621261055
transform 1 0 15264 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_155
timestamp 1621261055
transform 1 0 16032 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_163
timestamp 1621261055
transform 1 0 16800 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_303
timestamp 1621261055
transform 1 0 19680 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_171
timestamp 1621261055
transform 1 0 17568 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_179
timestamp 1621261055
transform 1 0 18336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_187
timestamp 1621261055
transform 1 0 19104 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_191
timestamp 1621261055
transform 1 0 19488 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_194
timestamp 1621261055
transform 1 0 19776 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_202
timestamp 1621261055
transform 1 0 20544 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_210
timestamp 1621261055
transform 1 0 21312 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_218
timestamp 1621261055
transform 1 0 22080 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_226
timestamp 1621261055
transform 1 0 22848 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_304
timestamp 1621261055
transform 1 0 24960 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_234
timestamp 1621261055
transform 1 0 23616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_242
timestamp 1621261055
transform 1 0 24384 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_246
timestamp 1621261055
transform 1 0 24768 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_249
timestamp 1621261055
transform 1 0 25056 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_257
timestamp 1621261055
transform 1 0 25824 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_265
timestamp 1621261055
transform 1 0 26592 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_273
timestamp 1621261055
transform 1 0 27360 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_281
timestamp 1621261055
transform 1 0 28128 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_289
timestamp 1621261055
transform 1 0 28896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_297
timestamp 1621261055
transform 1 0 29664 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_305
timestamp 1621261055
transform 1 0 30240 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_301
timestamp 1621261055
transform 1 0 30048 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_304
timestamp 1621261055
transform 1 0 30336 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_312
timestamp 1621261055
transform 1 0 31104 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_320
timestamp 1621261055
transform 1 0 31872 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_328
timestamp 1621261055
transform 1 0 32640 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _033_
timestamp 1621261055
transform 1 0 34656 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_306
timestamp 1621261055
transform 1 0 35520 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_27
timestamp 1621261055
transform 1 0 34464 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_336
timestamp 1621261055
transform 1 0 33408 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_344
timestamp 1621261055
transform 1 0 34176 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_346
timestamp 1621261055
transform 1 0 34368 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_12_352
timestamp 1621261055
transform 1 0 34944 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_356
timestamp 1621261055
transform 1 0 35328 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_359
timestamp 1621261055
transform 1 0 35616 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_367
timestamp 1621261055
transform 1 0 36384 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_375
timestamp 1621261055
transform 1 0 37152 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_383
timestamp 1621261055
transform 1 0 37920 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_391
timestamp 1621261055
transform 1 0 38688 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_307
timestamp 1621261055
transform 1 0 40800 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_399
timestamp 1621261055
transform 1 0 39456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_407
timestamp 1621261055
transform 1 0 40224 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_411
timestamp 1621261055
transform 1 0 40608 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_414
timestamp 1621261055
transform 1 0 40896 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_422
timestamp 1621261055
transform 1 0 41664 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _062_
timestamp 1621261055
transform 1 0 42432 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_12_433
timestamp 1621261055
transform 1 0 42720 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_441
timestamp 1621261055
transform 1 0 43488 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_449
timestamp 1621261055
transform 1 0 44256 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_457
timestamp 1621261055
transform 1 0 45024 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _176_
timestamp 1621261055
transform 1 0 48192 0 -1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_308
timestamp 1621261055
transform 1 0 46080 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_465
timestamp 1621261055
transform 1 0 45792 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_12_467
timestamp 1621261055
transform 1 0 45984 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_469
timestamp 1621261055
transform 1 0 46176 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_477
timestamp 1621261055
transform 1 0 46944 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_485
timestamp 1621261055
transform 1 0 47712 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_12_489
timestamp 1621261055
transform 1 0 48096 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_493
timestamp 1621261055
transform 1 0 48480 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_309
timestamp 1621261055
transform 1 0 51360 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_12_501
timestamp 1621261055
transform 1 0 49248 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_509
timestamp 1621261055
transform 1 0 50016 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_12_517
timestamp 1621261055
transform 1 0 50784 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_521
timestamp 1621261055
transform 1 0 51168 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_12_524
timestamp 1621261055
transform 1 0 51456 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_532
timestamp 1621261055
transform 1 0 52224 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_540
timestamp 1621261055
transform 1 0 52992 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_548
timestamp 1621261055
transform 1 0 53760 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_12_556
timestamp 1621261055
transform 1 0 54528 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_568
timestamp 1621261055
transform 1 0 55680 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_12_564
timestamp 1621261055
transform 1 0 55296 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_12_574
timestamp 1621261055
transform 1 0 56256 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output470
timestamp 1621261055
transform 1 0 55872 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_310
timestamp 1621261055
transform 1 0 56640 0 -1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_12_579
timestamp 1621261055
transform 1 0 56736 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_129
timestamp 1621261055
transform -1 0 57696 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_128
timestamp 1621261055
transform -1 0 57120 0 -1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output465
timestamp 1621261055
transform -1 0 57504 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_12_589
timestamp 1621261055
transform 1 0 57696 0 -1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_25
timestamp 1621261055
transform -1 0 58848 0 -1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_26
timestamp 1621261055
transform 1 0 1152 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_4
timestamp 1621261055
transform 1 0 1536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_12
timestamp 1621261055
transform 1 0 2304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_20
timestamp 1621261055
transform 1 0 3072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_28
timestamp 1621261055
transform 1 0 3840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_311
timestamp 1621261055
transform 1 0 6432 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_53
timestamp 1621261055
transform 1 0 7488 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_36
timestamp 1621261055
transform 1 0 4608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_44
timestamp 1621261055
transform 1 0 5376 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_52
timestamp 1621261055
transform 1 0 6144 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_54
timestamp 1621261055
transform 1 0 6336 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_56
timestamp 1621261055
transform 1 0 6528 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_64
timestamp 1621261055
transform 1 0 7296 0 1 11322
box -38 -49 230 715
use HAX1  HAX1
timestamp 1623617396
transform 1 0 7680 0 1 11322
box 0 -48 3168 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_312
timestamp 1621261055
transform 1 0 11712 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_57
timestamp 1621261055
transform 1 0 10848 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_103
timestamp 1621261055
transform 1 0 11040 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_107
timestamp 1621261055
transform 1 0 11424 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_109
timestamp 1621261055
transform 1 0 11616 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_111
timestamp 1621261055
transform 1 0 11808 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_119
timestamp 1621261055
transform 1 0 12576 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_127
timestamp 1621261055
transform 1 0 13344 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_313
timestamp 1621261055
transform 1 0 16992 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_135
timestamp 1621261055
transform 1 0 14112 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_143
timestamp 1621261055
transform 1 0 14880 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_151
timestamp 1621261055
transform 1 0 15648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_159
timestamp 1621261055
transform 1 0 16416 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_163
timestamp 1621261055
transform 1 0 16800 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_166
timestamp 1621261055
transform 1 0 17088 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_174
timestamp 1621261055
transform 1 0 17856 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_182
timestamp 1621261055
transform 1 0 18624 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_190
timestamp 1621261055
transform 1 0 19392 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_198
timestamp 1621261055
transform 1 0 20160 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_314
timestamp 1621261055
transform 1 0 22272 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_206
timestamp 1621261055
transform 1 0 20928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_214
timestamp 1621261055
transform 1 0 21696 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_218
timestamp 1621261055
transform 1 0 22080 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_221
timestamp 1621261055
transform 1 0 22368 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_229
timestamp 1621261055
transform 1 0 23136 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _132_
timestamp 1621261055
transform 1 0 24864 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_13_237
timestamp 1621261055
transform 1 0 23904 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_245
timestamp 1621261055
transform 1 0 24672 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_250
timestamp 1621261055
transform 1 0 25152 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_258
timestamp 1621261055
transform 1 0 25920 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_315
timestamp 1621261055
transform 1 0 27552 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_266
timestamp 1621261055
transform 1 0 26688 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_13_274
timestamp 1621261055
transform 1 0 27456 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_276
timestamp 1621261055
transform 1 0 27648 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_284
timestamp 1621261055
transform 1 0 28416 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_292
timestamp 1621261055
transform 1 0 29184 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_316
timestamp 1621261055
transform 1 0 32832 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_300
timestamp 1621261055
transform 1 0 29952 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_308
timestamp 1621261055
transform 1 0 30720 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_316
timestamp 1621261055
transform 1 0 31488 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_324
timestamp 1621261055
transform 1 0 32256 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_328
timestamp 1621261055
transform 1 0 32640 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _028_
timestamp 1621261055
transform 1 0 34176 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_16
timestamp 1621261055
transform 1 0 33984 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_331
timestamp 1621261055
transform 1 0 32928 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_339
timestamp 1621261055
transform 1 0 33696 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_13_341
timestamp 1621261055
transform 1 0 33888 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_347
timestamp 1621261055
transform 1 0 34464 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_355
timestamp 1621261055
transform 1 0 35232 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_363
timestamp 1621261055
transform 1 0 36000 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_317
timestamp 1621261055
transform 1 0 38112 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_371
timestamp 1621261055
transform 1 0 36768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_379
timestamp 1621261055
transform 1 0 37536 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_383
timestamp 1621261055
transform 1 0 37920 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_386
timestamp 1621261055
transform 1 0 38208 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_394
timestamp 1621261055
transform 1 0 38976 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_402
timestamp 1621261055
transform 1 0 39744 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_410
timestamp 1621261055
transform 1 0 40512 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_418
timestamp 1621261055
transform 1 0 41280 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_426
timestamp 1621261055
transform 1 0 42048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _210_
timestamp 1621261055
transform 1 0 44064 0 1 11322
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_318
timestamp 1621261055
transform 1 0 43392 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_13_434
timestamp 1621261055
transform 1 0 42816 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_438
timestamp 1621261055
transform 1 0 43200 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_441
timestamp 1621261055
transform 1 0 43488 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_445
timestamp 1621261055
transform 1 0 43872 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_450
timestamp 1621261055
transform 1 0 44352 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_458
timestamp 1621261055
transform 1 0 45120 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_319
timestamp 1621261055
transform 1 0 48672 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_466
timestamp 1621261055
transform 1 0 45888 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_474
timestamp 1621261055
transform 1 0 46656 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_482
timestamp 1621261055
transform 1 0 47424 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_490
timestamp 1621261055
transform 1 0 48192 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_13_494
timestamp 1621261055
transform 1 0 48576 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_496
timestamp 1621261055
transform 1 0 48768 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_504
timestamp 1621261055
transform 1 0 49536 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_512
timestamp 1621261055
transform 1 0 50304 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_520
timestamp 1621261055
transform 1 0 51072 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_528
timestamp 1621261055
transform 1 0 51840 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_320
timestamp 1621261055
transform 1 0 53952 0 1 11322
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_13_536
timestamp 1621261055
transform 1 0 52608 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_13_544
timestamp 1621261055
transform 1 0 53376 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_548
timestamp 1621261055
transform 1 0 53760 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_13_551
timestamp 1621261055
transform 1 0 54048 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_13_559
timestamp 1621261055
transform 1 0 54816 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output467
timestamp 1621261055
transform 1 0 57120 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output474
timestamp 1621261055
transform -1 0 56736 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_142
timestamp 1621261055
transform -1 0 56352 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_567
timestamp 1621261055
transform 1 0 55584 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_571
timestamp 1621261055
transform 1 0 55968 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_13_579
timestamp 1621261055
transform 1 0 56736 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_13_587
timestamp 1621261055
transform 1 0 57504 0 1 11322
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_27
timestamp 1621261055
transform -1 0 58848 0 1 11322
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_13_595
timestamp 1621261055
transform 1 0 58272 0 1 11322
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_28
timestamp 1621261055
transform 1 0 1152 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_321
timestamp 1621261055
transform 1 0 3840 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_4
timestamp 1621261055
transform 1 0 1536 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_12
timestamp 1621261055
transform 1 0 2304 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_20
timestamp 1621261055
transform 1 0 3072 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_29
timestamp 1621261055
transform 1 0 3936 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_37
timestamp 1621261055
transform 1 0 4704 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_45
timestamp 1621261055
transform 1 0 5472 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_53
timestamp 1621261055
transform 1 0 6240 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_61
timestamp 1621261055
transform 1 0 7008 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_322
timestamp 1621261055
transform 1 0 9120 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_69
timestamp 1621261055
transform 1 0 7776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_77
timestamp 1621261055
transform 1 0 8544 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_81
timestamp 1621261055
transform 1 0 8928 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_84
timestamp 1621261055
transform 1 0 9216 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_92
timestamp 1621261055
transform 1 0 9984 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_100
timestamp 1621261055
transform 1 0 10752 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_108
timestamp 1621261055
transform 1 0 11520 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_116
timestamp 1621261055
transform 1 0 12288 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_124
timestamp 1621261055
transform 1 0 13056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_132
timestamp 1621261055
transform 1 0 13824 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_323
timestamp 1621261055
transform 1 0 14400 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_136
timestamp 1621261055
transform 1 0 14208 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_139
timestamp 1621261055
transform 1 0 14496 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_147
timestamp 1621261055
transform 1 0 15264 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_155
timestamp 1621261055
transform 1 0 16032 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_163
timestamp 1621261055
transform 1 0 16800 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_324
timestamp 1621261055
transform 1 0 19680 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_171
timestamp 1621261055
transform 1 0 17568 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_179
timestamp 1621261055
transform 1 0 18336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_187
timestamp 1621261055
transform 1 0 19104 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_191
timestamp 1621261055
transform 1 0 19488 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_194
timestamp 1621261055
transform 1 0 19776 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_202
timestamp 1621261055
transform 1 0 20544 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_210
timestamp 1621261055
transform 1 0 21312 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_218
timestamp 1621261055
transform 1 0 22080 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_226
timestamp 1621261055
transform 1 0 22848 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_325
timestamp 1621261055
transform 1 0 24960 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_234
timestamp 1621261055
transform 1 0 23616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_242
timestamp 1621261055
transform 1 0 24384 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_246
timestamp 1621261055
transform 1 0 24768 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_249
timestamp 1621261055
transform 1 0 25056 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_257
timestamp 1621261055
transform 1 0 25824 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_265
timestamp 1621261055
transform 1 0 26592 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_273
timestamp 1621261055
transform 1 0 27360 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_281
timestamp 1621261055
transform 1 0 28128 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_289
timestamp 1621261055
transform 1 0 28896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_297
timestamp 1621261055
transform 1 0 29664 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_326
timestamp 1621261055
transform 1 0 30240 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_301
timestamp 1621261055
transform 1 0 30048 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_304
timestamp 1621261055
transform 1 0 30336 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_312
timestamp 1621261055
transform 1 0 31104 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_320
timestamp 1621261055
transform 1 0 31872 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_328
timestamp 1621261055
transform 1 0 32640 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_327
timestamp 1621261055
transform 1 0 35520 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_336
timestamp 1621261055
transform 1 0 33408 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_344
timestamp 1621261055
transform 1 0 34176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_352
timestamp 1621261055
transform 1 0 34944 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_356
timestamp 1621261055
transform 1 0 35328 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_359
timestamp 1621261055
transform 1 0 35616 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _119_
timestamp 1621261055
transform 1 0 37344 0 -1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_14_367
timestamp 1621261055
transform 1 0 36384 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_375
timestamp 1621261055
transform 1 0 37152 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_380
timestamp 1621261055
transform 1 0 37632 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_388
timestamp 1621261055
transform 1 0 38400 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_396
timestamp 1621261055
transform 1 0 39168 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_328
timestamp 1621261055
transform 1 0 40800 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_404
timestamp 1621261055
transform 1 0 39936 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_14_412
timestamp 1621261055
transform 1 0 40704 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_414
timestamp 1621261055
transform 1 0 40896 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_422
timestamp 1621261055
transform 1 0 41664 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_430
timestamp 1621261055
transform 1 0 42432 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_438
timestamp 1621261055
transform 1 0 43200 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_446
timestamp 1621261055
transform 1 0 43968 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_454
timestamp 1621261055
transform 1 0 44736 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_462
timestamp 1621261055
transform 1 0 45504 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_329
timestamp 1621261055
transform 1 0 46080 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_466
timestamp 1621261055
transform 1 0 45888 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_469
timestamp 1621261055
transform 1 0 46176 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_477
timestamp 1621261055
transform 1 0 46944 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_485
timestamp 1621261055
transform 1 0 47712 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_493
timestamp 1621261055
transform 1 0 48480 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_330
timestamp 1621261055
transform 1 0 51360 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_14_501
timestamp 1621261055
transform 1 0 49248 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_509
timestamp 1621261055
transform 1 0 50016 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_14_517
timestamp 1621261055
transform 1 0 50784 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_521
timestamp 1621261055
transform 1 0 51168 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_14_524
timestamp 1621261055
transform 1 0 51456 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_532
timestamp 1621261055
transform 1 0 52224 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_540
timestamp 1621261055
transform 1 0 52992 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_548
timestamp 1621261055
transform 1 0 53760 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_556
timestamp 1621261055
transform 1 0 54528 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_14_564
timestamp 1621261055
transform 1 0 55296 0 -1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_576
timestamp 1621261055
transform 1 0 56448 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_572
timestamp 1621261055
transform 1 0 56064 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_331
timestamp 1621261055
transform 1 0 56640 0 -1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_14_583
timestamp 1621261055
transform 1 0 57120 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_14_579
timestamp 1621261055
transform 1 0 56736 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_133
timestamp 1621261055
transform -1 0 57504 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output468
timestamp 1621261055
transform -1 0 57888 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_14_593
timestamp 1621261055
transform 1 0 58080 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_134
timestamp 1621261055
transform -1 0 58080 0 -1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_29
timestamp 1621261055
transform -1 0 58848 0 -1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_4
timestamp 1621261055
transform 1 0 1536 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_4
timestamp 1621261055
transform 1 0 1536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_32
timestamp 1621261055
transform 1 0 1152 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_30
timestamp 1621261055
transform 1 0 1152 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_12
timestamp 1621261055
transform 1 0 2304 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_12
timestamp 1621261055
transform 1 0 2304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_20
timestamp 1621261055
transform 1 0 3072 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_20
timestamp 1621261055
transform 1 0 3072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_29
timestamp 1621261055
transform 1 0 3936 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_28
timestamp 1621261055
transform 1 0 3840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_342
timestamp 1621261055
transform 1 0 3840 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_37
timestamp 1621261055
transform 1 0 4704 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_36
timestamp 1621261055
transform 1 0 4608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_45
timestamp 1621261055
transform 1 0 5472 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_44
timestamp 1621261055
transform 1 0 5376 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_53
timestamp 1621261055
transform 1 0 6240 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_56
timestamp 1621261055
transform 1 0 6528 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_15_54
timestamp 1621261055
transform 1 0 6336 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_52
timestamp 1621261055
transform 1 0 6144 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_332
timestamp 1621261055
transform 1 0 6432 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_61
timestamp 1621261055
transform 1 0 7008 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_64
timestamp 1621261055
transform 1 0 7296 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_59
timestamp 1621261055
transform 1 0 7488 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_16_69
timestamp 1621261055
transform 1 0 7776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_74
timestamp 1621261055
transform 1 0 8256 0 1 12654
box -38 -49 806 715
use INV  INV
timestamp 1623617396
transform 1 0 7680 0 1 12654
box 0 -48 576 714
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_81
timestamp 1621261055
transform 1 0 8928 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_77
timestamp 1621261055
transform 1 0 8544 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_82
timestamp 1621261055
transform 1 0 9024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_343
timestamp 1621261055
transform 1 0 9120 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_92
timestamp 1621261055
transform 1 0 9984 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_84
timestamp 1621261055
transform 1 0 9216 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_90
timestamp 1621261055
transform 1 0 9792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_98
timestamp 1621261055
transform 1 0 10560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_100
timestamp 1621261055
transform 1 0 10752 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_106
timestamp 1621261055
transform 1 0 11328 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_116
timestamp 1621261055
transform 1 0 12288 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_108
timestamp 1621261055
transform 1 0 11520 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_111
timestamp 1621261055
transform 1 0 11808 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_333
timestamp 1621261055
transform 1 0 11712 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_124
timestamp 1621261055
transform 1 0 13056 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_119
timestamp 1621261055
transform 1 0 12576 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_132
timestamp 1621261055
transform 1 0 13824 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_127
timestamp 1621261055
transform 1 0 13344 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_139
timestamp 1621261055
transform 1 0 14496 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_136
timestamp 1621261055
transform 1 0 14208 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_135
timestamp 1621261055
transform 1 0 14112 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_344
timestamp 1621261055
transform 1 0 14400 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_147
timestamp 1621261055
transform 1 0 15264 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_143
timestamp 1621261055
transform 1 0 14880 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_155
timestamp 1621261055
transform 1 0 16032 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_151
timestamp 1621261055
transform 1 0 15648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_163
timestamp 1621261055
transform 1 0 16800 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_163
timestamp 1621261055
transform 1 0 16800 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_159
timestamp 1621261055
transform 1 0 16416 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_334
timestamp 1621261055
transform 1 0 16992 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_171
timestamp 1621261055
transform 1 0 17568 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_166
timestamp 1621261055
transform 1 0 17088 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_179
timestamp 1621261055
transform 1 0 18336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_182
timestamp 1621261055
transform 1 0 18624 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_174
timestamp 1621261055
transform 1 0 17856 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_191
timestamp 1621261055
transform 1 0 19488 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_187
timestamp 1621261055
transform 1 0 19104 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_190
timestamp 1621261055
transform 1 0 19392 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_194
timestamp 1621261055
transform 1 0 19776 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_198
timestamp 1621261055
transform 1 0 20160 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_345
timestamp 1621261055
transform 1 0 19680 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_202
timestamp 1621261055
transform 1 0 20544 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_206
timestamp 1621261055
transform 1 0 20928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_210
timestamp 1621261055
transform 1 0 21312 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_214
timestamp 1621261055
transform 1 0 21696 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_218
timestamp 1621261055
transform 1 0 22080 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_221
timestamp 1621261055
transform 1 0 22368 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_218
timestamp 1621261055
transform 1 0 22080 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_335
timestamp 1621261055
transform 1 0 22272 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_226
timestamp 1621261055
transform 1 0 22848 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_229
timestamp 1621261055
transform 1 0 23136 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_234
timestamp 1621261055
transform 1 0 23616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_237
timestamp 1621261055
transform 1 0 23904 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_246
timestamp 1621261055
transform 1 0 24768 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_242
timestamp 1621261055
transform 1 0 24384 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_245
timestamp 1621261055
transform 1 0 24672 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_346
timestamp 1621261055
transform 1 0 24960 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_256
timestamp 1621261055
transform 1 0 25728 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_249
timestamp 1621261055
transform 1 0 25056 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_253
timestamp 1621261055
transform 1 0 25440 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_41
timestamp 1621261055
transform -1 0 25440 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _045_
timestamp 1621261055
transform -1 0 25728 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_264
timestamp 1621261055
transform 1 0 26496 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_261
timestamp 1621261055
transform 1 0 26208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_272
timestamp 1621261055
transform 1 0 27264 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_269
timestamp 1621261055
transform 1 0 26976 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_280
timestamp 1621261055
transform 1 0 28032 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_276
timestamp 1621261055
transform 1 0 27648 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_273
timestamp 1621261055
transform 1 0 27360 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_336
timestamp 1621261055
transform 1 0 27552 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_288
timestamp 1621261055
transform 1 0 28800 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_284
timestamp 1621261055
transform 1 0 28416 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_296
timestamp 1621261055
transform 1 0 29568 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_292
timestamp 1621261055
transform 1 0 29184 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_304
timestamp 1621261055
transform 1 0 30336 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_16_302
timestamp 1621261055
transform 1 0 30144 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_300
timestamp 1621261055
transform 1 0 29952 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_300
timestamp 1621261055
transform 1 0 29952 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_347
timestamp 1621261055
transform 1 0 30240 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_312
timestamp 1621261055
transform 1 0 31104 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_308
timestamp 1621261055
transform 1 0 30720 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_320
timestamp 1621261055
transform 1 0 31872 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_316
timestamp 1621261055
transform 1 0 31488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_328
timestamp 1621261055
transform 1 0 32640 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_328
timestamp 1621261055
transform 1 0 32640 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_324
timestamp 1621261055
transform 1 0 32256 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_337
timestamp 1621261055
transform 1 0 32832 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_336
timestamp 1621261055
transform 1 0 33408 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_331
timestamp 1621261055
transform 1 0 32928 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_344
timestamp 1621261055
transform 1 0 34176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_347
timestamp 1621261055
transform 1 0 34464 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_339
timestamp 1621261055
transform 1 0 33696 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_356
timestamp 1621261055
transform 1 0 35328 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_352
timestamp 1621261055
transform 1 0 34944 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_355
timestamp 1621261055
transform 1 0 35232 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_359
timestamp 1621261055
transform 1 0 35616 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_363
timestamp 1621261055
transform 1 0 36000 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_348
timestamp 1621261055
transform 1 0 35520 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_367
timestamp 1621261055
transform 1 0 36384 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_371
timestamp 1621261055
transform 1 0 36768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_375
timestamp 1621261055
transform 1 0 37152 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_379
timestamp 1621261055
transform 1 0 37536 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_383
timestamp 1621261055
transform 1 0 37920 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_386
timestamp 1621261055
transform 1 0 38208 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_383
timestamp 1621261055
transform 1 0 37920 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_338
timestamp 1621261055
transform 1 0 38112 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_391
timestamp 1621261055
transform 1 0 38688 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_394
timestamp 1621261055
transform 1 0 38976 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_399
timestamp 1621261055
transform 1 0 39456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_402
timestamp 1621261055
transform 1 0 39744 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_411
timestamp 1621261055
transform 1 0 40608 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_407
timestamp 1621261055
transform 1 0 40224 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_410
timestamp 1621261055
transform 1 0 40512 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_349
timestamp 1621261055
transform 1 0 40800 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_422
timestamp 1621261055
transform 1 0 41664 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_414
timestamp 1621261055
transform 1 0 40896 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_418
timestamp 1621261055
transform 1 0 41280 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_426
timestamp 1621261055
transform 1 0 42048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_430
timestamp 1621261055
transform 1 0 42432 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_434
timestamp 1621261055
transform 1 0 42816 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_16_446
timestamp 1621261055
transform 1 0 43968 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_438
timestamp 1621261055
transform 1 0 43200 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_441
timestamp 1621261055
transform 1 0 43488 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_438
timestamp 1621261055
transform 1 0 43200 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_339
timestamp 1621261055
transform 1 0 43392 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_454
timestamp 1621261055
transform 1 0 44736 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_449
timestamp 1621261055
transform 1 0 44256 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_16_462
timestamp 1621261055
transform 1 0 45504 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_457
timestamp 1621261055
transform 1 0 45024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_469
timestamp 1621261055
transform 1 0 46176 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_466
timestamp 1621261055
transform 1 0 45888 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_15_465
timestamp 1621261055
transform 1 0 45792 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_350
timestamp 1621261055
transform 1 0 46080 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_477
timestamp 1621261055
transform 1 0 46944 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_473
timestamp 1621261055
transform 1 0 46560 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_485
timestamp 1621261055
transform 1 0 47712 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_481
timestamp 1621261055
transform 1 0 47328 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_493
timestamp 1621261055
transform 1 0 48480 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_493
timestamp 1621261055
transform 1 0 48480 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_489
timestamp 1621261055
transform 1 0 48096 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_340
timestamp 1621261055
transform 1 0 48672 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_501
timestamp 1621261055
transform 1 0 49248 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_496
timestamp 1621261055
transform 1 0 48768 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_509
timestamp 1621261055
transform 1 0 50016 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_512
timestamp 1621261055
transform 1 0 50304 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_504
timestamp 1621261055
transform 1 0 49536 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_521
timestamp 1621261055
transform 1 0 51168 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_517
timestamp 1621261055
transform 1 0 50784 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_520
timestamp 1621261055
transform 1 0 51072 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_524
timestamp 1621261055
transform 1 0 51456 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_528
timestamp 1621261055
transform 1 0 51840 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_351
timestamp 1621261055
transform 1 0 51360 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_16_532
timestamp 1621261055
transform 1 0 52224 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_536
timestamp 1621261055
transform 1 0 52608 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_540
timestamp 1621261055
transform 1 0 52992 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_15_544
timestamp 1621261055
transform 1 0 53376 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_16_552
timestamp 1621261055
transform 1 0 54144 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_16_548
timestamp 1621261055
transform 1 0 53760 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_551
timestamp 1621261055
transform 1 0 54048 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_548
timestamp 1621261055
transform 1 0 53760 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_341
timestamp 1621261055
transform 1 0 53952 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _105_
timestamp 1621261055
transform 1 0 54240 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_556
timestamp 1621261055
transform 1 0 54528 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_559
timestamp 1621261055
transform 1 0 54816 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_16_564
timestamp 1621261055
transform 1 0 55296 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_15_567
timestamp 1621261055
transform 1 0 55584 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_576
timestamp 1621261055
transform 1 0 56448 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_572
timestamp 1621261055
transform 1 0 56064 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_575
timestamp 1621261055
transform 1 0 56352 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_81
timestamp 1621261055
transform -1 0 56736 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_352
timestamp 1621261055
transform 1 0 56640 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_16_583
timestamp 1621261055
transform 1 0 57120 0 -1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_16_579
timestamp 1621261055
transform 1 0 56736 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_15_582
timestamp 1621261055
transform 1 0 57024 0 1 12654
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _161_
timestamp 1621261055
transform 1 0 57312 0 -1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _057_
timestamp 1621261055
transform -1 0 57024 0 1 12654
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_16_588
timestamp 1621261055
transform 1 0 57600 0 -1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_15_594
timestamp 1621261055
transform 1 0 58176 0 1 12654
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_15_590
timestamp 1621261055
transform 1 0 57792 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_31
timestamp 1621261055
transform -1 0 58848 0 1 12654
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_33
timestamp 1621261055
transform -1 0 58848 0 -1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_15_596
timestamp 1621261055
transform 1 0 58368 0 1 12654
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_16_596
timestamp 1621261055
transform 1 0 58368 0 -1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_34
timestamp 1621261055
transform 1 0 1152 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_4
timestamp 1621261055
transform 1 0 1536 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_12
timestamp 1621261055
transform 1 0 2304 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_20
timestamp 1621261055
transform 1 0 3072 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_28
timestamp 1621261055
transform 1 0 3840 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_353
timestamp 1621261055
transform 1 0 6432 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_63
timestamp 1621261055
transform 1 0 7488 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_36
timestamp 1621261055
transform 1 0 4608 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_44
timestamp 1621261055
transform 1 0 5376 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_52
timestamp 1621261055
transform 1 0 6144 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_54
timestamp 1621261055
transform 1 0 6336 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_56
timestamp 1621261055
transform 1 0 6528 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_64
timestamp 1621261055
transform 1 0 7296 0 1 13986
box -38 -49 230 715
use INVX1  INVX1
timestamp 1623617396
transform 1 0 7680 0 1 13986
box 0 -48 576 714
use sky130_fd_sc_ls__conb_1  _108_
timestamp 1621261055
transform 1 0 9408 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_17_74
timestamp 1621261055
transform 1 0 8256 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_82
timestamp 1621261055
transform 1 0 9024 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_17_89
timestamp 1621261055
transform 1 0 9696 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_97
timestamp 1621261055
transform 1 0 10464 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_354
timestamp 1621261055
transform 1 0 11712 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_105
timestamp 1621261055
transform 1 0 11232 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_17_109
timestamp 1621261055
transform 1 0 11616 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_111
timestamp 1621261055
transform 1 0 11808 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_119
timestamp 1621261055
transform 1 0 12576 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_127
timestamp 1621261055
transform 1 0 13344 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _130_
timestamp 1621261055
transform 1 0 14400 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_355
timestamp 1621261055
transform 1 0 16992 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_135
timestamp 1621261055
transform 1 0 14112 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_137
timestamp 1621261055
transform 1 0 14304 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_141
timestamp 1621261055
transform 1 0 14688 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_149
timestamp 1621261055
transform 1 0 15456 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_157
timestamp 1621261055
transform 1 0 16224 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_166
timestamp 1621261055
transform 1 0 17088 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_174
timestamp 1621261055
transform 1 0 17856 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_182
timestamp 1621261055
transform 1 0 18624 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_190
timestamp 1621261055
transform 1 0 19392 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_198
timestamp 1621261055
transform 1 0 20160 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_356
timestamp 1621261055
transform 1 0 22272 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_206
timestamp 1621261055
transform 1 0 20928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_214
timestamp 1621261055
transform 1 0 21696 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_218
timestamp 1621261055
transform 1 0 22080 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_221
timestamp 1621261055
transform 1 0 22368 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_229
timestamp 1621261055
transform 1 0 23136 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_237
timestamp 1621261055
transform 1 0 23904 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_245
timestamp 1621261055
transform 1 0 24672 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_253
timestamp 1621261055
transform 1 0 25440 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_261
timestamp 1621261055
transform 1 0 26208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _023_
timestamp 1621261055
transform 1 0 28032 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_357
timestamp 1621261055
transform 1 0 27552 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_0
timestamp 1621261055
transform 1 0 27840 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_17_269
timestamp 1621261055
transform 1 0 26976 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_273
timestamp 1621261055
transform 1 0 27360 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_276
timestamp 1621261055
transform 1 0 27648 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_283
timestamp 1621261055
transform 1 0 28320 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_291
timestamp 1621261055
transform 1 0 29088 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_358
timestamp 1621261055
transform 1 0 32832 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_299
timestamp 1621261055
transform 1 0 29856 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_307
timestamp 1621261055
transform 1 0 30624 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_315
timestamp 1621261055
transform 1 0 31392 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_323
timestamp 1621261055
transform 1 0 32160 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_327
timestamp 1621261055
transform 1 0 32544 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_17_329
timestamp 1621261055
transform 1 0 32736 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_331
timestamp 1621261055
transform 1 0 32928 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_339
timestamp 1621261055
transform 1 0 33696 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_347
timestamp 1621261055
transform 1 0 34464 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_355
timestamp 1621261055
transform 1 0 35232 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_363
timestamp 1621261055
transform 1 0 36000 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_359
timestamp 1621261055
transform 1 0 38112 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_371
timestamp 1621261055
transform 1 0 36768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_379
timestamp 1621261055
transform 1 0 37536 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_383
timestamp 1621261055
transform 1 0 37920 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_386
timestamp 1621261055
transform 1 0 38208 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_394
timestamp 1621261055
transform 1 0 38976 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_402
timestamp 1621261055
transform 1 0 39744 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_410
timestamp 1621261055
transform 1 0 40512 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_418
timestamp 1621261055
transform 1 0 41280 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_426
timestamp 1621261055
transform 1 0 42048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_360
timestamp 1621261055
transform 1 0 43392 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_17_434
timestamp 1621261055
transform 1 0 42816 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_438
timestamp 1621261055
transform 1 0 43200 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_441
timestamp 1621261055
transform 1 0 43488 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_449
timestamp 1621261055
transform 1 0 44256 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_457
timestamp 1621261055
transform 1 0 45024 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_361
timestamp 1621261055
transform 1 0 48672 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_465
timestamp 1621261055
transform 1 0 45792 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_473
timestamp 1621261055
transform 1 0 46560 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_481
timestamp 1621261055
transform 1 0 47328 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_489
timestamp 1621261055
transform 1 0 48096 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_493
timestamp 1621261055
transform 1 0 48480 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _216_
timestamp 1621261055
transform 1 0 49632 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_17_496
timestamp 1621261055
transform 1 0 48768 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_17_504
timestamp 1621261055
transform 1 0 49536 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_508
timestamp 1621261055
transform 1 0 49920 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_516
timestamp 1621261055
transform 1 0 50688 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_524
timestamp 1621261055
transform 1 0 51456 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_362
timestamp 1621261055
transform 1 0 53952 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_17_532
timestamp 1621261055
transform 1 0 52224 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_540
timestamp 1621261055
transform 1 0 52992 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_548
timestamp 1621261055
transform 1 0 53760 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_551
timestamp 1621261055
transform 1 0 54048 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_559
timestamp 1621261055
transform 1 0 54816 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _175_
timestamp 1621261055
transform 1 0 56160 0 1 13986
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_17_567
timestamp 1621261055
transform 1 0 55584 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_17_571
timestamp 1621261055
transform 1 0 55968 0 1 13986
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_17_576
timestamp 1621261055
transform 1 0 56448 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_17_584
timestamp 1621261055
transform 1 0 57216 0 1 13986
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_17_592
timestamp 1621261055
transform 1 0 57984 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_35
timestamp 1621261055
transform -1 0 58848 0 1 13986
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_17_596
timestamp 1621261055
transform 1 0 58368 0 1 13986
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _003_
timestamp 1621261055
transform -1 0 2784 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_36
timestamp 1621261055
transform 1 0 1152 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_363
timestamp 1621261055
transform 1 0 3840 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_10
timestamp 1621261055
transform -1 0 2496 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_4
timestamp 1621261055
transform 1 0 1536 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_17
timestamp 1621261055
transform 1 0 2784 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_25
timestamp 1621261055
transform 1 0 3552 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_27
timestamp 1621261055
transform 1 0 3744 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_29
timestamp 1621261055
transform 1 0 3936 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_37
timestamp 1621261055
transform 1 0 4704 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_45
timestamp 1621261055
transform 1 0 5472 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_53
timestamp 1621261055
transform 1 0 6240 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_61
timestamp 1621261055
transform 1 0 7008 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_364
timestamp 1621261055
transform 1 0 9120 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_69
timestamp 1621261055
transform 1 0 7776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_77
timestamp 1621261055
transform 1 0 8544 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_81
timestamp 1621261055
transform 1 0 8928 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_84
timestamp 1621261055
transform 1 0 9216 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_92
timestamp 1621261055
transform 1 0 9984 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_100
timestamp 1621261055
transform 1 0 10752 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_108
timestamp 1621261055
transform 1 0 11520 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_116
timestamp 1621261055
transform 1 0 12288 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_124
timestamp 1621261055
transform 1 0 13056 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_132
timestamp 1621261055
transform 1 0 13824 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_365
timestamp 1621261055
transform 1 0 14400 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_136
timestamp 1621261055
transform 1 0 14208 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_139
timestamp 1621261055
transform 1 0 14496 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_147
timestamp 1621261055
transform 1 0 15264 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_155
timestamp 1621261055
transform 1 0 16032 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_163
timestamp 1621261055
transform 1 0 16800 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_366
timestamp 1621261055
transform 1 0 19680 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_171
timestamp 1621261055
transform 1 0 17568 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_179
timestamp 1621261055
transform 1 0 18336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_187
timestamp 1621261055
transform 1 0 19104 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_191
timestamp 1621261055
transform 1 0 19488 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_194
timestamp 1621261055
transform 1 0 19776 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_202
timestamp 1621261055
transform 1 0 20544 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_210
timestamp 1621261055
transform 1 0 21312 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_218
timestamp 1621261055
transform 1 0 22080 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_226
timestamp 1621261055
transform 1 0 22848 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _091_
timestamp 1621261055
transform 1 0 25440 0 -1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_367
timestamp 1621261055
transform 1 0 24960 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_234
timestamp 1621261055
transform 1 0 23616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_242
timestamp 1621261055
transform 1 0 24384 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_246
timestamp 1621261055
transform 1 0 24768 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_18_249
timestamp 1621261055
transform 1 0 25056 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_18_256
timestamp 1621261055
transform 1 0 25728 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_264
timestamp 1621261055
transform 1 0 26496 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_272
timestamp 1621261055
transform 1 0 27264 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_280
timestamp 1621261055
transform 1 0 28032 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_288
timestamp 1621261055
transform 1 0 28800 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_296
timestamp 1621261055
transform 1 0 29568 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_368
timestamp 1621261055
transform 1 0 30240 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_300
timestamp 1621261055
transform 1 0 29952 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_18_302
timestamp 1621261055
transform 1 0 30144 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_304
timestamp 1621261055
transform 1 0 30336 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_312
timestamp 1621261055
transform 1 0 31104 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_320
timestamp 1621261055
transform 1 0 31872 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_328
timestamp 1621261055
transform 1 0 32640 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_369
timestamp 1621261055
transform 1 0 35520 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_336
timestamp 1621261055
transform 1 0 33408 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_344
timestamp 1621261055
transform 1 0 34176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_352
timestamp 1621261055
transform 1 0 34944 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_356
timestamp 1621261055
transform 1 0 35328 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_359
timestamp 1621261055
transform 1 0 35616 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_367
timestamp 1621261055
transform 1 0 36384 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_375
timestamp 1621261055
transform 1 0 37152 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_383
timestamp 1621261055
transform 1 0 37920 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_391
timestamp 1621261055
transform 1 0 38688 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_370
timestamp 1621261055
transform 1 0 40800 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_399
timestamp 1621261055
transform 1 0 39456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_407
timestamp 1621261055
transform 1 0 40224 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_411
timestamp 1621261055
transform 1 0 40608 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_414
timestamp 1621261055
transform 1 0 40896 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_422
timestamp 1621261055
transform 1 0 41664 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_430
timestamp 1621261055
transform 1 0 42432 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_438
timestamp 1621261055
transform 1 0 43200 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_446
timestamp 1621261055
transform 1 0 43968 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_454
timestamp 1621261055
transform 1 0 44736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_462
timestamp 1621261055
transform 1 0 45504 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_371
timestamp 1621261055
transform 1 0 46080 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_466
timestamp 1621261055
transform 1 0 45888 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_469
timestamp 1621261055
transform 1 0 46176 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_477
timestamp 1621261055
transform 1 0 46944 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_485
timestamp 1621261055
transform 1 0 47712 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_493
timestamp 1621261055
transform 1 0 48480 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_372
timestamp 1621261055
transform 1 0 51360 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_501
timestamp 1621261055
transform 1 0 49248 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_509
timestamp 1621261055
transform 1 0 50016 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_517
timestamp 1621261055
transform 1 0 50784 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_521
timestamp 1621261055
transform 1 0 51168 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_524
timestamp 1621261055
transform 1 0 51456 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_532
timestamp 1621261055
transform 1 0 52224 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_540
timestamp 1621261055
transform 1 0 52992 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_548
timestamp 1621261055
transform 1 0 53760 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_556
timestamp 1621261055
transform 1 0 54528 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_373
timestamp 1621261055
transform 1 0 56640 0 -1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_18_564
timestamp 1621261055
transform 1 0 55296 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_18_572
timestamp 1621261055
transform 1 0 56064 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_576
timestamp 1621261055
transform 1 0 56448 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_18_579
timestamp 1621261055
transform 1 0 56736 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_18_587
timestamp 1621261055
transform 1 0 57504 0 -1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_37
timestamp 1621261055
transform -1 0 58848 0 -1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_18_595
timestamp 1621261055
transform 1 0 58272 0 -1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _061_
timestamp 1621261055
transform 1 0 3648 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_38
timestamp 1621261055
transform 1 0 1152 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_4
timestamp 1621261055
transform 1 0 1536 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_12
timestamp 1621261055
transform 1 0 2304 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_20
timestamp 1621261055
transform 1 0 3072 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_24
timestamp 1621261055
transform 1 0 3456 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_29
timestamp 1621261055
transform 1 0 3936 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_374
timestamp 1621261055
transform 1 0 6432 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_65
timestamp 1621261055
transform 1 0 7488 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_37
timestamp 1621261055
transform 1 0 4704 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_45
timestamp 1621261055
transform 1 0 5472 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_53
timestamp 1621261055
transform 1 0 6240 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_56
timestamp 1621261055
transform 1 0 6528 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_64
timestamp 1621261055
transform 1 0 7296 0 1 15318
box -38 -49 230 715
use INVX2  INVX2
timestamp 1623617396
transform 1 0 7680 0 1 15318
box 0 -48 576 714
use sky130_fd_sc_ls__conb_1  _164_
timestamp 1621261055
transform 1 0 8640 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_19_74
timestamp 1621261055
transform 1 0 8256 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_81
timestamp 1621261055
transform 1 0 8928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_89
timestamp 1621261055
transform 1 0 9696 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_97
timestamp 1621261055
transform 1 0 10464 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_375
timestamp 1621261055
transform 1 0 11712 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_105
timestamp 1621261055
transform 1 0 11232 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_19_109
timestamp 1621261055
transform 1 0 11616 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_111
timestamp 1621261055
transform 1 0 11808 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_119
timestamp 1621261055
transform 1 0 12576 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_127
timestamp 1621261055
transform 1 0 13344 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _151_
timestamp 1621261055
transform 1 0 15936 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_376
timestamp 1621261055
transform 1 0 16992 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_135
timestamp 1621261055
transform 1 0 14112 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_143
timestamp 1621261055
transform 1 0 14880 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_151
timestamp 1621261055
transform 1 0 15648 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_153
timestamp 1621261055
transform 1 0 15840 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_157
timestamp 1621261055
transform 1 0 16224 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_166
timestamp 1621261055
transform 1 0 17088 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_174
timestamp 1621261055
transform 1 0 17856 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_182
timestamp 1621261055
transform 1 0 18624 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_190
timestamp 1621261055
transform 1 0 19392 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_198
timestamp 1621261055
transform 1 0 20160 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_377
timestamp 1621261055
transform 1 0 22272 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_206
timestamp 1621261055
transform 1 0 20928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_214
timestamp 1621261055
transform 1 0 21696 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_218
timestamp 1621261055
transform 1 0 22080 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_221
timestamp 1621261055
transform 1 0 22368 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_229
timestamp 1621261055
transform 1 0 23136 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_237
timestamp 1621261055
transform 1 0 23904 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_245
timestamp 1621261055
transform 1 0 24672 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_253
timestamp 1621261055
transform 1 0 25440 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_261
timestamp 1621261055
transform 1 0 26208 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _149_
timestamp 1621261055
transform 1 0 26592 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_378
timestamp 1621261055
transform 1 0 27552 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_268
timestamp 1621261055
transform 1 0 26880 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_272
timestamp 1621261055
transform 1 0 27264 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_274
timestamp 1621261055
transform 1 0 27456 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_276
timestamp 1621261055
transform 1 0 27648 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_284
timestamp 1621261055
transform 1 0 28416 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_292
timestamp 1621261055
transform 1 0 29184 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_379
timestamp 1621261055
transform 1 0 32832 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_300
timestamp 1621261055
transform 1 0 29952 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_308
timestamp 1621261055
transform 1 0 30720 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_316
timestamp 1621261055
transform 1 0 31488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_324
timestamp 1621261055
transform 1 0 32256 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_328
timestamp 1621261055
transform 1 0 32640 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_331
timestamp 1621261055
transform 1 0 32928 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_339
timestamp 1621261055
transform 1 0 33696 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_347
timestamp 1621261055
transform 1 0 34464 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_355
timestamp 1621261055
transform 1 0 35232 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_363
timestamp 1621261055
transform 1 0 36000 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_380
timestamp 1621261055
transform 1 0 38112 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_371
timestamp 1621261055
transform 1 0 36768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_379
timestamp 1621261055
transform 1 0 37536 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_383
timestamp 1621261055
transform 1 0 37920 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_386
timestamp 1621261055
transform 1 0 38208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_394
timestamp 1621261055
transform 1 0 38976 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_402
timestamp 1621261055
transform 1 0 39744 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_410
timestamp 1621261055
transform 1 0 40512 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_418
timestamp 1621261055
transform 1 0 41280 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_426
timestamp 1621261055
transform 1 0 42048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_381
timestamp 1621261055
transform 1 0 43392 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_19_434
timestamp 1621261055
transform 1 0 42816 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_438
timestamp 1621261055
transform 1 0 43200 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_19_441
timestamp 1621261055
transform 1 0 43488 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_449
timestamp 1621261055
transform 1 0 44256 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_457
timestamp 1621261055
transform 1 0 45024 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_382
timestamp 1621261055
transform 1 0 48672 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_465
timestamp 1621261055
transform 1 0 45792 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_473
timestamp 1621261055
transform 1 0 46560 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_481
timestamp 1621261055
transform 1 0 47328 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_489
timestamp 1621261055
transform 1 0 48096 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_493
timestamp 1621261055
transform 1 0 48480 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _148_
timestamp 1621261055
transform 1 0 49920 0 1 15318
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_19_496
timestamp 1621261055
transform 1 0 48768 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_504
timestamp 1621261055
transform 1 0 49536 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_19_511
timestamp 1621261055
transform 1 0 50208 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_519
timestamp 1621261055
transform 1 0 50976 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_527
timestamp 1621261055
transform 1 0 51744 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_383
timestamp 1621261055
transform 1 0 53952 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_535
timestamp 1621261055
transform 1 0 52512 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_543
timestamp 1621261055
transform 1 0 53280 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_547
timestamp 1621261055
transform 1 0 53664 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_19_549
timestamp 1621261055
transform 1 0 53856 0 1 15318
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_19_551
timestamp 1621261055
transform 1 0 54048 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_559
timestamp 1621261055
transform 1 0 54816 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_567
timestamp 1621261055
transform 1 0 55584 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_575
timestamp 1621261055
transform 1 0 56352 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_19_583
timestamp 1621261055
transform 1 0 57120 0 1 15318
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_19_591
timestamp 1621261055
transform 1 0 57888 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_39
timestamp 1621261055
transform -1 0 58848 0 1 15318
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_19_595
timestamp 1621261055
transform 1 0 58272 0 1 15318
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_8
timestamp 1621261055
transform 1 0 1920 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_20_4
timestamp 1621261055
transform 1 0 1536 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_40
timestamp 1621261055
transform 1 0 1152 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_20_16
timestamp 1621261055
transform 1 0 2688 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_20_10
timestamp 1621261055
transform 1 0 2112 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_33
timestamp 1621261055
transform -1 0 2400 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _019_
timestamp 1621261055
transform -1 0 2688 0 -1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_20_24
timestamp 1621261055
transform 1 0 3456 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_20_29
timestamp 1621261055
transform 1 0 3936 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_384
timestamp 1621261055
transform 1 0 3840 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_37
timestamp 1621261055
transform 1 0 4704 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_45
timestamp 1621261055
transform 1 0 5472 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_53
timestamp 1621261055
transform 1 0 6240 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_61
timestamp 1621261055
transform 1 0 7008 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_385
timestamp 1621261055
transform 1 0 9120 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_69
timestamp 1621261055
transform 1 0 7776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_77
timestamp 1621261055
transform 1 0 8544 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_81
timestamp 1621261055
transform 1 0 8928 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_84
timestamp 1621261055
transform 1 0 9216 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_92
timestamp 1621261055
transform 1 0 9984 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_100
timestamp 1621261055
transform 1 0 10752 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_108
timestamp 1621261055
transform 1 0 11520 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_116
timestamp 1621261055
transform 1 0 12288 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_124
timestamp 1621261055
transform 1 0 13056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_132
timestamp 1621261055
transform 1 0 13824 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_386
timestamp 1621261055
transform 1 0 14400 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_136
timestamp 1621261055
transform 1 0 14208 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_139
timestamp 1621261055
transform 1 0 14496 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_147
timestamp 1621261055
transform 1 0 15264 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_155
timestamp 1621261055
transform 1 0 16032 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_163
timestamp 1621261055
transform 1 0 16800 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_387
timestamp 1621261055
transform 1 0 19680 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_171
timestamp 1621261055
transform 1 0 17568 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_179
timestamp 1621261055
transform 1 0 18336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_187
timestamp 1621261055
transform 1 0 19104 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_191
timestamp 1621261055
transform 1 0 19488 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_194
timestamp 1621261055
transform 1 0 19776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_202
timestamp 1621261055
transform 1 0 20544 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_210
timestamp 1621261055
transform 1 0 21312 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_218
timestamp 1621261055
transform 1 0 22080 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_226
timestamp 1621261055
transform 1 0 22848 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_388
timestamp 1621261055
transform 1 0 24960 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_234
timestamp 1621261055
transform 1 0 23616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_242
timestamp 1621261055
transform 1 0 24384 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_246
timestamp 1621261055
transform 1 0 24768 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_249
timestamp 1621261055
transform 1 0 25056 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_257
timestamp 1621261055
transform 1 0 25824 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_265
timestamp 1621261055
transform 1 0 26592 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_273
timestamp 1621261055
transform 1 0 27360 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_281
timestamp 1621261055
transform 1 0 28128 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_289
timestamp 1621261055
transform 1 0 28896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_297
timestamp 1621261055
transform 1 0 29664 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_389
timestamp 1621261055
transform 1 0 30240 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_301
timestamp 1621261055
transform 1 0 30048 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_304
timestamp 1621261055
transform 1 0 30336 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_312
timestamp 1621261055
transform 1 0 31104 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_320
timestamp 1621261055
transform 1 0 31872 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_328
timestamp 1621261055
transform 1 0 32640 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_390
timestamp 1621261055
transform 1 0 35520 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_336
timestamp 1621261055
transform 1 0 33408 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_344
timestamp 1621261055
transform 1 0 34176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_352
timestamp 1621261055
transform 1 0 34944 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_356
timestamp 1621261055
transform 1 0 35328 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_359
timestamp 1621261055
transform 1 0 35616 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_367
timestamp 1621261055
transform 1 0 36384 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_375
timestamp 1621261055
transform 1 0 37152 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_383
timestamp 1621261055
transform 1 0 37920 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_391
timestamp 1621261055
transform 1 0 38688 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_391
timestamp 1621261055
transform 1 0 40800 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_399
timestamp 1621261055
transform 1 0 39456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_407
timestamp 1621261055
transform 1 0 40224 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_411
timestamp 1621261055
transform 1 0 40608 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_414
timestamp 1621261055
transform 1 0 40896 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_422
timestamp 1621261055
transform 1 0 41664 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_430
timestamp 1621261055
transform 1 0 42432 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_438
timestamp 1621261055
transform 1 0 43200 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_446
timestamp 1621261055
transform 1 0 43968 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_454
timestamp 1621261055
transform 1 0 44736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_462
timestamp 1621261055
transform 1 0 45504 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_392
timestamp 1621261055
transform 1 0 46080 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_466
timestamp 1621261055
transform 1 0 45888 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_469
timestamp 1621261055
transform 1 0 46176 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_477
timestamp 1621261055
transform 1 0 46944 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_485
timestamp 1621261055
transform 1 0 47712 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_493
timestamp 1621261055
transform 1 0 48480 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_393
timestamp 1621261055
transform 1 0 51360 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_501
timestamp 1621261055
transform 1 0 49248 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_509
timestamp 1621261055
transform 1 0 50016 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_20_517
timestamp 1621261055
transform 1 0 50784 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_521
timestamp 1621261055
transform 1 0 51168 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_524
timestamp 1621261055
transform 1 0 51456 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _181_
timestamp 1621261055
transform 1 0 53952 0 -1 16650
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_20_532
timestamp 1621261055
transform 1 0 52224 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_540
timestamp 1621261055
transform 1 0 52992 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_548
timestamp 1621261055
transform 1 0 53760 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_20_553
timestamp 1621261055
transform 1 0 54240 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_561
timestamp 1621261055
transform 1 0 55008 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_394
timestamp 1621261055
transform 1 0 56640 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_569
timestamp 1621261055
transform 1 0 55776 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_20_577
timestamp 1621261055
transform 1 0 56544 0 -1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_20_579
timestamp 1621261055
transform 1 0 56736 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_20_587
timestamp 1621261055
transform 1 0 57504 0 -1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_41
timestamp 1621261055
transform -1 0 58848 0 -1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_20_595
timestamp 1621261055
transform 1 0 58272 0 -1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_42
timestamp 1621261055
transform 1 0 1152 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_21_4
timestamp 1621261055
transform 1 0 1536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_12
timestamp 1621261055
transform 1 0 2304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_20
timestamp 1621261055
transform 1 0 3072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_28
timestamp 1621261055
transform 1 0 3840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_395
timestamp 1621261055
transform 1 0 6432 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_67
timestamp 1621261055
transform 1 0 7488 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_36
timestamp 1621261055
transform 1 0 4608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_44
timestamp 1621261055
transform 1 0 5376 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_52
timestamp 1621261055
transform 1 0 6144 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_21_54
timestamp 1621261055
transform 1 0 6336 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_56
timestamp 1621261055
transform 1 0 6528 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_64
timestamp 1621261055
transform 1 0 7296 0 1 16650
box -38 -49 230 715
use INVX4  INVX4
timestamp 1623617396
transform 1 0 7680 0 1 16650
box 0 -48 864 714
use sky130_fd_sc_ls__decap_8  FILLER_21_77
timestamp 1621261055
transform 1 0 8544 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_85
timestamp 1621261055
transform 1 0 9312 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_93
timestamp 1621261055
transform 1 0 10080 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_396
timestamp 1621261055
transform 1 0 11712 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_101
timestamp 1621261055
transform 1 0 10848 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_21_109
timestamp 1621261055
transform 1 0 11616 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_111
timestamp 1621261055
transform 1 0 11808 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_119
timestamp 1621261055
transform 1 0 12576 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_127
timestamp 1621261055
transform 1 0 13344 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_397
timestamp 1621261055
transform 1 0 16992 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_135
timestamp 1621261055
transform 1 0 14112 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_143
timestamp 1621261055
transform 1 0 14880 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_151
timestamp 1621261055
transform 1 0 15648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_159
timestamp 1621261055
transform 1 0 16416 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_163
timestamp 1621261055
transform 1 0 16800 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_166
timestamp 1621261055
transform 1 0 17088 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_174
timestamp 1621261055
transform 1 0 17856 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_182
timestamp 1621261055
transform 1 0 18624 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_190
timestamp 1621261055
transform 1 0 19392 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_198
timestamp 1621261055
transform 1 0 20160 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_398
timestamp 1621261055
transform 1 0 22272 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_206
timestamp 1621261055
transform 1 0 20928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_214
timestamp 1621261055
transform 1 0 21696 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_218
timestamp 1621261055
transform 1 0 22080 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_221
timestamp 1621261055
transform 1 0 22368 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_229
timestamp 1621261055
transform 1 0 23136 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_237
timestamp 1621261055
transform 1 0 23904 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_245
timestamp 1621261055
transform 1 0 24672 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_253
timestamp 1621261055
transform 1 0 25440 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_261
timestamp 1621261055
transform 1 0 26208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_399
timestamp 1621261055
transform 1 0 27552 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_269
timestamp 1621261055
transform 1 0 26976 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_273
timestamp 1621261055
transform 1 0 27360 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_276
timestamp 1621261055
transform 1 0 27648 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_284
timestamp 1621261055
transform 1 0 28416 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_292
timestamp 1621261055
transform 1 0 29184 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_400
timestamp 1621261055
transform 1 0 32832 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_300
timestamp 1621261055
transform 1 0 29952 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_308
timestamp 1621261055
transform 1 0 30720 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_316
timestamp 1621261055
transform 1 0 31488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_324
timestamp 1621261055
transform 1 0 32256 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_328
timestamp 1621261055
transform 1 0 32640 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_331
timestamp 1621261055
transform 1 0 32928 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_339
timestamp 1621261055
transform 1 0 33696 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_347
timestamp 1621261055
transform 1 0 34464 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_355
timestamp 1621261055
transform 1 0 35232 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_363
timestamp 1621261055
transform 1 0 36000 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_401
timestamp 1621261055
transform 1 0 38112 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_371
timestamp 1621261055
transform 1 0 36768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_379
timestamp 1621261055
transform 1 0 37536 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_383
timestamp 1621261055
transform 1 0 37920 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_386
timestamp 1621261055
transform 1 0 38208 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_394
timestamp 1621261055
transform 1 0 38976 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_402
timestamp 1621261055
transform 1 0 39744 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_410
timestamp 1621261055
transform 1 0 40512 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_418
timestamp 1621261055
transform 1 0 41280 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_426
timestamp 1621261055
transform 1 0 42048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_402
timestamp 1621261055
transform 1 0 43392 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_21_434
timestamp 1621261055
transform 1 0 42816 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_438
timestamp 1621261055
transform 1 0 43200 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_441
timestamp 1621261055
transform 1 0 43488 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_449
timestamp 1621261055
transform 1 0 44256 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_457
timestamp 1621261055
transform 1 0 45024 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_403
timestamp 1621261055
transform 1 0 48672 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_465
timestamp 1621261055
transform 1 0 45792 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_473
timestamp 1621261055
transform 1 0 46560 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_481
timestamp 1621261055
transform 1 0 47328 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_489
timestamp 1621261055
transform 1 0 48096 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_493
timestamp 1621261055
transform 1 0 48480 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_496
timestamp 1621261055
transform 1 0 48768 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_504
timestamp 1621261055
transform 1 0 49536 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_512
timestamp 1621261055
transform 1 0 50304 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_520
timestamp 1621261055
transform 1 0 51072 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_528
timestamp 1621261055
transform 1 0 51840 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_404
timestamp 1621261055
transform 1 0 53952 0 1 16650
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_21_536
timestamp 1621261055
transform 1 0 52608 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_544
timestamp 1621261055
transform 1 0 53376 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_548
timestamp 1621261055
transform 1 0 53760 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_21_551
timestamp 1621261055
transform 1 0 54048 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_559
timestamp 1621261055
transform 1 0 54816 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_567
timestamp 1621261055
transform 1 0 55584 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_575
timestamp 1621261055
transform 1 0 56352 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_21_583
timestamp 1621261055
transform 1 0 57120 0 1 16650
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_21_591
timestamp 1621261055
transform 1 0 57888 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_43
timestamp 1621261055
transform -1 0 58848 0 1 16650
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_21_595
timestamp 1621261055
transform 1 0 58272 0 1 16650
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_44
timestamp 1621261055
transform 1 0 1152 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_405
timestamp 1621261055
transform 1 0 3840 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_4
timestamp 1621261055
transform 1 0 1536 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_12
timestamp 1621261055
transform 1 0 2304 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_20
timestamp 1621261055
transform 1 0 3072 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_29
timestamp 1621261055
transform 1 0 3936 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _194_
timestamp 1621261055
transform 1 0 7200 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_22_37
timestamp 1621261055
transform 1 0 4704 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_45
timestamp 1621261055
transform 1 0 5472 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_53
timestamp 1621261055
transform 1 0 6240 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_61
timestamp 1621261055
transform 1 0 7008 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_66
timestamp 1621261055
transform 1 0 7488 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_406
timestamp 1621261055
transform 1 0 9120 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_74
timestamp 1621261055
transform 1 0 8256 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_22_82
timestamp 1621261055
transform 1 0 9024 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_84
timestamp 1621261055
transform 1 0 9216 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_92
timestamp 1621261055
transform 1 0 9984 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_100
timestamp 1621261055
transform 1 0 10752 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_108
timestamp 1621261055
transform 1 0 11520 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_116
timestamp 1621261055
transform 1 0 12288 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_124
timestamp 1621261055
transform 1 0 13056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_132
timestamp 1621261055
transform 1 0 13824 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_407
timestamp 1621261055
transform 1 0 14400 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_136
timestamp 1621261055
transform 1 0 14208 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_139
timestamp 1621261055
transform 1 0 14496 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_147
timestamp 1621261055
transform 1 0 15264 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_155
timestamp 1621261055
transform 1 0 16032 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_163
timestamp 1621261055
transform 1 0 16800 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_408
timestamp 1621261055
transform 1 0 19680 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_171
timestamp 1621261055
transform 1 0 17568 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_179
timestamp 1621261055
transform 1 0 18336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_187
timestamp 1621261055
transform 1 0 19104 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_191
timestamp 1621261055
transform 1 0 19488 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_194
timestamp 1621261055
transform 1 0 19776 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_202
timestamp 1621261055
transform 1 0 20544 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_210
timestamp 1621261055
transform 1 0 21312 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_218
timestamp 1621261055
transform 1 0 22080 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_226
timestamp 1621261055
transform 1 0 22848 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_409
timestamp 1621261055
transform 1 0 24960 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_234
timestamp 1621261055
transform 1 0 23616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_242
timestamp 1621261055
transform 1 0 24384 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_246
timestamp 1621261055
transform 1 0 24768 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_249
timestamp 1621261055
transform 1 0 25056 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_257
timestamp 1621261055
transform 1 0 25824 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_265
timestamp 1621261055
transform 1 0 26592 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_273
timestamp 1621261055
transform 1 0 27360 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_281
timestamp 1621261055
transform 1 0 28128 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_289
timestamp 1621261055
transform 1 0 28896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_297
timestamp 1621261055
transform 1 0 29664 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_410
timestamp 1621261055
transform 1 0 30240 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_301
timestamp 1621261055
transform 1 0 30048 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_304
timestamp 1621261055
transform 1 0 30336 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_312
timestamp 1621261055
transform 1 0 31104 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_320
timestamp 1621261055
transform 1 0 31872 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_328
timestamp 1621261055
transform 1 0 32640 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_411
timestamp 1621261055
transform 1 0 35520 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_336
timestamp 1621261055
transform 1 0 33408 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_344
timestamp 1621261055
transform 1 0 34176 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_352
timestamp 1621261055
transform 1 0 34944 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_356
timestamp 1621261055
transform 1 0 35328 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_359
timestamp 1621261055
transform 1 0 35616 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_367
timestamp 1621261055
transform 1 0 36384 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_375
timestamp 1621261055
transform 1 0 37152 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_383
timestamp 1621261055
transform 1 0 37920 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_391
timestamp 1621261055
transform 1 0 38688 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_412
timestamp 1621261055
transform 1 0 40800 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_399
timestamp 1621261055
transform 1 0 39456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_407
timestamp 1621261055
transform 1 0 40224 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_411
timestamp 1621261055
transform 1 0 40608 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_414
timestamp 1621261055
transform 1 0 40896 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_422
timestamp 1621261055
transform 1 0 41664 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_430
timestamp 1621261055
transform 1 0 42432 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_438
timestamp 1621261055
transform 1 0 43200 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_446
timestamp 1621261055
transform 1 0 43968 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_454
timestamp 1621261055
transform 1 0 44736 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_462
timestamp 1621261055
transform 1 0 45504 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _027_
timestamp 1621261055
transform -1 0 46944 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_413
timestamp 1621261055
transform 1 0 46080 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_14
timestamp 1621261055
transform -1 0 46656 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_466
timestamp 1621261055
transform 1 0 45888 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_469
timestamp 1621261055
transform 1 0 46176 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_22_471
timestamp 1621261055
transform 1 0 46368 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_477
timestamp 1621261055
transform 1 0 46944 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_485
timestamp 1621261055
transform 1 0 47712 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_493
timestamp 1621261055
transform 1 0 48480 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_414
timestamp 1621261055
transform 1 0 51360 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_501
timestamp 1621261055
transform 1 0 49248 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_509
timestamp 1621261055
transform 1 0 50016 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_517
timestamp 1621261055
transform 1 0 50784 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_521
timestamp 1621261055
transform 1 0 51168 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_22_524
timestamp 1621261055
transform 1 0 51456 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_532
timestamp 1621261055
transform 1 0 52224 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_540
timestamp 1621261055
transform 1 0 52992 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_548
timestamp 1621261055
transform 1 0 53760 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_22_556
timestamp 1621261055
transform 1 0 54528 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _068_
timestamp 1621261055
transform 1 0 57120 0 -1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_415
timestamp 1621261055
transform 1 0 56640 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_22_564
timestamp 1621261055
transform 1 0 55296 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_22_572
timestamp 1621261055
transform 1 0 56064 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_576
timestamp 1621261055
transform 1 0 56448 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_22_579
timestamp 1621261055
transform 1 0 56736 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_22_586
timestamp 1621261055
transform 1 0 57408 0 -1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_22_594
timestamp 1621261055
transform 1 0 58176 0 -1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_45
timestamp 1621261055
transform -1 0 58848 0 -1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_22_596
timestamp 1621261055
transform 1 0 58368 0 -1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_4
timestamp 1621261055
transform 1 0 1536 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_4
timestamp 1621261055
transform 1 0 1536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_48
timestamp 1621261055
transform 1 0 1152 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_46
timestamp 1621261055
transform 1 0 1152 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_12
timestamp 1621261055
transform 1 0 2304 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_12
timestamp 1621261055
transform 1 0 2304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_20
timestamp 1621261055
transform 1 0 3072 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_20
timestamp 1621261055
transform 1 0 3072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_29
timestamp 1621261055
transform 1 0 3936 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_28
timestamp 1621261055
transform 1 0 3840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_426
timestamp 1621261055
transform 1 0 3840 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _075_
timestamp 1621261055
transform 1 0 4320 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_36
timestamp 1621261055
transform 1 0 4608 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_36
timestamp 1621261055
transform 1 0 4608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_44
timestamp 1621261055
transform 1 0 5376 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_44
timestamp 1621261055
transform 1 0 5376 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_52
timestamp 1621261055
transform 1 0 6144 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_56
timestamp 1621261055
transform 1 0 6528 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_54
timestamp 1621261055
transform 1 0 6336 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_52
timestamp 1621261055
transform 1 0 6144 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_416
timestamp 1621261055
transform 1 0 6432 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_60
timestamp 1621261055
transform 1 0 6912 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_64
timestamp 1621261055
transform 1 0 7296 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_73
timestamp 1621261055
transform 1 0 7488 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_80
timestamp 1621261055
transform 1 0 8832 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_76
timestamp 1621261055
transform 1 0 8448 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_68
timestamp 1621261055
transform 1 0 7680 0 -1 19314
box -38 -49 806 715
use INVX8  INVX8
timestamp 1623617396
transform 1 0 7680 0 1 17982
box 0 -48 1440 714
use sky130_fd_sc_ls__decap_8  FILLER_24_92
timestamp 1621261055
transform 1 0 9984 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_84
timestamp 1621261055
transform 1 0 9216 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_24_82
timestamp 1621261055
transform 1 0 9024 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_90
timestamp 1621261055
transform 1 0 9792 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_83
timestamp 1621261055
transform 1 0 9120 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_2
timestamp 1621261055
transform -1 0 9504 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_427
timestamp 1621261055
transform 1 0 9120 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _000_
timestamp 1621261055
transform -1 0 9792 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_23_98
timestamp 1621261055
transform 1 0 10560 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_100
timestamp 1621261055
transform 1 0 10752 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_106
timestamp 1621261055
transform 1 0 11328 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_116
timestamp 1621261055
transform 1 0 12288 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_108
timestamp 1621261055
transform 1 0 11520 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_111
timestamp 1621261055
transform 1 0 11808 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_417
timestamp 1621261055
transform 1 0 11712 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_124
timestamp 1621261055
transform 1 0 13056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_119
timestamp 1621261055
transform 1 0 12576 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_132
timestamp 1621261055
transform 1 0 13824 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_127
timestamp 1621261055
transform 1 0 13344 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_139
timestamp 1621261055
transform 1 0 14496 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_136
timestamp 1621261055
transform 1 0 14208 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_135
timestamp 1621261055
transform 1 0 14112 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_428
timestamp 1621261055
transform 1 0 14400 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_146
timestamp 1621261055
transform 1 0 15168 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_143
timestamp 1621261055
transform 1 0 14880 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _084_
timestamp 1621261055
transform 1 0 14880 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_154
timestamp 1621261055
transform 1 0 15936 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_151
timestamp 1621261055
transform 1 0 15648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_162
timestamp 1621261055
transform 1 0 16704 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_163
timestamp 1621261055
transform 1 0 16800 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_159
timestamp 1621261055
transform 1 0 16416 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_418
timestamp 1621261055
transform 1 0 16992 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_170
timestamp 1621261055
transform 1 0 17472 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_166
timestamp 1621261055
transform 1 0 17088 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_178
timestamp 1621261055
transform 1 0 18240 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_182
timestamp 1621261055
transform 1 0 18624 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_174
timestamp 1621261055
transform 1 0 17856 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_190
timestamp 1621261055
transform 1 0 19392 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_186
timestamp 1621261055
transform 1 0 19008 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_190
timestamp 1621261055
transform 1 0 19392 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_194
timestamp 1621261055
transform 1 0 19776 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_24_192
timestamp 1621261055
transform 1 0 19584 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_198
timestamp 1621261055
transform 1 0 20160 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_429
timestamp 1621261055
transform 1 0 19680 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_202
timestamp 1621261055
transform 1 0 20544 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_206
timestamp 1621261055
transform 1 0 20928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_210
timestamp 1621261055
transform 1 0 21312 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_214
timestamp 1621261055
transform 1 0 21696 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_218
timestamp 1621261055
transform 1 0 22080 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_221
timestamp 1621261055
transform 1 0 22368 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_218
timestamp 1621261055
transform 1 0 22080 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_419
timestamp 1621261055
transform 1 0 22272 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_226
timestamp 1621261055
transform 1 0 22848 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_229
timestamp 1621261055
transform 1 0 23136 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_234
timestamp 1621261055
transform 1 0 23616 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_239
timestamp 1621261055
transform 1 0 24096 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_235
timestamp 1621261055
transform 1 0 23712 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_233
timestamp 1621261055
transform 1 0 23520 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _125_
timestamp 1621261055
transform 1 0 23808 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_246
timestamp 1621261055
transform 1 0 24768 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_242
timestamp 1621261055
transform 1 0 24384 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_247
timestamp 1621261055
transform 1 0 24864 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_430
timestamp 1621261055
transform 1 0 24960 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_257
timestamp 1621261055
transform 1 0 25824 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_249
timestamp 1621261055
transform 1 0 25056 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_255
timestamp 1621261055
transform 1 0 25632 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_263
timestamp 1621261055
transform 1 0 26400 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_265
timestamp 1621261055
transform 1 0 26592 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_271
timestamp 1621261055
transform 1 0 27168 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_281
timestamp 1621261055
transform 1 0 28128 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_273
timestamp 1621261055
transform 1 0 27360 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_276
timestamp 1621261055
transform 1 0 27648 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_420
timestamp 1621261055
transform 1 0 27552 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_289
timestamp 1621261055
transform 1 0 28896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_284
timestamp 1621261055
transform 1 0 28416 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_297
timestamp 1621261055
transform 1 0 29664 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_292
timestamp 1621261055
transform 1 0 29184 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_304
timestamp 1621261055
transform 1 0 30336 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_301
timestamp 1621261055
transform 1 0 30048 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_300
timestamp 1621261055
transform 1 0 29952 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_431
timestamp 1621261055
transform 1 0 30240 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_312
timestamp 1621261055
transform 1 0 31104 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_308
timestamp 1621261055
transform 1 0 30720 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_320
timestamp 1621261055
transform 1 0 31872 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_316
timestamp 1621261055
transform 1 0 31488 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_328
timestamp 1621261055
transform 1 0 32640 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_328
timestamp 1621261055
transform 1 0 32640 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_324
timestamp 1621261055
transform 1 0 32256 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_421
timestamp 1621261055
transform 1 0 32832 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_336
timestamp 1621261055
transform 1 0 33408 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_331
timestamp 1621261055
transform 1 0 32928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_344
timestamp 1621261055
transform 1 0 34176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_347
timestamp 1621261055
transform 1 0 34464 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_339
timestamp 1621261055
transform 1 0 33696 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_356
timestamp 1621261055
transform 1 0 35328 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_352
timestamp 1621261055
transform 1 0 34944 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_355
timestamp 1621261055
transform 1 0 35232 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_24_363
timestamp 1621261055
transform 1 0 36000 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_24_359
timestamp 1621261055
transform 1 0 35616 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_363
timestamp 1621261055
transform 1 0 36000 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_432
timestamp 1621261055
transform 1 0 35520 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_369
timestamp 1621261055
transform 1 0 36576 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_371
timestamp 1621261055
transform 1 0 36768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_4
timestamp 1621261055
transform 1 0 36096 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _001_
timestamp 1621261055
transform 1 0 36288 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_377
timestamp 1621261055
transform 1 0 37344 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_379
timestamp 1621261055
transform 1 0 37536 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_385
timestamp 1621261055
transform 1 0 38112 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_386
timestamp 1621261055
transform 1 0 38208 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_383
timestamp 1621261055
transform 1 0 37920 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_422
timestamp 1621261055
transform 1 0 38112 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_393
timestamp 1621261055
transform 1 0 38880 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_394
timestamp 1621261055
transform 1 0 38976 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_24_401
timestamp 1621261055
transform 1 0 39648 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_23_402
timestamp 1621261055
transform 1 0 39744 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _127_
timestamp 1621261055
transform 1 0 39744 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_405
timestamp 1621261055
transform 1 0 40032 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_410
timestamp 1621261055
transform 1 0 40512 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_433
timestamp 1621261055
transform 1 0 40800 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_422
timestamp 1621261055
transform 1 0 41664 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_414
timestamp 1621261055
transform 1 0 40896 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_418
timestamp 1621261055
transform 1 0 41280 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_426
timestamp 1621261055
transform 1 0 42048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_430
timestamp 1621261055
transform 1 0 42432 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_434
timestamp 1621261055
transform 1 0 42816 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_446
timestamp 1621261055
transform 1 0 43968 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_438
timestamp 1621261055
transform 1 0 43200 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_441
timestamp 1621261055
transform 1 0 43488 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_438
timestamp 1621261055
transform 1 0 43200 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_423
timestamp 1621261055
transform 1 0 43392 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _106_
timestamp 1621261055
transform 1 0 43872 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_24_454
timestamp 1621261055
transform 1 0 44736 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_450
timestamp 1621261055
transform 1 0 44352 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_448
timestamp 1621261055
transform 1 0 44160 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_93
timestamp 1621261055
transform -1 0 44640 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _041_
timestamp 1621261055
transform -1 0 44928 0 1 17982
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_24_462
timestamp 1621261055
transform 1 0 45504 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_456
timestamp 1621261055
transform 1 0 44928 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_469
timestamp 1621261055
transform 1 0 46176 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_466
timestamp 1621261055
transform 1 0 45888 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_23_464
timestamp 1621261055
transform 1 0 45696 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_434
timestamp 1621261055
transform 1 0 46080 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_477
timestamp 1621261055
transform 1 0 46944 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_472
timestamp 1621261055
transform 1 0 46464 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_485
timestamp 1621261055
transform 1 0 47712 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_488
timestamp 1621261055
transform 1 0 48000 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_480
timestamp 1621261055
transform 1 0 47232 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_493
timestamp 1621261055
transform 1 0 48480 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_23_494
timestamp 1621261055
transform 1 0 48576 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_492
timestamp 1621261055
transform 1 0 48384 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_424
timestamp 1621261055
transform 1 0 48672 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_501
timestamp 1621261055
transform 1 0 49248 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_496
timestamp 1621261055
transform 1 0 48768 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_509
timestamp 1621261055
transform 1 0 50016 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_512
timestamp 1621261055
transform 1 0 50304 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_504
timestamp 1621261055
transform 1 0 49536 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_521
timestamp 1621261055
transform 1 0 51168 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_517
timestamp 1621261055
transform 1 0 50784 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_520
timestamp 1621261055
transform 1 0 51072 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_524
timestamp 1621261055
transform 1 0 51456 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_528
timestamp 1621261055
transform 1 0 51840 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_435
timestamp 1621261055
transform 1 0 51360 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_532
timestamp 1621261055
transform 1 0 52224 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_536
timestamp 1621261055
transform 1 0 52608 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_540
timestamp 1621261055
transform 1 0 52992 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_23_544
timestamp 1621261055
transform 1 0 53376 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_24_548
timestamp 1621261055
transform 1 0 53760 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_551
timestamp 1621261055
transform 1 0 54048 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_548
timestamp 1621261055
transform 1 0 53760 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_425
timestamp 1621261055
transform 1 0 53952 0 1 17982
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_556
timestamp 1621261055
transform 1 0 54528 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_559
timestamp 1621261055
transform 1 0 54816 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_24_564
timestamp 1621261055
transform 1 0 55296 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_23_567
timestamp 1621261055
transform 1 0 55584 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_576
timestamp 1621261055
transform 1 0 56448 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_24_572
timestamp 1621261055
transform 1 0 56064 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_575
timestamp 1621261055
transform 1 0 56352 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_436
timestamp 1621261055
transform 1 0 56640 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_24_586
timestamp 1621261055
transform 1 0 57408 0 -1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_24_579
timestamp 1621261055
transform 1 0 56736 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_23_583
timestamp 1621261055
transform 1 0 57120 0 1 17982
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _115_
timestamp 1621261055
transform 1 0 57120 0 -1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_24_594
timestamp 1621261055
transform 1 0 58176 0 -1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_23_591
timestamp 1621261055
transform 1 0 57888 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_47
timestamp 1621261055
transform -1 0 58848 0 1 17982
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_49
timestamp 1621261055
transform -1 0 58848 0 -1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_23_595
timestamp 1621261055
transform 1 0 58272 0 1 17982
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_24_596
timestamp 1621261055
transform 1 0 58368 0 -1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_50
timestamp 1621261055
transform 1 0 1152 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_4
timestamp 1621261055
transform 1 0 1536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_12
timestamp 1621261055
transform 1 0 2304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_20
timestamp 1621261055
transform 1 0 3072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_28
timestamp 1621261055
transform 1 0 3840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_437
timestamp 1621261055
transform 1 0 6432 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_78
timestamp 1621261055
transform 1 0 7488 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_36
timestamp 1621261055
transform 1 0 4608 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_44
timestamp 1621261055
transform 1 0 5376 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_52
timestamp 1621261055
transform 1 0 6144 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_25_54
timestamp 1621261055
transform 1 0 6336 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_56
timestamp 1621261055
transform 1 0 6528 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_64
timestamp 1621261055
transform 1 0 7296 0 1 19314
box -38 -49 230 715
use MUX2X1  MUX2X1
timestamp 1623617396
transform 1 0 7680 0 1 19314
box 0 -48 1728 714
use sky130_fd_sc_ls__decap_8  FILLER_25_86
timestamp 1621261055
transform 1 0 9408 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_94
timestamp 1621261055
transform 1 0 10176 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_438
timestamp 1621261055
transform 1 0 11712 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_102
timestamp 1621261055
transform 1 0 10944 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_111
timestamp 1621261055
transform 1 0 11808 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_119
timestamp 1621261055
transform 1 0 12576 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_127
timestamp 1621261055
transform 1 0 13344 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_439
timestamp 1621261055
transform 1 0 16992 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_135
timestamp 1621261055
transform 1 0 14112 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_143
timestamp 1621261055
transform 1 0 14880 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_151
timestamp 1621261055
transform 1 0 15648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_159
timestamp 1621261055
transform 1 0 16416 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_163
timestamp 1621261055
transform 1 0 16800 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_166
timestamp 1621261055
transform 1 0 17088 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_174
timestamp 1621261055
transform 1 0 17856 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_182
timestamp 1621261055
transform 1 0 18624 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_190
timestamp 1621261055
transform 1 0 19392 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_198
timestamp 1621261055
transform 1 0 20160 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_440
timestamp 1621261055
transform 1 0 22272 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_206
timestamp 1621261055
transform 1 0 20928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_214
timestamp 1621261055
transform 1 0 21696 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_218
timestamp 1621261055
transform 1 0 22080 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_221
timestamp 1621261055
transform 1 0 22368 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_229
timestamp 1621261055
transform 1 0 23136 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_237
timestamp 1621261055
transform 1 0 23904 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_245
timestamp 1621261055
transform 1 0 24672 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_253
timestamp 1621261055
transform 1 0 25440 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_261
timestamp 1621261055
transform 1 0 26208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_441
timestamp 1621261055
transform 1 0 27552 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_269
timestamp 1621261055
transform 1 0 26976 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_273
timestamp 1621261055
transform 1 0 27360 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_276
timestamp 1621261055
transform 1 0 27648 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_284
timestamp 1621261055
transform 1 0 28416 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_292
timestamp 1621261055
transform 1 0 29184 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_442
timestamp 1621261055
transform 1 0 32832 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_300
timestamp 1621261055
transform 1 0 29952 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_308
timestamp 1621261055
transform 1 0 30720 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_316
timestamp 1621261055
transform 1 0 31488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_324
timestamp 1621261055
transform 1 0 32256 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_328
timestamp 1621261055
transform 1 0 32640 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_331
timestamp 1621261055
transform 1 0 32928 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_339
timestamp 1621261055
transform 1 0 33696 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_347
timestamp 1621261055
transform 1 0 34464 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_355
timestamp 1621261055
transform 1 0 35232 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_363
timestamp 1621261055
transform 1 0 36000 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_443
timestamp 1621261055
transform 1 0 38112 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_371
timestamp 1621261055
transform 1 0 36768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_379
timestamp 1621261055
transform 1 0 37536 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_383
timestamp 1621261055
transform 1 0 37920 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_386
timestamp 1621261055
transform 1 0 38208 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_394
timestamp 1621261055
transform 1 0 38976 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_402
timestamp 1621261055
transform 1 0 39744 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_410
timestamp 1621261055
transform 1 0 40512 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_418
timestamp 1621261055
transform 1 0 41280 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_426
timestamp 1621261055
transform 1 0 42048 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_444
timestamp 1621261055
transform 1 0 43392 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_25_434
timestamp 1621261055
transform 1 0 42816 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_438
timestamp 1621261055
transform 1 0 43200 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_25_441
timestamp 1621261055
transform 1 0 43488 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_449
timestamp 1621261055
transform 1 0 44256 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_457
timestamp 1621261055
transform 1 0 45024 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_461
timestamp 1621261055
transform 1 0 45408 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _113_
timestamp 1621261055
transform 1 0 45696 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_445
timestamp 1621261055
transform 1 0 48672 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_25_463
timestamp 1621261055
transform 1 0 45600 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_467
timestamp 1621261055
transform 1 0 45984 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_475
timestamp 1621261055
transform 1 0 46752 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_483
timestamp 1621261055
transform 1 0 47520 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_491
timestamp 1621261055
transform 1 0 48288 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_25_496
timestamp 1621261055
transform 1 0 48768 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_504
timestamp 1621261055
transform 1 0 49536 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_512
timestamp 1621261055
transform 1 0 50304 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_520
timestamp 1621261055
transform 1 0 51072 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_528
timestamp 1621261055
transform 1 0 51840 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _128_
timestamp 1621261055
transform 1 0 54528 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _157_
timestamp 1621261055
transform 1 0 52704 0 1 19314
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_446
timestamp 1621261055
transform 1 0 53952 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_25_536
timestamp 1621261055
transform 1 0 52608 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_540
timestamp 1621261055
transform 1 0 52992 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_548
timestamp 1621261055
transform 1 0 53760 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_25_551
timestamp 1621261055
transform 1 0 54048 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_25_555
timestamp 1621261055
transform 1 0 54432 0 1 19314
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_25_559
timestamp 1621261055
transform 1 0 54816 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_567
timestamp 1621261055
transform 1 0 55584 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_575
timestamp 1621261055
transform 1 0 56352 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_25_583
timestamp 1621261055
transform 1 0 57120 0 1 19314
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_25_591
timestamp 1621261055
transform 1 0 57888 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_51
timestamp 1621261055
transform -1 0 58848 0 1 19314
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_25_595
timestamp 1621261055
transform 1 0 58272 0 1 19314
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_52
timestamp 1621261055
transform 1 0 1152 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_447
timestamp 1621261055
transform 1 0 3840 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_4
timestamp 1621261055
transform 1 0 1536 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_12
timestamp 1621261055
transform 1 0 2304 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_20
timestamp 1621261055
transform 1 0 3072 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_29
timestamp 1621261055
transform 1 0 3936 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_37
timestamp 1621261055
transform 1 0 4704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_45
timestamp 1621261055
transform 1 0 5472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_53
timestamp 1621261055
transform 1 0 6240 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_61
timestamp 1621261055
transform 1 0 7008 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_69
timestamp 1621261055
transform 1 0 7776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_81
timestamp 1621261055
transform 1 0 8928 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_26_77
timestamp 1621261055
transform 1 0 8544 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_448
timestamp 1621261055
transform 1 0 9120 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_91
timestamp 1621261055
transform 1 0 9888 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_84
timestamp 1621261055
transform 1 0 9216 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_55
timestamp 1621261055
transform -1 0 9600 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _036_
timestamp 1621261055
transform -1 0 9888 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_99
timestamp 1621261055
transform 1 0 10656 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_26_95
timestamp 1621261055
transform 1 0 10272 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _096_
timestamp 1621261055
transform 1 0 10368 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_26_107
timestamp 1621261055
transform 1 0 11424 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_115
timestamp 1621261055
transform 1 0 12192 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_123
timestamp 1621261055
transform 1 0 12960 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_131
timestamp 1621261055
transform 1 0 13728 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _040_
timestamp 1621261055
transform -1 0 16704 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_449
timestamp 1621261055
transform 1 0 14400 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_91
timestamp 1621261055
transform -1 0 16416 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_135
timestamp 1621261055
transform 1 0 14112 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_137
timestamp 1621261055
transform 1 0 14304 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_139
timestamp 1621261055
transform 1 0 14496 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_147
timestamp 1621261055
transform 1 0 15264 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_155
timestamp 1621261055
transform 1 0 16032 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_162
timestamp 1621261055
transform 1 0 16704 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _213_
timestamp 1621261055
transform 1 0 18624 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_450
timestamp 1621261055
transform 1 0 19680 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_170
timestamp 1621261055
transform 1 0 17472 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_178
timestamp 1621261055
transform 1 0 18240 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_26_185
timestamp 1621261055
transform 1 0 18912 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_194
timestamp 1621261055
transform 1 0 19776 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_202
timestamp 1621261055
transform 1 0 20544 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_210
timestamp 1621261055
transform 1 0 21312 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_218
timestamp 1621261055
transform 1 0 22080 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_226
timestamp 1621261055
transform 1 0 22848 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_451
timestamp 1621261055
transform 1 0 24960 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_234
timestamp 1621261055
transform 1 0 23616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_242
timestamp 1621261055
transform 1 0 24384 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_246
timestamp 1621261055
transform 1 0 24768 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_249
timestamp 1621261055
transform 1 0 25056 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_257
timestamp 1621261055
transform 1 0 25824 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_265
timestamp 1621261055
transform 1 0 26592 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_273
timestamp 1621261055
transform 1 0 27360 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_281
timestamp 1621261055
transform 1 0 28128 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_289
timestamp 1621261055
transform 1 0 28896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_297
timestamp 1621261055
transform 1 0 29664 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_452
timestamp 1621261055
transform 1 0 30240 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_301
timestamp 1621261055
transform 1 0 30048 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_304
timestamp 1621261055
transform 1 0 30336 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_312
timestamp 1621261055
transform 1 0 31104 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_320
timestamp 1621261055
transform 1 0 31872 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_328
timestamp 1621261055
transform 1 0 32640 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_453
timestamp 1621261055
transform 1 0 35520 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_336
timestamp 1621261055
transform 1 0 33408 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_344
timestamp 1621261055
transform 1 0 34176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_352
timestamp 1621261055
transform 1 0 34944 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_356
timestamp 1621261055
transform 1 0 35328 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_359
timestamp 1621261055
transform 1 0 35616 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_367
timestamp 1621261055
transform 1 0 36384 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_375
timestamp 1621261055
transform 1 0 37152 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_383
timestamp 1621261055
transform 1 0 37920 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_391
timestamp 1621261055
transform 1 0 38688 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_454
timestamp 1621261055
transform 1 0 40800 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_399
timestamp 1621261055
transform 1 0 39456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_407
timestamp 1621261055
transform 1 0 40224 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_411
timestamp 1621261055
transform 1 0 40608 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_414
timestamp 1621261055
transform 1 0 40896 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_422
timestamp 1621261055
transform 1 0 41664 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _056_
timestamp 1621261055
transform 1 0 44640 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _185_
timestamp 1621261055
transform 1 0 42528 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_76
timestamp 1621261055
transform 1 0 44448 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_430
timestamp 1621261055
transform 1 0 42432 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_434
timestamp 1621261055
transform 1 0 42816 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_442
timestamp 1621261055
transform 1 0 43584 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_26_450
timestamp 1621261055
transform 1 0 44352 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_456
timestamp 1621261055
transform 1 0 44928 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _134_
timestamp 1621261055
transform 1 0 46944 0 -1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_455
timestamp 1621261055
transform 1 0 46080 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_26_464
timestamp 1621261055
transform 1 0 45696 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_26_469
timestamp 1621261055
transform 1 0 46176 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_480
timestamp 1621261055
transform 1 0 47232 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_488
timestamp 1621261055
transform 1 0 48000 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_456
timestamp 1621261055
transform 1 0 51360 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_496
timestamp 1621261055
transform 1 0 48768 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_504
timestamp 1621261055
transform 1 0 49536 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_512
timestamp 1621261055
transform 1 0 50304 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_520
timestamp 1621261055
transform 1 0 51072 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_26_522
timestamp 1621261055
transform 1 0 51264 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_524
timestamp 1621261055
transform 1 0 51456 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_532
timestamp 1621261055
transform 1 0 52224 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_540
timestamp 1621261055
transform 1 0 52992 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_548
timestamp 1621261055
transform 1 0 53760 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_556
timestamp 1621261055
transform 1 0 54528 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_457
timestamp 1621261055
transform 1 0 56640 0 -1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_26_564
timestamp 1621261055
transform 1 0 55296 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_26_572
timestamp 1621261055
transform 1 0 56064 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_576
timestamp 1621261055
transform 1 0 56448 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_26_579
timestamp 1621261055
transform 1 0 56736 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_26_587
timestamp 1621261055
transform 1 0 57504 0 -1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_53
timestamp 1621261055
transform -1 0 58848 0 -1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_26_595
timestamp 1621261055
transform 1 0 58272 0 -1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_54
timestamp 1621261055
transform 1 0 1152 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_27_4
timestamp 1621261055
transform 1 0 1536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_12
timestamp 1621261055
transform 1 0 2304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_20
timestamp 1621261055
transform 1 0 3072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_28
timestamp 1621261055
transform 1 0 3840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_36
timestamp 1621261055
transform 1 0 4608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_44
timestamp 1621261055
transform 1 0 5376 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_56
timestamp 1621261055
transform 1 0 6528 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_27_54
timestamp 1621261055
transform 1 0 6336 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_52
timestamp 1621261055
transform 1 0 6144 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_458
timestamp 1621261055
transform 1 0 6432 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_27_65
timestamp 1621261055
transform 1 0 7392 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_63
timestamp 1621261055
transform 1 0 7200 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_85
timestamp 1621261055
transform 1 0 7488 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _063_
timestamp 1621261055
transform 1 0 6912 0 1 20646
box -38 -49 326 715
use NAND2X1  NAND2X1
timestamp 1623617396
transform 1 0 7680 0 1 20646
box 0 -48 864 714
use sky130_fd_sc_ls__decap_8  FILLER_27_77
timestamp 1621261055
transform 1 0 8544 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_85
timestamp 1621261055
transform 1 0 9312 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_93
timestamp 1621261055
transform 1 0 10080 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_459
timestamp 1621261055
transform 1 0 11712 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_101
timestamp 1621261055
transform 1 0 10848 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_27_109
timestamp 1621261055
transform 1 0 11616 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_111
timestamp 1621261055
transform 1 0 11808 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_119
timestamp 1621261055
transform 1 0 12576 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_127
timestamp 1621261055
transform 1 0 13344 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_460
timestamp 1621261055
transform 1 0 16992 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_135
timestamp 1621261055
transform 1 0 14112 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_143
timestamp 1621261055
transform 1 0 14880 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_151
timestamp 1621261055
transform 1 0 15648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_159
timestamp 1621261055
transform 1 0 16416 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_163
timestamp 1621261055
transform 1 0 16800 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_166
timestamp 1621261055
transform 1 0 17088 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_174
timestamp 1621261055
transform 1 0 17856 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_182
timestamp 1621261055
transform 1 0 18624 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_190
timestamp 1621261055
transform 1 0 19392 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_198
timestamp 1621261055
transform 1 0 20160 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_461
timestamp 1621261055
transform 1 0 22272 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_206
timestamp 1621261055
transform 1 0 20928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_214
timestamp 1621261055
transform 1 0 21696 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_218
timestamp 1621261055
transform 1 0 22080 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_221
timestamp 1621261055
transform 1 0 22368 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_229
timestamp 1621261055
transform 1 0 23136 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_237
timestamp 1621261055
transform 1 0 23904 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_245
timestamp 1621261055
transform 1 0 24672 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_253
timestamp 1621261055
transform 1 0 25440 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_261
timestamp 1621261055
transform 1 0 26208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_462
timestamp 1621261055
transform 1 0 27552 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_27_269
timestamp 1621261055
transform 1 0 26976 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_273
timestamp 1621261055
transform 1 0 27360 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_276
timestamp 1621261055
transform 1 0 27648 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_284
timestamp 1621261055
transform 1 0 28416 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_292
timestamp 1621261055
transform 1 0 29184 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_463
timestamp 1621261055
transform 1 0 32832 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_300
timestamp 1621261055
transform 1 0 29952 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_308
timestamp 1621261055
transform 1 0 30720 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_316
timestamp 1621261055
transform 1 0 31488 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_324
timestamp 1621261055
transform 1 0 32256 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_328
timestamp 1621261055
transform 1 0 32640 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _092_
timestamp 1621261055
transform 1 0 34176 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_27_331
timestamp 1621261055
transform 1 0 32928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_339
timestamp 1621261055
transform 1 0 33696 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_27_343
timestamp 1621261055
transform 1 0 34080 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_347
timestamp 1621261055
transform 1 0 34464 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_355
timestamp 1621261055
transform 1 0 35232 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_363
timestamp 1621261055
transform 1 0 36000 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_464
timestamp 1621261055
transform 1 0 38112 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_371
timestamp 1621261055
transform 1 0 36768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_379
timestamp 1621261055
transform 1 0 37536 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_383
timestamp 1621261055
transform 1 0 37920 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_386
timestamp 1621261055
transform 1 0 38208 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_394
timestamp 1621261055
transform 1 0 38976 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _026_
timestamp 1621261055
transform 1 0 41184 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_27_402
timestamp 1621261055
transform 1 0 39744 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_410
timestamp 1621261055
transform 1 0 40512 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_414
timestamp 1621261055
transform 1 0 40896 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_416
timestamp 1621261055
transform 1 0 41088 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_420
timestamp 1621261055
transform 1 0 41472 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_428
timestamp 1621261055
transform 1 0 42240 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _025_
timestamp 1621261055
transform -1 0 44160 0 1 20646
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_465
timestamp 1621261055
transform 1 0 43392 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_8
timestamp 1621261055
transform -1 0 43872 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_27_436
timestamp 1621261055
transform 1 0 43008 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_441
timestamp 1621261055
transform 1 0 43488 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_448
timestamp 1621261055
transform 1 0 44160 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_456
timestamp 1621261055
transform 1 0 44928 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_466
timestamp 1621261055
transform 1 0 48672 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_464
timestamp 1621261055
transform 1 0 45696 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_472
timestamp 1621261055
transform 1 0 46464 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_480
timestamp 1621261055
transform 1 0 47232 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_488
timestamp 1621261055
transform 1 0 48000 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_492
timestamp 1621261055
transform 1 0 48384 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_27_494
timestamp 1621261055
transform 1 0 48576 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_496
timestamp 1621261055
transform 1 0 48768 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_504
timestamp 1621261055
transform 1 0 49536 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_512
timestamp 1621261055
transform 1 0 50304 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_520
timestamp 1621261055
transform 1 0 51072 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_528
timestamp 1621261055
transform 1 0 51840 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_467
timestamp 1621261055
transform 1 0 53952 0 1 20646
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_27_536
timestamp 1621261055
transform 1 0 52608 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_544
timestamp 1621261055
transform 1 0 53376 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_548
timestamp 1621261055
transform 1 0 53760 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_27_551
timestamp 1621261055
transform 1 0 54048 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_559
timestamp 1621261055
transform 1 0 54816 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_567
timestamp 1621261055
transform 1 0 55584 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_575
timestamp 1621261055
transform 1 0 56352 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_27_583
timestamp 1621261055
transform 1 0 57120 0 1 20646
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_27_591
timestamp 1621261055
transform 1 0 57888 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_55
timestamp 1621261055
transform -1 0 58848 0 1 20646
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_27_595
timestamp 1621261055
transform 1 0 58272 0 1 20646
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_56
timestamp 1621261055
transform 1 0 1152 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_468
timestamp 1621261055
transform 1 0 3840 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_4
timestamp 1621261055
transform 1 0 1536 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_12
timestamp 1621261055
transform 1 0 2304 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_20
timestamp 1621261055
transform 1 0 3072 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_29
timestamp 1621261055
transform 1 0 3936 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_37
timestamp 1621261055
transform 1 0 4704 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_45
timestamp 1621261055
transform 1 0 5472 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_53
timestamp 1621261055
transform 1 0 6240 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_61
timestamp 1621261055
transform 1 0 7008 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_469
timestamp 1621261055
transform 1 0 9120 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_69
timestamp 1621261055
transform 1 0 7776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_77
timestamp 1621261055
transform 1 0 8544 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_81
timestamp 1621261055
transform 1 0 8928 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_84
timestamp 1621261055
transform 1 0 9216 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_92
timestamp 1621261055
transform 1 0 9984 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_100
timestamp 1621261055
transform 1 0 10752 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_108
timestamp 1621261055
transform 1 0 11520 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_116
timestamp 1621261055
transform 1 0 12288 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_124
timestamp 1621261055
transform 1 0 13056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_132
timestamp 1621261055
transform 1 0 13824 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_470
timestamp 1621261055
transform 1 0 14400 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_136
timestamp 1621261055
transform 1 0 14208 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_139
timestamp 1621261055
transform 1 0 14496 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_147
timestamp 1621261055
transform 1 0 15264 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_155
timestamp 1621261055
transform 1 0 16032 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_163
timestamp 1621261055
transform 1 0 16800 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_471
timestamp 1621261055
transform 1 0 19680 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_171
timestamp 1621261055
transform 1 0 17568 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_179
timestamp 1621261055
transform 1 0 18336 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_187
timestamp 1621261055
transform 1 0 19104 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_191
timestamp 1621261055
transform 1 0 19488 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_194
timestamp 1621261055
transform 1 0 19776 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_202
timestamp 1621261055
transform 1 0 20544 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_210
timestamp 1621261055
transform 1 0 21312 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_218
timestamp 1621261055
transform 1 0 22080 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_226
timestamp 1621261055
transform 1 0 22848 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_472
timestamp 1621261055
transform 1 0 24960 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_234
timestamp 1621261055
transform 1 0 23616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_242
timestamp 1621261055
transform 1 0 24384 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_246
timestamp 1621261055
transform 1 0 24768 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_249
timestamp 1621261055
transform 1 0 25056 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_257
timestamp 1621261055
transform 1 0 25824 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_265
timestamp 1621261055
transform 1 0 26592 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_273
timestamp 1621261055
transform 1 0 27360 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_281
timestamp 1621261055
transform 1 0 28128 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_289
timestamp 1621261055
transform 1 0 28896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_297
timestamp 1621261055
transform 1 0 29664 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_28_304
timestamp 1621261055
transform 1 0 30336 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_301
timestamp 1621261055
transform 1 0 30048 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_473
timestamp 1621261055
transform 1 0 30240 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_28_310
timestamp 1621261055
transform 1 0 30912 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_308
timestamp 1621261055
transform 1 0 30720 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_12
timestamp 1621261055
transform -1 0 31200 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _004_
timestamp 1621261055
transform -1 0 31488 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_320
timestamp 1621261055
transform 1 0 31872 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_28_316
timestamp 1621261055
transform 1 0 31488 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _139_
timestamp 1621261055
transform 1 0 32064 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_28_325
timestamp 1621261055
transform 1 0 32352 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_474
timestamp 1621261055
transform 1 0 35520 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_333
timestamp 1621261055
transform 1 0 33120 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_341
timestamp 1621261055
transform 1 0 33888 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_349
timestamp 1621261055
transform 1 0 34656 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_28_357
timestamp 1621261055
transform 1 0 35424 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_359
timestamp 1621261055
transform 1 0 35616 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_367
timestamp 1621261055
transform 1 0 36384 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_375
timestamp 1621261055
transform 1 0 37152 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_383
timestamp 1621261055
transform 1 0 37920 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_391
timestamp 1621261055
transform 1 0 38688 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_475
timestamp 1621261055
transform 1 0 40800 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_399
timestamp 1621261055
transform 1 0 39456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_407
timestamp 1621261055
transform 1 0 40224 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_411
timestamp 1621261055
transform 1 0 40608 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_414
timestamp 1621261055
transform 1 0 40896 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_422
timestamp 1621261055
transform 1 0 41664 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_430
timestamp 1621261055
transform 1 0 42432 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_438
timestamp 1621261055
transform 1 0 43200 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_446
timestamp 1621261055
transform 1 0 43968 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_454
timestamp 1621261055
transform 1 0 44736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_462
timestamp 1621261055
transform 1 0 45504 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_476
timestamp 1621261055
transform 1 0 46080 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_466
timestamp 1621261055
transform 1 0 45888 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_469
timestamp 1621261055
transform 1 0 46176 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_477
timestamp 1621261055
transform 1 0 46944 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_485
timestamp 1621261055
transform 1 0 47712 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_493
timestamp 1621261055
transform 1 0 48480 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_477
timestamp 1621261055
transform 1 0 51360 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_501
timestamp 1621261055
transform 1 0 49248 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_509
timestamp 1621261055
transform 1 0 50016 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_517
timestamp 1621261055
transform 1 0 50784 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_521
timestamp 1621261055
transform 1 0 51168 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_524
timestamp 1621261055
transform 1 0 51456 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_532
timestamp 1621261055
transform 1 0 52224 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_540
timestamp 1621261055
transform 1 0 52992 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_548
timestamp 1621261055
transform 1 0 53760 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_28_556
timestamp 1621261055
transform 1 0 54528 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _131_
timestamp 1621261055
transform 1 0 57792 0 -1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_478
timestamp 1621261055
transform 1 0 56640 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_28_564
timestamp 1621261055
transform 1 0 55296 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_28_572
timestamp 1621261055
transform 1 0 56064 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_576
timestamp 1621261055
transform 1 0 56448 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_28_579
timestamp 1621261055
transform 1 0 56736 0 -1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_28_587
timestamp 1621261055
transform 1 0 57504 0 -1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_28_589
timestamp 1621261055
transform 1 0 57696 0 -1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_28_593
timestamp 1621261055
transform 1 0 58080 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_57
timestamp 1621261055
transform -1 0 58848 0 -1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _117_
timestamp 1621261055
transform 1 0 2400 0 1 21978
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_58
timestamp 1621261055
transform 1 0 1152 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_29_4
timestamp 1621261055
transform 1 0 1536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_29_12
timestamp 1621261055
transform 1 0 2304 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_16
timestamp 1621261055
transform 1 0 2688 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_24
timestamp 1621261055
transform 1 0 3456 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_32
timestamp 1621261055
transform 1 0 4224 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_479
timestamp 1621261055
transform 1 0 6432 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_40
timestamp 1621261055
transform 1 0 4992 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_48
timestamp 1621261055
transform 1 0 5760 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_52
timestamp 1621261055
transform 1 0 6144 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_29_54
timestamp 1621261055
transform 1 0 6336 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_56
timestamp 1621261055
transform 1 0 6528 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_64
timestamp 1621261055
transform 1 0 7296 0 1 21978
box -38 -49 422 715
use NAND3X1  NAND3X1
timestamp 1623617396
transform 1 0 7680 0 1 21978
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_8  FILLER_29_80
timestamp 1621261055
transform 1 0 8832 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_88
timestamp 1621261055
transform 1 0 9600 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_96
timestamp 1621261055
transform 1 0 10368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_480
timestamp 1621261055
transform 1 0 11712 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_104
timestamp 1621261055
transform 1 0 11136 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_108
timestamp 1621261055
transform 1 0 11520 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_111
timestamp 1621261055
transform 1 0 11808 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_119
timestamp 1621261055
transform 1 0 12576 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_127
timestamp 1621261055
transform 1 0 13344 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_481
timestamp 1621261055
transform 1 0 16992 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_135
timestamp 1621261055
transform 1 0 14112 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_143
timestamp 1621261055
transform 1 0 14880 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_151
timestamp 1621261055
transform 1 0 15648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_159
timestamp 1621261055
transform 1 0 16416 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_163
timestamp 1621261055
transform 1 0 16800 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_166
timestamp 1621261055
transform 1 0 17088 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_174
timestamp 1621261055
transform 1 0 17856 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_182
timestamp 1621261055
transform 1 0 18624 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_190
timestamp 1621261055
transform 1 0 19392 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_198
timestamp 1621261055
transform 1 0 20160 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_482
timestamp 1621261055
transform 1 0 22272 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_206
timestamp 1621261055
transform 1 0 20928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_214
timestamp 1621261055
transform 1 0 21696 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_218
timestamp 1621261055
transform 1 0 22080 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_221
timestamp 1621261055
transform 1 0 22368 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_229
timestamp 1621261055
transform 1 0 23136 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_237
timestamp 1621261055
transform 1 0 23904 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_245
timestamp 1621261055
transform 1 0 24672 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_253
timestamp 1621261055
transform 1 0 25440 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_261
timestamp 1621261055
transform 1 0 26208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_483
timestamp 1621261055
transform 1 0 27552 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_269
timestamp 1621261055
transform 1 0 26976 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_273
timestamp 1621261055
transform 1 0 27360 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_276
timestamp 1621261055
transform 1 0 27648 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_284
timestamp 1621261055
transform 1 0 28416 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_292
timestamp 1621261055
transform 1 0 29184 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_484
timestamp 1621261055
transform 1 0 32832 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_300
timestamp 1621261055
transform 1 0 29952 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_308
timestamp 1621261055
transform 1 0 30720 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_316
timestamp 1621261055
transform 1 0 31488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_324
timestamp 1621261055
transform 1 0 32256 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_328
timestamp 1621261055
transform 1 0 32640 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_331
timestamp 1621261055
transform 1 0 32928 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_339
timestamp 1621261055
transform 1 0 33696 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_347
timestamp 1621261055
transform 1 0 34464 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_355
timestamp 1621261055
transform 1 0 35232 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_363
timestamp 1621261055
transform 1 0 36000 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_485
timestamp 1621261055
transform 1 0 38112 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_371
timestamp 1621261055
transform 1 0 36768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_379
timestamp 1621261055
transform 1 0 37536 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_383
timestamp 1621261055
transform 1 0 37920 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_386
timestamp 1621261055
transform 1 0 38208 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_394
timestamp 1621261055
transform 1 0 38976 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_402
timestamp 1621261055
transform 1 0 39744 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_410
timestamp 1621261055
transform 1 0 40512 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_418
timestamp 1621261055
transform 1 0 41280 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_426
timestamp 1621261055
transform 1 0 42048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_486
timestamp 1621261055
transform 1 0 43392 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_29_434
timestamp 1621261055
transform 1 0 42816 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_438
timestamp 1621261055
transform 1 0 43200 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_441
timestamp 1621261055
transform 1 0 43488 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_449
timestamp 1621261055
transform 1 0 44256 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_457
timestamp 1621261055
transform 1 0 45024 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_487
timestamp 1621261055
transform 1 0 48672 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_465
timestamp 1621261055
transform 1 0 45792 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_473
timestamp 1621261055
transform 1 0 46560 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_481
timestamp 1621261055
transform 1 0 47328 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_489
timestamp 1621261055
transform 1 0 48096 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_493
timestamp 1621261055
transform 1 0 48480 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_496
timestamp 1621261055
transform 1 0 48768 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_504
timestamp 1621261055
transform 1 0 49536 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_512
timestamp 1621261055
transform 1 0 50304 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_520
timestamp 1621261055
transform 1 0 51072 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_528
timestamp 1621261055
transform 1 0 51840 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_488
timestamp 1621261055
transform 1 0 53952 0 1 21978
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_29_536
timestamp 1621261055
transform 1 0 52608 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_544
timestamp 1621261055
transform 1 0 53376 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_548
timestamp 1621261055
transform 1 0 53760 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_29_551
timestamp 1621261055
transform 1 0 54048 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_559
timestamp 1621261055
transform 1 0 54816 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_567
timestamp 1621261055
transform 1 0 55584 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_575
timestamp 1621261055
transform 1 0 56352 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_29_583
timestamp 1621261055
transform 1 0 57120 0 1 21978
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_29_591
timestamp 1621261055
transform 1 0 57888 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_59
timestamp 1621261055
transform -1 0 58848 0 1 21978
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_29_595
timestamp 1621261055
transform 1 0 58272 0 1 21978
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_31_4
timestamp 1621261055
transform 1 0 1536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_4
timestamp 1621261055
transform 1 0 1536 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_62
timestamp 1621261055
transform 1 0 1152 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_60
timestamp 1621261055
transform 1 0 1152 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_12
timestamp 1621261055
transform 1 0 2304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_12
timestamp 1621261055
transform 1 0 2304 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_20
timestamp 1621261055
transform 1 0 3072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_20
timestamp 1621261055
transform 1 0 3072 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_28
timestamp 1621261055
transform 1 0 3840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_29
timestamp 1621261055
transform 1 0 3936 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_489
timestamp 1621261055
transform 1 0 3840 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_36
timestamp 1621261055
transform 1 0 4608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_37
timestamp 1621261055
transform 1 0 4704 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_44
timestamp 1621261055
transform 1 0 5376 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_45
timestamp 1621261055
transform 1 0 5472 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_56
timestamp 1621261055
transform 1 0 6528 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_54
timestamp 1621261055
transform 1 0 6336 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_52
timestamp 1621261055
transform 1 0 6144 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_53
timestamp 1621261055
transform 1 0 6240 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_500
timestamp 1621261055
transform 1 0 6432 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_31_64
timestamp 1621261055
transform 1 0 7296 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_61
timestamp 1621261055
transform 1 0 7008 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_73
timestamp 1621261055
transform 1 0 8160 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_69
timestamp 1621261055
transform 1 0 7776 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _199_
timestamp 1621261055
transform 1 0 7872 0 -1 23310
box -38 -49 326 715
use NOR2X1  NOR2X1
timestamp 1623617396
transform 1 0 7680 0 1 23310
box 0 -48 864 714
use sky130_fd_sc_ls__decap_8  FILLER_31_77
timestamp 1621261055
transform 1 0 8544 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_84
timestamp 1621261055
transform 1 0 9216 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_81
timestamp 1621261055
transform 1 0 8928 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_490
timestamp 1621261055
transform 1 0 9120 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_93
timestamp 1621261055
transform 1 0 10080 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_85
timestamp 1621261055
transform 1 0 9312 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_92
timestamp 1621261055
transform 1 0 9984 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_101
timestamp 1621261055
transform 1 0 10848 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_100
timestamp 1621261055
transform 1 0 10752 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_111
timestamp 1621261055
transform 1 0 11808 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_109
timestamp 1621261055
transform 1 0 11616 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_30_116
timestamp 1621261055
transform 1 0 12288 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_108
timestamp 1621261055
transform 1 0 11520 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_501
timestamp 1621261055
transform 1 0 11712 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_119
timestamp 1621261055
transform 1 0 12576 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_124
timestamp 1621261055
transform 1 0 13056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_127
timestamp 1621261055
transform 1 0 13344 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_132
timestamp 1621261055
transform 1 0 13824 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_135
timestamp 1621261055
transform 1 0 14112 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_139
timestamp 1621261055
transform 1 0 14496 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_136
timestamp 1621261055
transform 1 0 14208 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_491
timestamp 1621261055
transform 1 0 14400 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_143
timestamp 1621261055
transform 1 0 14880 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_147
timestamp 1621261055
transform 1 0 15264 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_151
timestamp 1621261055
transform 1 0 15648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_155
timestamp 1621261055
transform 1 0 16032 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_163
timestamp 1621261055
transform 1 0 16800 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_159
timestamp 1621261055
transform 1 0 16416 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_163
timestamp 1621261055
transform 1 0 16800 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_502
timestamp 1621261055
transform 1 0 16992 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_166
timestamp 1621261055
transform 1 0 17088 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_171
timestamp 1621261055
transform 1 0 17568 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_182
timestamp 1621261055
transform 1 0 18624 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_174
timestamp 1621261055
transform 1 0 17856 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_179
timestamp 1621261055
transform 1 0 18336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_190
timestamp 1621261055
transform 1 0 19392 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_191
timestamp 1621261055
transform 1 0 19488 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_187
timestamp 1621261055
transform 1 0 19104 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_198
timestamp 1621261055
transform 1 0 20160 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_194
timestamp 1621261055
transform 1 0 19776 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_492
timestamp 1621261055
transform 1 0 19680 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_206
timestamp 1621261055
transform 1 0 20928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_202
timestamp 1621261055
transform 1 0 20544 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_214
timestamp 1621261055
transform 1 0 21696 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_210
timestamp 1621261055
transform 1 0 21312 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_221
timestamp 1621261055
transform 1 0 22368 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_218
timestamp 1621261055
transform 1 0 22080 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_218
timestamp 1621261055
transform 1 0 22080 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_503
timestamp 1621261055
transform 1 0 22272 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_229
timestamp 1621261055
transform 1 0 23136 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_226
timestamp 1621261055
transform 1 0 22848 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_237
timestamp 1621261055
transform 1 0 23904 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_234
timestamp 1621261055
transform 1 0 23616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_245
timestamp 1621261055
transform 1 0 24672 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_246
timestamp 1621261055
transform 1 0 24768 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_242
timestamp 1621261055
transform 1 0 24384 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_493
timestamp 1621261055
transform 1 0 24960 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_253
timestamp 1621261055
transform 1 0 25440 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_257
timestamp 1621261055
transform 1 0 25824 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_249
timestamp 1621261055
transform 1 0 25056 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_261
timestamp 1621261055
transform 1 0 26208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_269
timestamp 1621261055
transform 1 0 26976 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_265
timestamp 1621261055
transform 1 0 26592 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_276
timestamp 1621261055
transform 1 0 27648 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_273
timestamp 1621261055
transform 1 0 27360 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_281
timestamp 1621261055
transform 1 0 28128 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_273
timestamp 1621261055
transform 1 0 27360 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_504
timestamp 1621261055
transform 1 0 27552 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_284
timestamp 1621261055
transform 1 0 28416 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_286
timestamp 1621261055
transform 1 0 28608 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _135_
timestamp 1621261055
transform 1 0 28320 0 -1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_292
timestamp 1621261055
transform 1 0 29184 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_294
timestamp 1621261055
transform 1 0 29376 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_300
timestamp 1621261055
transform 1 0 29952 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_304
timestamp 1621261055
transform 1 0 30336 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_30_302
timestamp 1621261055
transform 1 0 30144 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_494
timestamp 1621261055
transform 1 0 30240 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_308
timestamp 1621261055
transform 1 0 30720 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_312
timestamp 1621261055
transform 1 0 31104 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_316
timestamp 1621261055
transform 1 0 31488 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_320
timestamp 1621261055
transform 1 0 31872 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_328
timestamp 1621261055
transform 1 0 32640 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_31_324
timestamp 1621261055
transform 1 0 32256 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_328
timestamp 1621261055
transform 1 0 32640 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_505
timestamp 1621261055
transform 1 0 32832 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_331
timestamp 1621261055
transform 1 0 32928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_336
timestamp 1621261055
transform 1 0 33408 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_347
timestamp 1621261055
transform 1 0 34464 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_339
timestamp 1621261055
transform 1 0 33696 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_344
timestamp 1621261055
transform 1 0 34176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_355
timestamp 1621261055
transform 1 0 35232 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_356
timestamp 1621261055
transform 1 0 35328 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_352
timestamp 1621261055
transform 1 0 34944 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_363
timestamp 1621261055
transform 1 0 36000 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_359
timestamp 1621261055
transform 1 0 35616 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_495
timestamp 1621261055
transform 1 0 35520 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_371
timestamp 1621261055
transform 1 0 36768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_367
timestamp 1621261055
transform 1 0 36384 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_379
timestamp 1621261055
transform 1 0 37536 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_375
timestamp 1621261055
transform 1 0 37152 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_386
timestamp 1621261055
transform 1 0 38208 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_383
timestamp 1621261055
transform 1 0 37920 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_383
timestamp 1621261055
transform 1 0 37920 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_506
timestamp 1621261055
transform 1 0 38112 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_394
timestamp 1621261055
transform 1 0 38976 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_391
timestamp 1621261055
transform 1 0 38688 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_402
timestamp 1621261055
transform 1 0 39744 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_399
timestamp 1621261055
transform 1 0 39456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_410
timestamp 1621261055
transform 1 0 40512 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_411
timestamp 1621261055
transform 1 0 40608 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_407
timestamp 1621261055
transform 1 0 40224 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_496
timestamp 1621261055
transform 1 0 40800 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_418
timestamp 1621261055
transform 1 0 41280 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_422
timestamp 1621261055
transform 1 0 41664 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_414
timestamp 1621261055
transform 1 0 40896 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_426
timestamp 1621261055
transform 1 0 42048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_434
timestamp 1621261055
transform 1 0 42816 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_430
timestamp 1621261055
transform 1 0 42432 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_441
timestamp 1621261055
transform 1 0 43488 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_438
timestamp 1621261055
transform 1 0 43200 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_446
timestamp 1621261055
transform 1 0 43968 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_438
timestamp 1621261055
transform 1 0 43200 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_507
timestamp 1621261055
transform 1 0 43392 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _173_
timestamp 1621261055
transform 1 0 43872 0 1 23310
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_31_448
timestamp 1621261055
transform 1 0 44160 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_454
timestamp 1621261055
transform 1 0 44736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_456
timestamp 1621261055
transform 1 0 44928 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_30_462
timestamp 1621261055
transform 1 0 45504 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_464
timestamp 1621261055
transform 1 0 45696 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_469
timestamp 1621261055
transform 1 0 46176 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_466
timestamp 1621261055
transform 1 0 45888 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_497
timestamp 1621261055
transform 1 0 46080 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_472
timestamp 1621261055
transform 1 0 46464 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_477
timestamp 1621261055
transform 1 0 46944 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_488
timestamp 1621261055
transform 1 0 48000 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_480
timestamp 1621261055
transform 1 0 47232 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_485
timestamp 1621261055
transform 1 0 47712 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_31_494
timestamp 1621261055
transform 1 0 48576 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_492
timestamp 1621261055
transform 1 0 48384 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_493
timestamp 1621261055
transform 1 0 48480 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_508
timestamp 1621261055
transform 1 0 48672 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_496
timestamp 1621261055
transform 1 0 48768 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_501
timestamp 1621261055
transform 1 0 49248 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_512
timestamp 1621261055
transform 1 0 50304 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_504
timestamp 1621261055
transform 1 0 49536 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_509
timestamp 1621261055
transform 1 0 50016 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_520
timestamp 1621261055
transform 1 0 51072 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_521
timestamp 1621261055
transform 1 0 51168 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_517
timestamp 1621261055
transform 1 0 50784 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_31_528
timestamp 1621261055
transform 1 0 51840 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_524
timestamp 1621261055
transform 1 0 51456 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_498
timestamp 1621261055
transform 1 0 51360 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_536
timestamp 1621261055
transform 1 0 52608 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_532
timestamp 1621261055
transform 1 0 52224 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_544
timestamp 1621261055
transform 1 0 53376 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_30_540
timestamp 1621261055
transform 1 0 52992 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_551
timestamp 1621261055
transform 1 0 54048 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_548
timestamp 1621261055
transform 1 0 53760 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_30_548
timestamp 1621261055
transform 1 0 53760 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_509
timestamp 1621261055
transform 1 0 53952 0 1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_559
timestamp 1621261055
transform 1 0 54816 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_556
timestamp 1621261055
transform 1 0 54528 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_567
timestamp 1621261055
transform 1 0 55584 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_564
timestamp 1621261055
transform 1 0 55296 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_31_575
timestamp 1621261055
transform 1 0 56352 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_576
timestamp 1621261055
transform 1 0 56448 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_30_572
timestamp 1621261055
transform 1 0 56064 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_499
timestamp 1621261055
transform 1 0 56640 0 -1 23310
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_31_583
timestamp 1621261055
transform 1 0 57120 0 1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_587
timestamp 1621261055
transform 1 0 57504 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_30_579
timestamp 1621261055
transform 1 0 56736 0 -1 23310
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_31_591
timestamp 1621261055
transform 1 0 57888 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_61
timestamp 1621261055
transform -1 0 58848 0 -1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_63
timestamp 1621261055
transform -1 0 58848 0 1 23310
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_30_595
timestamp 1621261055
transform 1 0 58272 0 -1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_31_595
timestamp 1621261055
transform 1 0 58272 0 1 23310
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_8
timestamp 1621261055
transform 1 0 1920 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_32_4
timestamp 1621261055
transform 1 0 1536 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_64
timestamp 1621261055
transform 1 0 1152 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_15
timestamp 1621261055
transform 1 0 2592 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_39
timestamp 1621261055
transform 1 0 2112 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _043_
timestamp 1621261055
transform 1 0 2304 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_32_23
timestamp 1621261055
transform 1 0 3360 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_32_29
timestamp 1621261055
transform 1 0 3936 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_32_27
timestamp 1621261055
transform 1 0 3744 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_510
timestamp 1621261055
transform 1 0 3840 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_37
timestamp 1621261055
transform 1 0 4704 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_45
timestamp 1621261055
transform 1 0 5472 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_53
timestamp 1621261055
transform 1 0 6240 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_61
timestamp 1621261055
transform 1 0 7008 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_511
timestamp 1621261055
transform 1 0 9120 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_69
timestamp 1621261055
transform 1 0 7776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_77
timestamp 1621261055
transform 1 0 8544 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_81
timestamp 1621261055
transform 1 0 8928 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_84
timestamp 1621261055
transform 1 0 9216 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_92
timestamp 1621261055
transform 1 0 9984 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _077_
timestamp 1621261055
transform 1 0 13152 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_32_100
timestamp 1621261055
transform 1 0 10752 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_108
timestamp 1621261055
transform 1 0 11520 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_116
timestamp 1621261055
transform 1 0 12288 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_32_124
timestamp 1621261055
transform 1 0 13056 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_128
timestamp 1621261055
transform 1 0 13440 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_512
timestamp 1621261055
transform 1 0 14400 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_136
timestamp 1621261055
transform 1 0 14208 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_139
timestamp 1621261055
transform 1 0 14496 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_147
timestamp 1621261055
transform 1 0 15264 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_155
timestamp 1621261055
transform 1 0 16032 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_163
timestamp 1621261055
transform 1 0 16800 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_513
timestamp 1621261055
transform 1 0 19680 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_171
timestamp 1621261055
transform 1 0 17568 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_179
timestamp 1621261055
transform 1 0 18336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_187
timestamp 1621261055
transform 1 0 19104 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_191
timestamp 1621261055
transform 1 0 19488 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_194
timestamp 1621261055
transform 1 0 19776 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_202
timestamp 1621261055
transform 1 0 20544 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_210
timestamp 1621261055
transform 1 0 21312 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_218
timestamp 1621261055
transform 1 0 22080 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_226
timestamp 1621261055
transform 1 0 22848 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_514
timestamp 1621261055
transform 1 0 24960 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_234
timestamp 1621261055
transform 1 0 23616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_242
timestamp 1621261055
transform 1 0 24384 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_246
timestamp 1621261055
transform 1 0 24768 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_249
timestamp 1621261055
transform 1 0 25056 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_257
timestamp 1621261055
transform 1 0 25824 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_265
timestamp 1621261055
transform 1 0 26592 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_273
timestamp 1621261055
transform 1 0 27360 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_281
timestamp 1621261055
transform 1 0 28128 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_289
timestamp 1621261055
transform 1 0 28896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_297
timestamp 1621261055
transform 1 0 29664 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_515
timestamp 1621261055
transform 1 0 30240 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_301
timestamp 1621261055
transform 1 0 30048 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_304
timestamp 1621261055
transform 1 0 30336 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_312
timestamp 1621261055
transform 1 0 31104 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_320
timestamp 1621261055
transform 1 0 31872 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_328
timestamp 1621261055
transform 1 0 32640 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_516
timestamp 1621261055
transform 1 0 35520 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_336
timestamp 1621261055
transform 1 0 33408 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_344
timestamp 1621261055
transform 1 0 34176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_352
timestamp 1621261055
transform 1 0 34944 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_356
timestamp 1621261055
transform 1 0 35328 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_359
timestamp 1621261055
transform 1 0 35616 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _039_
timestamp 1621261055
transform -1 0 37152 0 -1 24642
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_89
timestamp 1621261055
transform -1 0 36864 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_367
timestamp 1621261055
transform 1 0 36384 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_32_369
timestamp 1621261055
transform 1 0 36576 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_375
timestamp 1621261055
transform 1 0 37152 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_383
timestamp 1621261055
transform 1 0 37920 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_391
timestamp 1621261055
transform 1 0 38688 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_517
timestamp 1621261055
transform 1 0 40800 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_399
timestamp 1621261055
transform 1 0 39456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_407
timestamp 1621261055
transform 1 0 40224 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_411
timestamp 1621261055
transform 1 0 40608 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_414
timestamp 1621261055
transform 1 0 40896 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_422
timestamp 1621261055
transform 1 0 41664 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_430
timestamp 1621261055
transform 1 0 42432 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_438
timestamp 1621261055
transform 1 0 43200 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_446
timestamp 1621261055
transform 1 0 43968 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_454
timestamp 1621261055
transform 1 0 44736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_462
timestamp 1621261055
transform 1 0 45504 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_518
timestamp 1621261055
transform 1 0 46080 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_466
timestamp 1621261055
transform 1 0 45888 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_469
timestamp 1621261055
transform 1 0 46176 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_477
timestamp 1621261055
transform 1 0 46944 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_485
timestamp 1621261055
transform 1 0 47712 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_493
timestamp 1621261055
transform 1 0 48480 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_519
timestamp 1621261055
transform 1 0 51360 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_501
timestamp 1621261055
transform 1 0 49248 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_509
timestamp 1621261055
transform 1 0 50016 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_517
timestamp 1621261055
transform 1 0 50784 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_521
timestamp 1621261055
transform 1 0 51168 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_524
timestamp 1621261055
transform 1 0 51456 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_532
timestamp 1621261055
transform 1 0 52224 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_540
timestamp 1621261055
transform 1 0 52992 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_548
timestamp 1621261055
transform 1 0 53760 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_556
timestamp 1621261055
transform 1 0 54528 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_520
timestamp 1621261055
transform 1 0 56640 0 -1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_32_564
timestamp 1621261055
transform 1 0 55296 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_32_572
timestamp 1621261055
transform 1 0 56064 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_576
timestamp 1621261055
transform 1 0 56448 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_32_579
timestamp 1621261055
transform 1 0 56736 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_32_587
timestamp 1621261055
transform 1 0 57504 0 -1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_65
timestamp 1621261055
transform -1 0 58848 0 -1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_32_595
timestamp 1621261055
transform 1 0 58272 0 -1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_66
timestamp 1621261055
transform 1 0 1152 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_33_4
timestamp 1621261055
transform 1 0 1536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_12
timestamp 1621261055
transform 1 0 2304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_20
timestamp 1621261055
transform 1 0 3072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_28
timestamp 1621261055
transform 1 0 3840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_521
timestamp 1621261055
transform 1 0 6432 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_36
timestamp 1621261055
transform 1 0 4608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_44
timestamp 1621261055
transform 1 0 5376 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_52
timestamp 1621261055
transform 1 0 6144 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_33_54
timestamp 1621261055
transform 1 0 6336 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_56
timestamp 1621261055
transform 1 0 6528 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_64
timestamp 1621261055
transform 1 0 7296 0 1 24642
box -38 -49 422 715
use OAI21X1  OAI21X1
timestamp 1623617396
transform 1 0 7680 0 1 24642
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_8  FILLER_33_80
timestamp 1621261055
transform 1 0 8832 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_88
timestamp 1621261055
transform 1 0 9600 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_96
timestamp 1621261055
transform 1 0 10368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_522
timestamp 1621261055
transform 1 0 11712 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_104
timestamp 1621261055
transform 1 0 11136 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_108
timestamp 1621261055
transform 1 0 11520 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_111
timestamp 1621261055
transform 1 0 11808 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_119
timestamp 1621261055
transform 1 0 12576 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_127
timestamp 1621261055
transform 1 0 13344 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_523
timestamp 1621261055
transform 1 0 16992 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_135
timestamp 1621261055
transform 1 0 14112 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_143
timestamp 1621261055
transform 1 0 14880 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_151
timestamp 1621261055
transform 1 0 15648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_159
timestamp 1621261055
transform 1 0 16416 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_163
timestamp 1621261055
transform 1 0 16800 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_166
timestamp 1621261055
transform 1 0 17088 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_174
timestamp 1621261055
transform 1 0 17856 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_182
timestamp 1621261055
transform 1 0 18624 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_190
timestamp 1621261055
transform 1 0 19392 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_198
timestamp 1621261055
transform 1 0 20160 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_524
timestamp 1621261055
transform 1 0 22272 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_206
timestamp 1621261055
transform 1 0 20928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_214
timestamp 1621261055
transform 1 0 21696 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_218
timestamp 1621261055
transform 1 0 22080 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_221
timestamp 1621261055
transform 1 0 22368 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_229
timestamp 1621261055
transform 1 0 23136 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_237
timestamp 1621261055
transform 1 0 23904 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_245
timestamp 1621261055
transform 1 0 24672 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_253
timestamp 1621261055
transform 1 0 25440 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_261
timestamp 1621261055
transform 1 0 26208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_525
timestamp 1621261055
transform 1 0 27552 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_269
timestamp 1621261055
transform 1 0 26976 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_273
timestamp 1621261055
transform 1 0 27360 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_276
timestamp 1621261055
transform 1 0 27648 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_284
timestamp 1621261055
transform 1 0 28416 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_292
timestamp 1621261055
transform 1 0 29184 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_526
timestamp 1621261055
transform 1 0 32832 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_300
timestamp 1621261055
transform 1 0 29952 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_308
timestamp 1621261055
transform 1 0 30720 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_316
timestamp 1621261055
transform 1 0 31488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_324
timestamp 1621261055
transform 1 0 32256 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_328
timestamp 1621261055
transform 1 0 32640 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_331
timestamp 1621261055
transform 1 0 32928 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_339
timestamp 1621261055
transform 1 0 33696 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_347
timestamp 1621261055
transform 1 0 34464 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_355
timestamp 1621261055
transform 1 0 35232 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_363
timestamp 1621261055
transform 1 0 36000 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_527
timestamp 1621261055
transform 1 0 38112 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_371
timestamp 1621261055
transform 1 0 36768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_379
timestamp 1621261055
transform 1 0 37536 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_383
timestamp 1621261055
transform 1 0 37920 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_386
timestamp 1621261055
transform 1 0 38208 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_394
timestamp 1621261055
transform 1 0 38976 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_402
timestamp 1621261055
transform 1 0 39744 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_410
timestamp 1621261055
transform 1 0 40512 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_418
timestamp 1621261055
transform 1 0 41280 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_426
timestamp 1621261055
transform 1 0 42048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_528
timestamp 1621261055
transform 1 0 43392 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_33_434
timestamp 1621261055
transform 1 0 42816 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_438
timestamp 1621261055
transform 1 0 43200 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_441
timestamp 1621261055
transform 1 0 43488 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_449
timestamp 1621261055
transform 1 0 44256 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_457
timestamp 1621261055
transform 1 0 45024 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_529
timestamp 1621261055
transform 1 0 48672 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_465
timestamp 1621261055
transform 1 0 45792 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_473
timestamp 1621261055
transform 1 0 46560 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_481
timestamp 1621261055
transform 1 0 47328 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_489
timestamp 1621261055
transform 1 0 48096 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_493
timestamp 1621261055
transform 1 0 48480 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_496
timestamp 1621261055
transform 1 0 48768 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_504
timestamp 1621261055
transform 1 0 49536 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_512
timestamp 1621261055
transform 1 0 50304 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_520
timestamp 1621261055
transform 1 0 51072 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_528
timestamp 1621261055
transform 1 0 51840 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_530
timestamp 1621261055
transform 1 0 53952 0 1 24642
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_33_536
timestamp 1621261055
transform 1 0 52608 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_544
timestamp 1621261055
transform 1 0 53376 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_548
timestamp 1621261055
transform 1 0 53760 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_33_551
timestamp 1621261055
transform 1 0 54048 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_559
timestamp 1621261055
transform 1 0 54816 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_567
timestamp 1621261055
transform 1 0 55584 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_575
timestamp 1621261055
transform 1 0 56352 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_33_583
timestamp 1621261055
transform 1 0 57120 0 1 24642
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_33_591
timestamp 1621261055
transform 1 0 57888 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_67
timestamp 1621261055
transform -1 0 58848 0 1 24642
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_33_595
timestamp 1621261055
transform 1 0 58272 0 1 24642
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_68
timestamp 1621261055
transform 1 0 1152 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_531
timestamp 1621261055
transform 1 0 3840 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_4
timestamp 1621261055
transform 1 0 1536 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_12
timestamp 1621261055
transform 1 0 2304 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_20
timestamp 1621261055
transform 1 0 3072 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_29
timestamp 1621261055
transform 1 0 3936 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_37
timestamp 1621261055
transform 1 0 4704 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_45
timestamp 1621261055
transform 1 0 5472 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_53
timestamp 1621261055
transform 1 0 6240 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_61
timestamp 1621261055
transform 1 0 7008 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_532
timestamp 1621261055
transform 1 0 9120 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_69
timestamp 1621261055
transform 1 0 7776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_77
timestamp 1621261055
transform 1 0 8544 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_81
timestamp 1621261055
transform 1 0 8928 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_84
timestamp 1621261055
transform 1 0 9216 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_92
timestamp 1621261055
transform 1 0 9984 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_100
timestamp 1621261055
transform 1 0 10752 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_108
timestamp 1621261055
transform 1 0 11520 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_116
timestamp 1621261055
transform 1 0 12288 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_124
timestamp 1621261055
transform 1 0 13056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_132
timestamp 1621261055
transform 1 0 13824 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_533
timestamp 1621261055
transform 1 0 14400 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_136
timestamp 1621261055
transform 1 0 14208 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_139
timestamp 1621261055
transform 1 0 14496 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_147
timestamp 1621261055
transform 1 0 15264 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_155
timestamp 1621261055
transform 1 0 16032 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_163
timestamp 1621261055
transform 1 0 16800 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_534
timestamp 1621261055
transform 1 0 19680 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_171
timestamp 1621261055
transform 1 0 17568 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_179
timestamp 1621261055
transform 1 0 18336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_187
timestamp 1621261055
transform 1 0 19104 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_191
timestamp 1621261055
transform 1 0 19488 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_194
timestamp 1621261055
transform 1 0 19776 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_202
timestamp 1621261055
transform 1 0 20544 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_210
timestamp 1621261055
transform 1 0 21312 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_218
timestamp 1621261055
transform 1 0 22080 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_226
timestamp 1621261055
transform 1 0 22848 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_535
timestamp 1621261055
transform 1 0 24960 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_234
timestamp 1621261055
transform 1 0 23616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_242
timestamp 1621261055
transform 1 0 24384 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_246
timestamp 1621261055
transform 1 0 24768 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_249
timestamp 1621261055
transform 1 0 25056 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_257
timestamp 1621261055
transform 1 0 25824 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_265
timestamp 1621261055
transform 1 0 26592 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_273
timestamp 1621261055
transform 1 0 27360 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_281
timestamp 1621261055
transform 1 0 28128 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_289
timestamp 1621261055
transform 1 0 28896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_297
timestamp 1621261055
transform 1 0 29664 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_536
timestamp 1621261055
transform 1 0 30240 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_301
timestamp 1621261055
transform 1 0 30048 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_304
timestamp 1621261055
transform 1 0 30336 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_312
timestamp 1621261055
transform 1 0 31104 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_320
timestamp 1621261055
transform 1 0 31872 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_328
timestamp 1621261055
transform 1 0 32640 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_537
timestamp 1621261055
transform 1 0 35520 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_336
timestamp 1621261055
transform 1 0 33408 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_344
timestamp 1621261055
transform 1 0 34176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_352
timestamp 1621261055
transform 1 0 34944 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_356
timestamp 1621261055
transform 1 0 35328 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_359
timestamp 1621261055
transform 1 0 35616 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_367
timestamp 1621261055
transform 1 0 36384 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_375
timestamp 1621261055
transform 1 0 37152 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_383
timestamp 1621261055
transform 1 0 37920 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_391
timestamp 1621261055
transform 1 0 38688 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_538
timestamp 1621261055
transform 1 0 40800 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_399
timestamp 1621261055
transform 1 0 39456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_407
timestamp 1621261055
transform 1 0 40224 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_411
timestamp 1621261055
transform 1 0 40608 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_414
timestamp 1621261055
transform 1 0 40896 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_422
timestamp 1621261055
transform 1 0 41664 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_430
timestamp 1621261055
transform 1 0 42432 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_438
timestamp 1621261055
transform 1 0 43200 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_446
timestamp 1621261055
transform 1 0 43968 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_454
timestamp 1621261055
transform 1 0 44736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_462
timestamp 1621261055
transform 1 0 45504 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_539
timestamp 1621261055
transform 1 0 46080 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_466
timestamp 1621261055
transform 1 0 45888 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_469
timestamp 1621261055
transform 1 0 46176 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_477
timestamp 1621261055
transform 1 0 46944 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_485
timestamp 1621261055
transform 1 0 47712 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_493
timestamp 1621261055
transform 1 0 48480 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_540
timestamp 1621261055
transform 1 0 51360 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_501
timestamp 1621261055
transform 1 0 49248 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_509
timestamp 1621261055
transform 1 0 50016 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_517
timestamp 1621261055
transform 1 0 50784 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_521
timestamp 1621261055
transform 1 0 51168 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_524
timestamp 1621261055
transform 1 0 51456 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_532
timestamp 1621261055
transform 1 0 52224 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_540
timestamp 1621261055
transform 1 0 52992 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_548
timestamp 1621261055
transform 1 0 53760 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_556
timestamp 1621261055
transform 1 0 54528 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_541
timestamp 1621261055
transform 1 0 56640 0 -1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_34_564
timestamp 1621261055
transform 1 0 55296 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_34_572
timestamp 1621261055
transform 1 0 56064 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_576
timestamp 1621261055
transform 1 0 56448 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_34_579
timestamp 1621261055
transform 1 0 56736 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_34_587
timestamp 1621261055
transform 1 0 57504 0 -1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_69
timestamp 1621261055
transform -1 0 58848 0 -1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_34_595
timestamp 1621261055
transform 1 0 58272 0 -1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_70
timestamp 1621261055
transform 1 0 1152 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_4
timestamp 1621261055
transform 1 0 1536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_12
timestamp 1621261055
transform 1 0 2304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_20
timestamp 1621261055
transform 1 0 3072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_28
timestamp 1621261055
transform 1 0 3840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_542
timestamp 1621261055
transform 1 0 6432 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_36
timestamp 1621261055
transform 1 0 4608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_44
timestamp 1621261055
transform 1 0 5376 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_52
timestamp 1621261055
transform 1 0 6144 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_54
timestamp 1621261055
transform 1 0 6336 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_56
timestamp 1621261055
transform 1 0 6528 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_64
timestamp 1621261055
transform 1 0 7296 0 1 25974
box -38 -49 422 715
use OAI22X1  OAI22X1
timestamp 1623617396
transform 1 0 7680 0 1 25974
box 0 -48 1440 714
use sky130_fd_sc_ls__decap_8  FILLER_35_83
timestamp 1621261055
transform 1 0 9120 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_91
timestamp 1621261055
transform 1 0 9888 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_99
timestamp 1621261055
transform 1 0 10656 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_543
timestamp 1621261055
transform 1 0 11712 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_107
timestamp 1621261055
transform 1 0 11424 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_109
timestamp 1621261055
transform 1 0 11616 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_111
timestamp 1621261055
transform 1 0 11808 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_119
timestamp 1621261055
transform 1 0 12576 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_127
timestamp 1621261055
transform 1 0 13344 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_544
timestamp 1621261055
transform 1 0 16992 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_135
timestamp 1621261055
transform 1 0 14112 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_143
timestamp 1621261055
transform 1 0 14880 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_151
timestamp 1621261055
transform 1 0 15648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_159
timestamp 1621261055
transform 1 0 16416 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_163
timestamp 1621261055
transform 1 0 16800 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_166
timestamp 1621261055
transform 1 0 17088 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_174
timestamp 1621261055
transform 1 0 17856 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_182
timestamp 1621261055
transform 1 0 18624 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_190
timestamp 1621261055
transform 1 0 19392 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_198
timestamp 1621261055
transform 1 0 20160 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_545
timestamp 1621261055
transform 1 0 22272 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_206
timestamp 1621261055
transform 1 0 20928 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_214
timestamp 1621261055
transform 1 0 21696 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_218
timestamp 1621261055
transform 1 0 22080 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_221
timestamp 1621261055
transform 1 0 22368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_229
timestamp 1621261055
transform 1 0 23136 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_237
timestamp 1621261055
transform 1 0 23904 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_245
timestamp 1621261055
transform 1 0 24672 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_253
timestamp 1621261055
transform 1 0 25440 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_261
timestamp 1621261055
transform 1 0 26208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_546
timestamp 1621261055
transform 1 0 27552 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_269
timestamp 1621261055
transform 1 0 26976 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_273
timestamp 1621261055
transform 1 0 27360 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_276
timestamp 1621261055
transform 1 0 27648 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_284
timestamp 1621261055
transform 1 0 28416 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_292
timestamp 1621261055
transform 1 0 29184 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_547
timestamp 1621261055
transform 1 0 32832 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_300
timestamp 1621261055
transform 1 0 29952 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_308
timestamp 1621261055
transform 1 0 30720 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_316
timestamp 1621261055
transform 1 0 31488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_324
timestamp 1621261055
transform 1 0 32256 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_328
timestamp 1621261055
transform 1 0 32640 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _184_
timestamp 1621261055
transform 1 0 33312 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_35_331
timestamp 1621261055
transform 1 0 32928 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_35_338
timestamp 1621261055
transform 1 0 33600 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_346
timestamp 1621261055
transform 1 0 34368 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_354
timestamp 1621261055
transform 1 0 35136 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_362
timestamp 1621261055
transform 1 0 35904 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _006_
timestamp 1621261055
transform -1 0 36864 0 1 25974
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_548
timestamp 1621261055
transform 1 0 38112 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_18
timestamp 1621261055
transform -1 0 36576 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_35_366
timestamp 1621261055
transform 1 0 36288 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_372
timestamp 1621261055
transform 1 0 36864 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_380
timestamp 1621261055
transform 1 0 37632 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_35_384
timestamp 1621261055
transform 1 0 38016 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_386
timestamp 1621261055
transform 1 0 38208 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_394
timestamp 1621261055
transform 1 0 38976 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_402
timestamp 1621261055
transform 1 0 39744 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_410
timestamp 1621261055
transform 1 0 40512 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_418
timestamp 1621261055
transform 1 0 41280 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_426
timestamp 1621261055
transform 1 0 42048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_549
timestamp 1621261055
transform 1 0 43392 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_35_434
timestamp 1621261055
transform 1 0 42816 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_438
timestamp 1621261055
transform 1 0 43200 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_441
timestamp 1621261055
transform 1 0 43488 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_449
timestamp 1621261055
transform 1 0 44256 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_457
timestamp 1621261055
transform 1 0 45024 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_550
timestamp 1621261055
transform 1 0 48672 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_465
timestamp 1621261055
transform 1 0 45792 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_473
timestamp 1621261055
transform 1 0 46560 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_481
timestamp 1621261055
transform 1 0 47328 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_489
timestamp 1621261055
transform 1 0 48096 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_493
timestamp 1621261055
transform 1 0 48480 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_496
timestamp 1621261055
transform 1 0 48768 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_504
timestamp 1621261055
transform 1 0 49536 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_512
timestamp 1621261055
transform 1 0 50304 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_520
timestamp 1621261055
transform 1 0 51072 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_528
timestamp 1621261055
transform 1 0 51840 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_551
timestamp 1621261055
transform 1 0 53952 0 1 25974
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_35_536
timestamp 1621261055
transform 1 0 52608 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_544
timestamp 1621261055
transform 1 0 53376 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_548
timestamp 1621261055
transform 1 0 53760 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_35_551
timestamp 1621261055
transform 1 0 54048 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_559
timestamp 1621261055
transform 1 0 54816 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_567
timestamp 1621261055
transform 1 0 55584 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_575
timestamp 1621261055
transform 1 0 56352 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_35_583
timestamp 1621261055
transform 1 0 57120 0 1 25974
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_35_591
timestamp 1621261055
transform 1 0 57888 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_71
timestamp 1621261055
transform -1 0 58848 0 1 25974
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_35_595
timestamp 1621261055
transform 1 0 58272 0 1 25974
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_72
timestamp 1621261055
transform 1 0 1152 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_552
timestamp 1621261055
transform 1 0 3840 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_4
timestamp 1621261055
transform 1 0 1536 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_12
timestamp 1621261055
transform 1 0 2304 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_20
timestamp 1621261055
transform 1 0 3072 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_29
timestamp 1621261055
transform 1 0 3936 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_37
timestamp 1621261055
transform 1 0 4704 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_45
timestamp 1621261055
transform 1 0 5472 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_53
timestamp 1621261055
transform 1 0 6240 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_61
timestamp 1621261055
transform 1 0 7008 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_553
timestamp 1621261055
transform 1 0 9120 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_69
timestamp 1621261055
transform 1 0 7776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_77
timestamp 1621261055
transform 1 0 8544 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_81
timestamp 1621261055
transform 1 0 8928 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_84
timestamp 1621261055
transform 1 0 9216 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_92
timestamp 1621261055
transform 1 0 9984 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_100
timestamp 1621261055
transform 1 0 10752 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_108
timestamp 1621261055
transform 1 0 11520 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_116
timestamp 1621261055
transform 1 0 12288 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_124
timestamp 1621261055
transform 1 0 13056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_132
timestamp 1621261055
transform 1 0 13824 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_554
timestamp 1621261055
transform 1 0 14400 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_136
timestamp 1621261055
transform 1 0 14208 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_139
timestamp 1621261055
transform 1 0 14496 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_147
timestamp 1621261055
transform 1 0 15264 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_155
timestamp 1621261055
transform 1 0 16032 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_163
timestamp 1621261055
transform 1 0 16800 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_555
timestamp 1621261055
transform 1 0 19680 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_171
timestamp 1621261055
transform 1 0 17568 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_179
timestamp 1621261055
transform 1 0 18336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_187
timestamp 1621261055
transform 1 0 19104 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_191
timestamp 1621261055
transform 1 0 19488 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_194
timestamp 1621261055
transform 1 0 19776 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_202
timestamp 1621261055
transform 1 0 20544 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_210
timestamp 1621261055
transform 1 0 21312 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_218
timestamp 1621261055
transform 1 0 22080 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_226
timestamp 1621261055
transform 1 0 22848 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_556
timestamp 1621261055
transform 1 0 24960 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_234
timestamp 1621261055
transform 1 0 23616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_242
timestamp 1621261055
transform 1 0 24384 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_246
timestamp 1621261055
transform 1 0 24768 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_249
timestamp 1621261055
transform 1 0 25056 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_257
timestamp 1621261055
transform 1 0 25824 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_265
timestamp 1621261055
transform 1 0 26592 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_273
timestamp 1621261055
transform 1 0 27360 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_281
timestamp 1621261055
transform 1 0 28128 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_289
timestamp 1621261055
transform 1 0 28896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_297
timestamp 1621261055
transform 1 0 29664 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_557
timestamp 1621261055
transform 1 0 30240 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_301
timestamp 1621261055
transform 1 0 30048 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_304
timestamp 1621261055
transform 1 0 30336 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_312
timestamp 1621261055
transform 1 0 31104 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_320
timestamp 1621261055
transform 1 0 31872 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_328
timestamp 1621261055
transform 1 0 32640 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_558
timestamp 1621261055
transform 1 0 35520 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_336
timestamp 1621261055
transform 1 0 33408 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_344
timestamp 1621261055
transform 1 0 34176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_352
timestamp 1621261055
transform 1 0 34944 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_356
timestamp 1621261055
transform 1 0 35328 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_359
timestamp 1621261055
transform 1 0 35616 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_367
timestamp 1621261055
transform 1 0 36384 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_375
timestamp 1621261055
transform 1 0 37152 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_383
timestamp 1621261055
transform 1 0 37920 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_391
timestamp 1621261055
transform 1 0 38688 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_559
timestamp 1621261055
transform 1 0 40800 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_399
timestamp 1621261055
transform 1 0 39456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_407
timestamp 1621261055
transform 1 0 40224 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_411
timestamp 1621261055
transform 1 0 40608 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_414
timestamp 1621261055
transform 1 0 40896 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_422
timestamp 1621261055
transform 1 0 41664 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_430
timestamp 1621261055
transform 1 0 42432 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_438
timestamp 1621261055
transform 1 0 43200 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_446
timestamp 1621261055
transform 1 0 43968 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_454
timestamp 1621261055
transform 1 0 44736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_462
timestamp 1621261055
transform 1 0 45504 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_560
timestamp 1621261055
transform 1 0 46080 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_466
timestamp 1621261055
transform 1 0 45888 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_469
timestamp 1621261055
transform 1 0 46176 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_477
timestamp 1621261055
transform 1 0 46944 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_485
timestamp 1621261055
transform 1 0 47712 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_493
timestamp 1621261055
transform 1 0 48480 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_561
timestamp 1621261055
transform 1 0 51360 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_501
timestamp 1621261055
transform 1 0 49248 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_509
timestamp 1621261055
transform 1 0 50016 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_517
timestamp 1621261055
transform 1 0 50784 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_521
timestamp 1621261055
transform 1 0 51168 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_524
timestamp 1621261055
transform 1 0 51456 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_532
timestamp 1621261055
transform 1 0 52224 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_540
timestamp 1621261055
transform 1 0 52992 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_548
timestamp 1621261055
transform 1 0 53760 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_556
timestamp 1621261055
transform 1 0 54528 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_562
timestamp 1621261055
transform 1 0 56640 0 -1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_36_564
timestamp 1621261055
transform 1 0 55296 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_36_572
timestamp 1621261055
transform 1 0 56064 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_576
timestamp 1621261055
transform 1 0 56448 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_36_579
timestamp 1621261055
transform 1 0 56736 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_36_587
timestamp 1621261055
transform 1 0 57504 0 -1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_73
timestamp 1621261055
transform -1 0 58848 0 -1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_36_595
timestamp 1621261055
transform 1 0 58272 0 -1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_74
timestamp 1621261055
transform 1 0 1152 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_4
timestamp 1621261055
transform 1 0 1536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_12
timestamp 1621261055
transform 1 0 2304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_20
timestamp 1621261055
transform 1 0 3072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_28
timestamp 1621261055
transform 1 0 3840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_563
timestamp 1621261055
transform 1 0 6432 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_36
timestamp 1621261055
transform 1 0 4608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_44
timestamp 1621261055
transform 1 0 5376 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_52
timestamp 1621261055
transform 1 0 6144 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_54
timestamp 1621261055
transform 1 0 6336 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_56
timestamp 1621261055
transform 1 0 6528 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_64
timestamp 1621261055
transform 1 0 7296 0 1 27306
box -38 -49 422 715
use OR2X1  OR2X1
timestamp 1623617396
transform 1 0 7680 0 1 27306
box 0 -48 1152 714
use sky130_fd_sc_ls__decap_8  FILLER_37_80
timestamp 1621261055
transform 1 0 8832 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_88
timestamp 1621261055
transform 1 0 9600 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_96
timestamp 1621261055
transform 1 0 10368 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_564
timestamp 1621261055
transform 1 0 11712 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_104
timestamp 1621261055
transform 1 0 11136 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_108
timestamp 1621261055
transform 1 0 11520 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_111
timestamp 1621261055
transform 1 0 11808 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_119
timestamp 1621261055
transform 1 0 12576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_127
timestamp 1621261055
transform 1 0 13344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _158_
timestamp 1621261055
transform 1 0 16032 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_565
timestamp 1621261055
transform 1 0 16992 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_135
timestamp 1621261055
transform 1 0 14112 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_143
timestamp 1621261055
transform 1 0 14880 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_151
timestamp 1621261055
transform 1 0 15648 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_37_158
timestamp 1621261055
transform 1 0 16320 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_162
timestamp 1621261055
transform 1 0 16704 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_164
timestamp 1621261055
transform 1 0 16896 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_166
timestamp 1621261055
transform 1 0 17088 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_174
timestamp 1621261055
transform 1 0 17856 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_182
timestamp 1621261055
transform 1 0 18624 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_190
timestamp 1621261055
transform 1 0 19392 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_198
timestamp 1621261055
transform 1 0 20160 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _166_
timestamp 1621261055
transform 1 0 22752 0 1 27306
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_566
timestamp 1621261055
transform 1 0 22272 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_206
timestamp 1621261055
transform 1 0 20928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_214
timestamp 1621261055
transform 1 0 21696 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_218
timestamp 1621261055
transform 1 0 22080 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_37_221
timestamp 1621261055
transform 1 0 22368 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_37_228
timestamp 1621261055
transform 1 0 23040 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_236
timestamp 1621261055
transform 1 0 23808 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_244
timestamp 1621261055
transform 1 0 24576 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_252
timestamp 1621261055
transform 1 0 25344 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_260
timestamp 1621261055
transform 1 0 26112 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_567
timestamp 1621261055
transform 1 0 27552 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_268
timestamp 1621261055
transform 1 0 26880 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_272
timestamp 1621261055
transform 1 0 27264 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_37_274
timestamp 1621261055
transform 1 0 27456 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_276
timestamp 1621261055
transform 1 0 27648 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_284
timestamp 1621261055
transform 1 0 28416 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_292
timestamp 1621261055
transform 1 0 29184 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_568
timestamp 1621261055
transform 1 0 32832 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_300
timestamp 1621261055
transform 1 0 29952 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_308
timestamp 1621261055
transform 1 0 30720 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_316
timestamp 1621261055
transform 1 0 31488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_324
timestamp 1621261055
transform 1 0 32256 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_328
timestamp 1621261055
transform 1 0 32640 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_331
timestamp 1621261055
transform 1 0 32928 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_339
timestamp 1621261055
transform 1 0 33696 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_347
timestamp 1621261055
transform 1 0 34464 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_355
timestamp 1621261055
transform 1 0 35232 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_363
timestamp 1621261055
transform 1 0 36000 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_569
timestamp 1621261055
transform 1 0 38112 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_371
timestamp 1621261055
transform 1 0 36768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_379
timestamp 1621261055
transform 1 0 37536 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_383
timestamp 1621261055
transform 1 0 37920 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_386
timestamp 1621261055
transform 1 0 38208 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_394
timestamp 1621261055
transform 1 0 38976 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_402
timestamp 1621261055
transform 1 0 39744 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_410
timestamp 1621261055
transform 1 0 40512 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_418
timestamp 1621261055
transform 1 0 41280 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_426
timestamp 1621261055
transform 1 0 42048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_570
timestamp 1621261055
transform 1 0 43392 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_37_434
timestamp 1621261055
transform 1 0 42816 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_438
timestamp 1621261055
transform 1 0 43200 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_441
timestamp 1621261055
transform 1 0 43488 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_449
timestamp 1621261055
transform 1 0 44256 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_457
timestamp 1621261055
transform 1 0 45024 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_571
timestamp 1621261055
transform 1 0 48672 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_465
timestamp 1621261055
transform 1 0 45792 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_473
timestamp 1621261055
transform 1 0 46560 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_481
timestamp 1621261055
transform 1 0 47328 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_489
timestamp 1621261055
transform 1 0 48096 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_493
timestamp 1621261055
transform 1 0 48480 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_496
timestamp 1621261055
transform 1 0 48768 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_504
timestamp 1621261055
transform 1 0 49536 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_512
timestamp 1621261055
transform 1 0 50304 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_520
timestamp 1621261055
transform 1 0 51072 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_528
timestamp 1621261055
transform 1 0 51840 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_572
timestamp 1621261055
transform 1 0 53952 0 1 27306
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_37_536
timestamp 1621261055
transform 1 0 52608 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_544
timestamp 1621261055
transform 1 0 53376 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_548
timestamp 1621261055
transform 1 0 53760 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_37_551
timestamp 1621261055
transform 1 0 54048 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_559
timestamp 1621261055
transform 1 0 54816 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_567
timestamp 1621261055
transform 1 0 55584 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_575
timestamp 1621261055
transform 1 0 56352 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_37_583
timestamp 1621261055
transform 1 0 57120 0 1 27306
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_37_591
timestamp 1621261055
transform 1 0 57888 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_75
timestamp 1621261055
transform -1 0 58848 0 1 27306
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_37_595
timestamp 1621261055
transform 1 0 58272 0 1 27306
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_39_4
timestamp 1621261055
transform 1 0 1536 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_4
timestamp 1621261055
transform 1 0 1536 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_6
timestamp 1621261055
transform -1 0 1824 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_78
timestamp 1621261055
transform 1 0 1152 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_76
timestamp 1621261055
transform 1 0 1152 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _002_
timestamp 1621261055
transform -1 0 2112 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_10
timestamp 1621261055
transform 1 0 2112 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_12
timestamp 1621261055
transform 1 0 2304 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_26
timestamp 1621261055
transform 1 0 3648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_18
timestamp 1621261055
transform 1 0 2880 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_20
timestamp 1621261055
transform 1 0 3072 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_29
timestamp 1621261055
transform 1 0 3936 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_573
timestamp 1621261055
transform 1 0 3840 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_34
timestamp 1621261055
transform 1 0 4416 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_37
timestamp 1621261055
transform 1 0 4704 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_50
timestamp 1621261055
transform 1 0 5952 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_42
timestamp 1621261055
transform 1 0 5184 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_45
timestamp 1621261055
transform 1 0 5472 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_56
timestamp 1621261055
transform 1 0 6528 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_54
timestamp 1621261055
transform 1 0 6336 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_53
timestamp 1621261055
transform 1 0 6240 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_584
timestamp 1621261055
transform 1 0 6432 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_39_64
timestamp 1621261055
transform 1 0 7296 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_61
timestamp 1621261055
transform 1 0 7008 0 -1 28638
box -38 -49 806 715
use XNOR2X1  XNOR2X1
timestamp 1623617396
transform 1 0 7680 0 1 28638
box 0 -48 2016 714
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_574
timestamp 1621261055
transform 1 0 9120 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_69
timestamp 1621261055
transform 1 0 7776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_77
timestamp 1621261055
transform 1 0 8544 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_81
timestamp 1621261055
transform 1 0 8928 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_84
timestamp 1621261055
transform 1 0 9216 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_92
timestamp 1621261055
transform 1 0 9984 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_89
timestamp 1621261055
transform 1 0 9696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_97
timestamp 1621261055
transform 1 0 10464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_105
timestamp 1621261055
transform 1 0 11232 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_100
timestamp 1621261055
transform 1 0 10752 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_111
timestamp 1621261055
transform 1 0 11808 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_109
timestamp 1621261055
transform 1 0 11616 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_116
timestamp 1621261055
transform 1 0 12288 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_108
timestamp 1621261055
transform 1 0 11520 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_585
timestamp 1621261055
transform 1 0 11712 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_119
timestamp 1621261055
transform 1 0 12576 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_124
timestamp 1621261055
transform 1 0 13056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_127
timestamp 1621261055
transform 1 0 13344 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_132
timestamp 1621261055
transform 1 0 13824 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_135
timestamp 1621261055
transform 1 0 14112 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_139
timestamp 1621261055
transform 1 0 14496 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_136
timestamp 1621261055
transform 1 0 14208 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_575
timestamp 1621261055
transform 1 0 14400 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_143
timestamp 1621261055
transform 1 0 14880 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_147
timestamp 1621261055
transform 1 0 15264 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_151
timestamp 1621261055
transform 1 0 15648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_155
timestamp 1621261055
transform 1 0 16032 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_163
timestamp 1621261055
transform 1 0 16800 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_159
timestamp 1621261055
transform 1 0 16416 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_163
timestamp 1621261055
transform 1 0 16800 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_586
timestamp 1621261055
transform 1 0 16992 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_166
timestamp 1621261055
transform 1 0 17088 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_171
timestamp 1621261055
transform 1 0 17568 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_182
timestamp 1621261055
transform 1 0 18624 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_174
timestamp 1621261055
transform 1 0 17856 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_179
timestamp 1621261055
transform 1 0 18336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_190
timestamp 1621261055
transform 1 0 19392 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_191
timestamp 1621261055
transform 1 0 19488 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_187
timestamp 1621261055
transform 1 0 19104 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_198
timestamp 1621261055
transform 1 0 20160 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_194
timestamp 1621261055
transform 1 0 19776 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_576
timestamp 1621261055
transform 1 0 19680 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_206
timestamp 1621261055
transform 1 0 20928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_202
timestamp 1621261055
transform 1 0 20544 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_214
timestamp 1621261055
transform 1 0 21696 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_210
timestamp 1621261055
transform 1 0 21312 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_221
timestamp 1621261055
transform 1 0 22368 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_218
timestamp 1621261055
transform 1 0 22080 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_38_220
timestamp 1621261055
transform 1 0 22272 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_218
timestamp 1621261055
transform 1 0 22080 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_35
timestamp 1621261055
transform -1 0 22560 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_587
timestamp 1621261055
transform 1 0 22272 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _035_
timestamp 1621261055
transform -1 0 22848 0 -1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_229
timestamp 1621261055
transform 1 0 23136 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_226
timestamp 1621261055
transform 1 0 22848 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_237
timestamp 1621261055
transform 1 0 23904 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_234
timestamp 1621261055
transform 1 0 23616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_245
timestamp 1621261055
transform 1 0 24672 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_246
timestamp 1621261055
transform 1 0 24768 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_242
timestamp 1621261055
transform 1 0 24384 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_577
timestamp 1621261055
transform 1 0 24960 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_253
timestamp 1621261055
transform 1 0 25440 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_257
timestamp 1621261055
transform 1 0 25824 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_249
timestamp 1621261055
transform 1 0 25056 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_261
timestamp 1621261055
transform 1 0 26208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_269
timestamp 1621261055
transform 1 0 26976 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_265
timestamp 1621261055
transform 1 0 26592 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_276
timestamp 1621261055
transform 1 0 27648 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_273
timestamp 1621261055
transform 1 0 27360 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_281
timestamp 1621261055
transform 1 0 28128 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_273
timestamp 1621261055
transform 1 0 27360 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_588
timestamp 1621261055
transform 1 0 27552 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_284
timestamp 1621261055
transform 1 0 28416 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_289
timestamp 1621261055
transform 1 0 28896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_292
timestamp 1621261055
transform 1 0 29184 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_297
timestamp 1621261055
transform 1 0 29664 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_300
timestamp 1621261055
transform 1 0 29952 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_304
timestamp 1621261055
transform 1 0 30336 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_301
timestamp 1621261055
transform 1 0 30048 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_578
timestamp 1621261055
transform 1 0 30240 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_308
timestamp 1621261055
transform 1 0 30720 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_312
timestamp 1621261055
transform 1 0 31104 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_316
timestamp 1621261055
transform 1 0 31488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_320
timestamp 1621261055
transform 1 0 31872 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_328
timestamp 1621261055
transform 1 0 32640 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_324
timestamp 1621261055
transform 1 0 32256 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_328
timestamp 1621261055
transform 1 0 32640 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_589
timestamp 1621261055
transform 1 0 32832 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_331
timestamp 1621261055
transform 1 0 32928 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_336
timestamp 1621261055
transform 1 0 33408 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_347
timestamp 1621261055
transform 1 0 34464 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_339
timestamp 1621261055
transform 1 0 33696 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_344
timestamp 1621261055
transform 1 0 34176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_355
timestamp 1621261055
transform 1 0 35232 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_356
timestamp 1621261055
transform 1 0 35328 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_352
timestamp 1621261055
transform 1 0 34944 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_363
timestamp 1621261055
transform 1 0 36000 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_359
timestamp 1621261055
transform 1 0 35616 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_579
timestamp 1621261055
transform 1 0 35520 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_371
timestamp 1621261055
transform 1 0 36768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_367
timestamp 1621261055
transform 1 0 36384 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_379
timestamp 1621261055
transform 1 0 37536 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_375
timestamp 1621261055
transform 1 0 37152 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_386
timestamp 1621261055
transform 1 0 38208 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_383
timestamp 1621261055
transform 1 0 37920 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_383
timestamp 1621261055
transform 1 0 37920 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_590
timestamp 1621261055
transform 1 0 38112 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_394
timestamp 1621261055
transform 1 0 38976 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_391
timestamp 1621261055
transform 1 0 38688 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_402
timestamp 1621261055
transform 1 0 39744 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_399
timestamp 1621261055
transform 1 0 39456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_410
timestamp 1621261055
transform 1 0 40512 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_411
timestamp 1621261055
transform 1 0 40608 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_407
timestamp 1621261055
transform 1 0 40224 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_580
timestamp 1621261055
transform 1 0 40800 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_418
timestamp 1621261055
transform 1 0 41280 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_422
timestamp 1621261055
transform 1 0 41664 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_414
timestamp 1621261055
transform 1 0 40896 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_426
timestamp 1621261055
transform 1 0 42048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_434
timestamp 1621261055
transform 1 0 42816 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_430
timestamp 1621261055
transform 1 0 42432 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_441
timestamp 1621261055
transform 1 0 43488 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_438
timestamp 1621261055
transform 1 0 43200 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_38_446
timestamp 1621261055
transform 1 0 43968 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_438
timestamp 1621261055
transform 1 0 43200 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_591
timestamp 1621261055
transform 1 0 43392 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_39_453
timestamp 1621261055
transform 1 0 44640 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_39_449
timestamp 1621261055
transform 1 0 44256 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_454
timestamp 1621261055
transform 1 0 44736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _124_
timestamp 1621261055
transform 1 0 44736 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_457
timestamp 1621261055
transform 1 0 45024 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_38_462
timestamp 1621261055
transform 1 0 45504 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_465
timestamp 1621261055
transform 1 0 45792 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_469
timestamp 1621261055
transform 1 0 46176 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_466
timestamp 1621261055
transform 1 0 45888 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_581
timestamp 1621261055
transform 1 0 46080 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_473
timestamp 1621261055
transform 1 0 46560 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_477
timestamp 1621261055
transform 1 0 46944 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_481
timestamp 1621261055
transform 1 0 47328 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_485
timestamp 1621261055
transform 1 0 47712 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_493
timestamp 1621261055
transform 1 0 48480 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_489
timestamp 1621261055
transform 1 0 48096 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_493
timestamp 1621261055
transform 1 0 48480 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_592
timestamp 1621261055
transform 1 0 48672 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_496
timestamp 1621261055
transform 1 0 48768 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_501
timestamp 1621261055
transform 1 0 49248 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_508
timestamp 1621261055
transform 1 0 49920 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_39_504
timestamp 1621261055
transform 1 0 49536 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_509
timestamp 1621261055
transform 1 0 50016 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _103_
timestamp 1621261055
transform 1 0 50112 0 1 28638
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_39_521
timestamp 1621261055
transform 1 0 51168 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_513
timestamp 1621261055
transform 1 0 50400 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_521
timestamp 1621261055
transform 1 0 51168 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_517
timestamp 1621261055
transform 1 0 50784 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_38_524
timestamp 1621261055
transform 1 0 51456 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_582
timestamp 1621261055
transform 1 0 51360 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_529
timestamp 1621261055
transform 1 0 51936 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_532
timestamp 1621261055
transform 1 0 52224 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_545
timestamp 1621261055
transform 1 0 53472 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_39_537
timestamp 1621261055
transform 1 0 52704 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_540
timestamp 1621261055
transform 1 0 52992 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_551
timestamp 1621261055
transform 1 0 54048 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_39_549
timestamp 1621261055
transform 1 0 53856 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_38_548
timestamp 1621261055
transform 1 0 53760 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_593
timestamp 1621261055
transform 1 0 53952 0 1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_559
timestamp 1621261055
transform 1 0 54816 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_556
timestamp 1621261055
transform 1 0 54528 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_567
timestamp 1621261055
transform 1 0 55584 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_564
timestamp 1621261055
transform 1 0 55296 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_39_575
timestamp 1621261055
transform 1 0 56352 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_576
timestamp 1621261055
transform 1 0 56448 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_38_572
timestamp 1621261055
transform 1 0 56064 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_583
timestamp 1621261055
transform 1 0 56640 0 -1 28638
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_39_583
timestamp 1621261055
transform 1 0 57120 0 1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_587
timestamp 1621261055
transform 1 0 57504 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_38_579
timestamp 1621261055
transform 1 0 56736 0 -1 28638
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_39_591
timestamp 1621261055
transform 1 0 57888 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_77
timestamp 1621261055
transform -1 0 58848 0 -1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_79
timestamp 1621261055
transform -1 0 58848 0 1 28638
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_38_595
timestamp 1621261055
transform 1 0 58272 0 -1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_39_595
timestamp 1621261055
transform 1 0 58272 0 1 28638
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_80
timestamp 1621261055
transform 1 0 1152 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_594
timestamp 1621261055
transform 1 0 3840 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_4
timestamp 1621261055
transform 1 0 1536 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_12
timestamp 1621261055
transform 1 0 2304 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_20
timestamp 1621261055
transform 1 0 3072 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_29
timestamp 1621261055
transform 1 0 3936 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_37
timestamp 1621261055
transform 1 0 4704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_45
timestamp 1621261055
transform 1 0 5472 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_53
timestamp 1621261055
transform 1 0 6240 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_61
timestamp 1621261055
transform 1 0 7008 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_595
timestamp 1621261055
transform 1 0 9120 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_69
timestamp 1621261055
transform 1 0 7776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_77
timestamp 1621261055
transform 1 0 8544 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_81
timestamp 1621261055
transform 1 0 8928 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_84
timestamp 1621261055
transform 1 0 9216 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_92
timestamp 1621261055
transform 1 0 9984 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _140_
timestamp 1621261055
transform 1 0 12768 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_40_100
timestamp 1621261055
transform 1 0 10752 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_108
timestamp 1621261055
transform 1 0 11520 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_116
timestamp 1621261055
transform 1 0 12288 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_40_120
timestamp 1621261055
transform 1 0 12672 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_124
timestamp 1621261055
transform 1 0 13056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_132
timestamp 1621261055
transform 1 0 13824 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _047_
timestamp 1621261055
transform 1 0 14880 0 -1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_596
timestamp 1621261055
transform 1 0 14400 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_49
timestamp 1621261055
transform 1 0 14688 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_136
timestamp 1621261055
transform 1 0 14208 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_139
timestamp 1621261055
transform 1 0 14496 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_146
timestamp 1621261055
transform 1 0 15168 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_154
timestamp 1621261055
transform 1 0 15936 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_162
timestamp 1621261055
transform 1 0 16704 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_597
timestamp 1621261055
transform 1 0 19680 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_170
timestamp 1621261055
transform 1 0 17472 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_178
timestamp 1621261055
transform 1 0 18240 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_186
timestamp 1621261055
transform 1 0 19008 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_190
timestamp 1621261055
transform 1 0 19392 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_40_192
timestamp 1621261055
transform 1 0 19584 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_194
timestamp 1621261055
transform 1 0 19776 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_202
timestamp 1621261055
transform 1 0 20544 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_210
timestamp 1621261055
transform 1 0 21312 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_218
timestamp 1621261055
transform 1 0 22080 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_226
timestamp 1621261055
transform 1 0 22848 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_598
timestamp 1621261055
transform 1 0 24960 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_234
timestamp 1621261055
transform 1 0 23616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_242
timestamp 1621261055
transform 1 0 24384 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_246
timestamp 1621261055
transform 1 0 24768 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_249
timestamp 1621261055
transform 1 0 25056 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_257
timestamp 1621261055
transform 1 0 25824 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_265
timestamp 1621261055
transform 1 0 26592 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_273
timestamp 1621261055
transform 1 0 27360 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_281
timestamp 1621261055
transform 1 0 28128 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_289
timestamp 1621261055
transform 1 0 28896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_297
timestamp 1621261055
transform 1 0 29664 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_599
timestamp 1621261055
transform 1 0 30240 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_301
timestamp 1621261055
transform 1 0 30048 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_304
timestamp 1621261055
transform 1 0 30336 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_312
timestamp 1621261055
transform 1 0 31104 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_320
timestamp 1621261055
transform 1 0 31872 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_328
timestamp 1621261055
transform 1 0 32640 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_600
timestamp 1621261055
transform 1 0 35520 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_336
timestamp 1621261055
transform 1 0 33408 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_344
timestamp 1621261055
transform 1 0 34176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_352
timestamp 1621261055
transform 1 0 34944 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_356
timestamp 1621261055
transform 1 0 35328 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_359
timestamp 1621261055
transform 1 0 35616 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_367
timestamp 1621261055
transform 1 0 36384 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_375
timestamp 1621261055
transform 1 0 37152 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_383
timestamp 1621261055
transform 1 0 37920 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_391
timestamp 1621261055
transform 1 0 38688 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_601
timestamp 1621261055
transform 1 0 40800 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_399
timestamp 1621261055
transform 1 0 39456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_407
timestamp 1621261055
transform 1 0 40224 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_411
timestamp 1621261055
transform 1 0 40608 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_414
timestamp 1621261055
transform 1 0 40896 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_422
timestamp 1621261055
transform 1 0 41664 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_430
timestamp 1621261055
transform 1 0 42432 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_438
timestamp 1621261055
transform 1 0 43200 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_446
timestamp 1621261055
transform 1 0 43968 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_454
timestamp 1621261055
transform 1 0 44736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_462
timestamp 1621261055
transform 1 0 45504 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_602
timestamp 1621261055
transform 1 0 46080 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_466
timestamp 1621261055
transform 1 0 45888 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_469
timestamp 1621261055
transform 1 0 46176 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_477
timestamp 1621261055
transform 1 0 46944 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_485
timestamp 1621261055
transform 1 0 47712 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_493
timestamp 1621261055
transform 1 0 48480 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_603
timestamp 1621261055
transform 1 0 51360 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_501
timestamp 1621261055
transform 1 0 49248 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_509
timestamp 1621261055
transform 1 0 50016 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_517
timestamp 1621261055
transform 1 0 50784 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_521
timestamp 1621261055
transform 1 0 51168 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_524
timestamp 1621261055
transform 1 0 51456 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_532
timestamp 1621261055
transform 1 0 52224 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_540
timestamp 1621261055
transform 1 0 52992 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_548
timestamp 1621261055
transform 1 0 53760 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_556
timestamp 1621261055
transform 1 0 54528 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_604
timestamp 1621261055
transform 1 0 56640 0 -1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_40_564
timestamp 1621261055
transform 1 0 55296 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_40_572
timestamp 1621261055
transform 1 0 56064 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_576
timestamp 1621261055
transform 1 0 56448 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_40_579
timestamp 1621261055
transform 1 0 56736 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_40_587
timestamp 1621261055
transform 1 0 57504 0 -1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_81
timestamp 1621261055
transform -1 0 58848 0 -1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_40_595
timestamp 1621261055
transform 1 0 58272 0 -1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_82
timestamp 1621261055
transform 1 0 1152 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_4
timestamp 1621261055
transform 1 0 1536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_12
timestamp 1621261055
transform 1 0 2304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_20
timestamp 1621261055
transform 1 0 3072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_28
timestamp 1621261055
transform 1 0 3840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _008_
timestamp 1621261055
transform -1 0 7392 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_605
timestamp 1621261055
transform 1 0 6432 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_20
timestamp 1621261055
transform -1 0 7104 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_36
timestamp 1621261055
transform 1 0 4608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_44
timestamp 1621261055
transform 1 0 5376 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_52
timestamp 1621261055
transform 1 0 6144 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_41_54
timestamp 1621261055
transform 1 0 6336 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_56
timestamp 1621261055
transform 1 0 6528 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_41_65
timestamp 1621261055
transform 1 0 7392 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_73
timestamp 1621261055
transform 1 0 8160 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_81
timestamp 1621261055
transform 1 0 8928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_89
timestamp 1621261055
transform 1 0 9696 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_97
timestamp 1621261055
transform 1 0 10464 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_606
timestamp 1621261055
transform 1 0 11712 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_105
timestamp 1621261055
transform 1 0 11232 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_41_109
timestamp 1621261055
transform 1 0 11616 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_111
timestamp 1621261055
transform 1 0 11808 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_119
timestamp 1621261055
transform 1 0 12576 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_127
timestamp 1621261055
transform 1 0 13344 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_607
timestamp 1621261055
transform 1 0 16992 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_135
timestamp 1621261055
transform 1 0 14112 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_143
timestamp 1621261055
transform 1 0 14880 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_151
timestamp 1621261055
transform 1 0 15648 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_159
timestamp 1621261055
transform 1 0 16416 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_163
timestamp 1621261055
transform 1 0 16800 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_166
timestamp 1621261055
transform 1 0 17088 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_174
timestamp 1621261055
transform 1 0 17856 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_182
timestamp 1621261055
transform 1 0 18624 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_190
timestamp 1621261055
transform 1 0 19392 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_198
timestamp 1621261055
transform 1 0 20160 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_608
timestamp 1621261055
transform 1 0 22272 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_206
timestamp 1621261055
transform 1 0 20928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_214
timestamp 1621261055
transform 1 0 21696 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_218
timestamp 1621261055
transform 1 0 22080 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_221
timestamp 1621261055
transform 1 0 22368 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_229
timestamp 1621261055
transform 1 0 23136 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_237
timestamp 1621261055
transform 1 0 23904 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_245
timestamp 1621261055
transform 1 0 24672 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_253
timestamp 1621261055
transform 1 0 25440 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_261
timestamp 1621261055
transform 1 0 26208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _138_
timestamp 1621261055
transform 1 0 28128 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_609
timestamp 1621261055
transform 1 0 27552 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_269
timestamp 1621261055
transform 1 0 26976 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_273
timestamp 1621261055
transform 1 0 27360 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_41_276
timestamp 1621261055
transform 1 0 27648 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_41_280
timestamp 1621261055
transform 1 0 28032 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_284
timestamp 1621261055
transform 1 0 28416 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_292
timestamp 1621261055
transform 1 0 29184 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _196_
timestamp 1621261055
transform 1 0 31968 0 1 29970
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_610
timestamp 1621261055
transform 1 0 32832 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_300
timestamp 1621261055
transform 1 0 29952 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_308
timestamp 1621261055
transform 1 0 30720 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_316
timestamp 1621261055
transform 1 0 31488 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_41_320
timestamp 1621261055
transform 1 0 31872 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_324
timestamp 1621261055
transform 1 0 32256 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_328
timestamp 1621261055
transform 1 0 32640 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_331
timestamp 1621261055
transform 1 0 32928 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_339
timestamp 1621261055
transform 1 0 33696 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_347
timestamp 1621261055
transform 1 0 34464 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_355
timestamp 1621261055
transform 1 0 35232 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_363
timestamp 1621261055
transform 1 0 36000 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_611
timestamp 1621261055
transform 1 0 38112 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_371
timestamp 1621261055
transform 1 0 36768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_379
timestamp 1621261055
transform 1 0 37536 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_383
timestamp 1621261055
transform 1 0 37920 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_386
timestamp 1621261055
transform 1 0 38208 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_394
timestamp 1621261055
transform 1 0 38976 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_402
timestamp 1621261055
transform 1 0 39744 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_410
timestamp 1621261055
transform 1 0 40512 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_418
timestamp 1621261055
transform 1 0 41280 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_426
timestamp 1621261055
transform 1 0 42048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_612
timestamp 1621261055
transform 1 0 43392 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_41_434
timestamp 1621261055
transform 1 0 42816 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_438
timestamp 1621261055
transform 1 0 43200 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_441
timestamp 1621261055
transform 1 0 43488 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_449
timestamp 1621261055
transform 1 0 44256 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_457
timestamp 1621261055
transform 1 0 45024 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_613
timestamp 1621261055
transform 1 0 48672 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_465
timestamp 1621261055
transform 1 0 45792 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_473
timestamp 1621261055
transform 1 0 46560 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_481
timestamp 1621261055
transform 1 0 47328 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_489
timestamp 1621261055
transform 1 0 48096 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_493
timestamp 1621261055
transform 1 0 48480 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_496
timestamp 1621261055
transform 1 0 48768 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_504
timestamp 1621261055
transform 1 0 49536 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_512
timestamp 1621261055
transform 1 0 50304 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_520
timestamp 1621261055
transform 1 0 51072 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_528
timestamp 1621261055
transform 1 0 51840 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_614
timestamp 1621261055
transform 1 0 53952 0 1 29970
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_41_536
timestamp 1621261055
transform 1 0 52608 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_544
timestamp 1621261055
transform 1 0 53376 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_548
timestamp 1621261055
transform 1 0 53760 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_41_551
timestamp 1621261055
transform 1 0 54048 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_559
timestamp 1621261055
transform 1 0 54816 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_567
timestamp 1621261055
transform 1 0 55584 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_575
timestamp 1621261055
transform 1 0 56352 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_41_583
timestamp 1621261055
transform 1 0 57120 0 1 29970
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_41_591
timestamp 1621261055
transform 1 0 57888 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_83
timestamp 1621261055
transform -1 0 58848 0 1 29970
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_41_595
timestamp 1621261055
transform 1 0 58272 0 1 29970
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_84
timestamp 1621261055
transform 1 0 1152 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_615
timestamp 1621261055
transform 1 0 3840 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_4
timestamp 1621261055
transform 1 0 1536 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_12
timestamp 1621261055
transform 1 0 2304 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_20
timestamp 1621261055
transform 1 0 3072 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_29
timestamp 1621261055
transform 1 0 3936 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _202_
timestamp 1621261055
transform 1 0 6432 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_37
timestamp 1621261055
transform 1 0 4704 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_45
timestamp 1621261055
transform 1 0 5472 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_53
timestamp 1621261055
transform 1 0 6240 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_58
timestamp 1621261055
transform 1 0 6720 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_66
timestamp 1621261055
transform 1 0 7488 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_616
timestamp 1621261055
transform 1 0 9120 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_74
timestamp 1621261055
transform 1 0 8256 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_42_82
timestamp 1621261055
transform 1 0 9024 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_84
timestamp 1621261055
transform 1 0 9216 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_92
timestamp 1621261055
transform 1 0 9984 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _163_
timestamp 1621261055
transform 1 0 11520 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_100
timestamp 1621261055
transform 1 0 10752 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_111
timestamp 1621261055
transform 1 0 11808 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_119
timestamp 1621261055
transform 1 0 12576 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_127
timestamp 1621261055
transform 1 0 13344 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_617
timestamp 1621261055
transform 1 0 14400 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_135
timestamp 1621261055
transform 1 0 14112 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_42_137
timestamp 1621261055
transform 1 0 14304 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_139
timestamp 1621261055
transform 1 0 14496 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_147
timestamp 1621261055
transform 1 0 15264 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_155
timestamp 1621261055
transform 1 0 16032 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_163
timestamp 1621261055
transform 1 0 16800 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_618
timestamp 1621261055
transform 1 0 19680 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_171
timestamp 1621261055
transform 1 0 17568 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_179
timestamp 1621261055
transform 1 0 18336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_187
timestamp 1621261055
transform 1 0 19104 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_191
timestamp 1621261055
transform 1 0 19488 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_194
timestamp 1621261055
transform 1 0 19776 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_202
timestamp 1621261055
transform 1 0 20544 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_210
timestamp 1621261055
transform 1 0 21312 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_218
timestamp 1621261055
transform 1 0 22080 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_226
timestamp 1621261055
transform 1 0 22848 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_619
timestamp 1621261055
transform 1 0 24960 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_234
timestamp 1621261055
transform 1 0 23616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_242
timestamp 1621261055
transform 1 0 24384 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_246
timestamp 1621261055
transform 1 0 24768 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_249
timestamp 1621261055
transform 1 0 25056 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_257
timestamp 1621261055
transform 1 0 25824 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _110_
timestamp 1621261055
transform 1 0 27936 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_42_265
timestamp 1621261055
transform 1 0 26592 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_273
timestamp 1621261055
transform 1 0 27360 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_277
timestamp 1621261055
transform 1 0 27744 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_282
timestamp 1621261055
transform 1 0 28224 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_290
timestamp 1621261055
transform 1 0 28992 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_620
timestamp 1621261055
transform 1 0 30240 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_42_298
timestamp 1621261055
transform 1 0 29760 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_42_302
timestamp 1621261055
transform 1 0 30144 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_304
timestamp 1621261055
transform 1 0 30336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_312
timestamp 1621261055
transform 1 0 31104 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_320
timestamp 1621261055
transform 1 0 31872 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_328
timestamp 1621261055
transform 1 0 32640 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_621
timestamp 1621261055
transform 1 0 35520 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_336
timestamp 1621261055
transform 1 0 33408 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_344
timestamp 1621261055
transform 1 0 34176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_352
timestamp 1621261055
transform 1 0 34944 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_356
timestamp 1621261055
transform 1 0 35328 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_359
timestamp 1621261055
transform 1 0 35616 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_367
timestamp 1621261055
transform 1 0 36384 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_375
timestamp 1621261055
transform 1 0 37152 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_383
timestamp 1621261055
transform 1 0 37920 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_391
timestamp 1621261055
transform 1 0 38688 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _012_
timestamp 1621261055
transform 1 0 41280 0 -1 31302
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_622
timestamp 1621261055
transform 1 0 40800 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_399
timestamp 1621261055
transform 1 0 39456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_407
timestamp 1621261055
transform 1 0 40224 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_411
timestamp 1621261055
transform 1 0 40608 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_42_414
timestamp 1621261055
transform 1 0 40896 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_42_421
timestamp 1621261055
transform 1 0 41568 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_429
timestamp 1621261055
transform 1 0 42336 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_437
timestamp 1621261055
transform 1 0 43104 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_445
timestamp 1621261055
transform 1 0 43872 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_453
timestamp 1621261055
transform 1 0 44640 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_461
timestamp 1621261055
transform 1 0 45408 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_623
timestamp 1621261055
transform 1 0 46080 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_465
timestamp 1621261055
transform 1 0 45792 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_42_467
timestamp 1621261055
transform 1 0 45984 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_469
timestamp 1621261055
transform 1 0 46176 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_477
timestamp 1621261055
transform 1 0 46944 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_485
timestamp 1621261055
transform 1 0 47712 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_493
timestamp 1621261055
transform 1 0 48480 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_624
timestamp 1621261055
transform 1 0 51360 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_501
timestamp 1621261055
transform 1 0 49248 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_509
timestamp 1621261055
transform 1 0 50016 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_517
timestamp 1621261055
transform 1 0 50784 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_521
timestamp 1621261055
transform 1 0 51168 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_524
timestamp 1621261055
transform 1 0 51456 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_532
timestamp 1621261055
transform 1 0 52224 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_540
timestamp 1621261055
transform 1 0 52992 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_548
timestamp 1621261055
transform 1 0 53760 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_556
timestamp 1621261055
transform 1 0 54528 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_625
timestamp 1621261055
transform 1 0 56640 0 -1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_42_564
timestamp 1621261055
transform 1 0 55296 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_42_572
timestamp 1621261055
transform 1 0 56064 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_576
timestamp 1621261055
transform 1 0 56448 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_42_579
timestamp 1621261055
transform 1 0 56736 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_42_587
timestamp 1621261055
transform 1 0 57504 0 -1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_85
timestamp 1621261055
transform -1 0 58848 0 -1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_42_595
timestamp 1621261055
transform 1 0 58272 0 -1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_86
timestamp 1621261055
transform 1 0 1152 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_43_4
timestamp 1621261055
transform 1 0 1536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_12
timestamp 1621261055
transform 1 0 2304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_20
timestamp 1621261055
transform 1 0 3072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_28
timestamp 1621261055
transform 1 0 3840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_626
timestamp 1621261055
transform 1 0 6432 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_36
timestamp 1621261055
transform 1 0 4608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_44
timestamp 1621261055
transform 1 0 5376 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_52
timestamp 1621261055
transform 1 0 6144 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_43_54
timestamp 1621261055
transform 1 0 6336 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_56
timestamp 1621261055
transform 1 0 6528 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_64
timestamp 1621261055
transform 1 0 7296 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_72
timestamp 1621261055
transform 1 0 8064 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_80
timestamp 1621261055
transform 1 0 8832 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_88
timestamp 1621261055
transform 1 0 9600 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_96
timestamp 1621261055
transform 1 0 10368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_627
timestamp 1621261055
transform 1 0 11712 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_104
timestamp 1621261055
transform 1 0 11136 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_108
timestamp 1621261055
transform 1 0 11520 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_111
timestamp 1621261055
transform 1 0 11808 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_119
timestamp 1621261055
transform 1 0 12576 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_127
timestamp 1621261055
transform 1 0 13344 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_628
timestamp 1621261055
transform 1 0 16992 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_135
timestamp 1621261055
transform 1 0 14112 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_143
timestamp 1621261055
transform 1 0 14880 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_151
timestamp 1621261055
transform 1 0 15648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_159
timestamp 1621261055
transform 1 0 16416 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_163
timestamp 1621261055
transform 1 0 16800 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_166
timestamp 1621261055
transform 1 0 17088 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_174
timestamp 1621261055
transform 1 0 17856 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_182
timestamp 1621261055
transform 1 0 18624 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_190
timestamp 1621261055
transform 1 0 19392 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_198
timestamp 1621261055
transform 1 0 20160 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_629
timestamp 1621261055
transform 1 0 22272 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_206
timestamp 1621261055
transform 1 0 20928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_214
timestamp 1621261055
transform 1 0 21696 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_218
timestamp 1621261055
transform 1 0 22080 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_221
timestamp 1621261055
transform 1 0 22368 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_229
timestamp 1621261055
transform 1 0 23136 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_237
timestamp 1621261055
transform 1 0 23904 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_245
timestamp 1621261055
transform 1 0 24672 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_253
timestamp 1621261055
transform 1 0 25440 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_261
timestamp 1621261055
transform 1 0 26208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_630
timestamp 1621261055
transform 1 0 27552 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_269
timestamp 1621261055
transform 1 0 26976 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_273
timestamp 1621261055
transform 1 0 27360 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_276
timestamp 1621261055
transform 1 0 27648 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_284
timestamp 1621261055
transform 1 0 28416 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_292
timestamp 1621261055
transform 1 0 29184 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_631
timestamp 1621261055
transform 1 0 32832 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_300
timestamp 1621261055
transform 1 0 29952 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_308
timestamp 1621261055
transform 1 0 30720 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_316
timestamp 1621261055
transform 1 0 31488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_324
timestamp 1621261055
transform 1 0 32256 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_328
timestamp 1621261055
transform 1 0 32640 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_331
timestamp 1621261055
transform 1 0 32928 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_339
timestamp 1621261055
transform 1 0 33696 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_347
timestamp 1621261055
transform 1 0 34464 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_355
timestamp 1621261055
transform 1 0 35232 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_363
timestamp 1621261055
transform 1 0 36000 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_632
timestamp 1621261055
transform 1 0 38112 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_371
timestamp 1621261055
transform 1 0 36768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_379
timestamp 1621261055
transform 1 0 37536 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_383
timestamp 1621261055
transform 1 0 37920 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_386
timestamp 1621261055
transform 1 0 38208 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_394
timestamp 1621261055
transform 1 0 38976 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_402
timestamp 1621261055
transform 1 0 39744 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_410
timestamp 1621261055
transform 1 0 40512 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_418
timestamp 1621261055
transform 1 0 41280 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_426
timestamp 1621261055
transform 1 0 42048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_633
timestamp 1621261055
transform 1 0 43392 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_43_434
timestamp 1621261055
transform 1 0 42816 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_438
timestamp 1621261055
transform 1 0 43200 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_441
timestamp 1621261055
transform 1 0 43488 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_449
timestamp 1621261055
transform 1 0 44256 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_457
timestamp 1621261055
transform 1 0 45024 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_634
timestamp 1621261055
transform 1 0 48672 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_465
timestamp 1621261055
transform 1 0 45792 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_473
timestamp 1621261055
transform 1 0 46560 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_481
timestamp 1621261055
transform 1 0 47328 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_489
timestamp 1621261055
transform 1 0 48096 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_493
timestamp 1621261055
transform 1 0 48480 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_496
timestamp 1621261055
transform 1 0 48768 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_504
timestamp 1621261055
transform 1 0 49536 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_512
timestamp 1621261055
transform 1 0 50304 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_520
timestamp 1621261055
transform 1 0 51072 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_528
timestamp 1621261055
transform 1 0 51840 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_635
timestamp 1621261055
transform 1 0 53952 0 1 31302
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_43_536
timestamp 1621261055
transform 1 0 52608 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_544
timestamp 1621261055
transform 1 0 53376 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_548
timestamp 1621261055
transform 1 0 53760 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_43_551
timestamp 1621261055
transform 1 0 54048 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_559
timestamp 1621261055
transform 1 0 54816 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_567
timestamp 1621261055
transform 1 0 55584 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_575
timestamp 1621261055
transform 1 0 56352 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_43_583
timestamp 1621261055
transform 1 0 57120 0 1 31302
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_43_591
timestamp 1621261055
transform 1 0 57888 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_87
timestamp 1621261055
transform -1 0 58848 0 1 31302
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_43_595
timestamp 1621261055
transform 1 0 58272 0 1 31302
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_8
timestamp 1621261055
transform 1 0 1920 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_44_4
timestamp 1621261055
transform 1 0 1536 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_88
timestamp 1621261055
transform 1 0 1152 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_13
timestamp 1621261055
transform 1 0 2400 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _180_
timestamp 1621261055
transform 1 0 2112 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_25
timestamp 1621261055
transform 1 0 3552 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_44_21
timestamp 1621261055
transform 1 0 3168 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_44_29
timestamp 1621261055
transform 1 0 3936 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_44_27
timestamp 1621261055
transform 1 0 3744 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_636
timestamp 1621261055
transform 1 0 3840 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _170_
timestamp 1621261055
transform 1 0 6432 0 -1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_44_37
timestamp 1621261055
transform 1 0 4704 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_45
timestamp 1621261055
transform 1 0 5472 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_53
timestamp 1621261055
transform 1 0 6240 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_58
timestamp 1621261055
transform 1 0 6720 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_66
timestamp 1621261055
transform 1 0 7488 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_637
timestamp 1621261055
transform 1 0 9120 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_74
timestamp 1621261055
transform 1 0 8256 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_44_82
timestamp 1621261055
transform 1 0 9024 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_84
timestamp 1621261055
transform 1 0 9216 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_92
timestamp 1621261055
transform 1 0 9984 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_100
timestamp 1621261055
transform 1 0 10752 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_108
timestamp 1621261055
transform 1 0 11520 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_116
timestamp 1621261055
transform 1 0 12288 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_124
timestamp 1621261055
transform 1 0 13056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_132
timestamp 1621261055
transform 1 0 13824 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_638
timestamp 1621261055
transform 1 0 14400 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_136
timestamp 1621261055
transform 1 0 14208 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_139
timestamp 1621261055
transform 1 0 14496 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_147
timestamp 1621261055
transform 1 0 15264 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_155
timestamp 1621261055
transform 1 0 16032 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_163
timestamp 1621261055
transform 1 0 16800 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_639
timestamp 1621261055
transform 1 0 19680 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_171
timestamp 1621261055
transform 1 0 17568 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_179
timestamp 1621261055
transform 1 0 18336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_187
timestamp 1621261055
transform 1 0 19104 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_191
timestamp 1621261055
transform 1 0 19488 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_194
timestamp 1621261055
transform 1 0 19776 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_202
timestamp 1621261055
transform 1 0 20544 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_210
timestamp 1621261055
transform 1 0 21312 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_218
timestamp 1621261055
transform 1 0 22080 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_226
timestamp 1621261055
transform 1 0 22848 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_640
timestamp 1621261055
transform 1 0 24960 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_234
timestamp 1621261055
transform 1 0 23616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_242
timestamp 1621261055
transform 1 0 24384 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_246
timestamp 1621261055
transform 1 0 24768 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_249
timestamp 1621261055
transform 1 0 25056 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_257
timestamp 1621261055
transform 1 0 25824 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_265
timestamp 1621261055
transform 1 0 26592 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_273
timestamp 1621261055
transform 1 0 27360 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_281
timestamp 1621261055
transform 1 0 28128 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_289
timestamp 1621261055
transform 1 0 28896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_297
timestamp 1621261055
transform 1 0 29664 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_641
timestamp 1621261055
transform 1 0 30240 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_301
timestamp 1621261055
transform 1 0 30048 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_304
timestamp 1621261055
transform 1 0 30336 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_312
timestamp 1621261055
transform 1 0 31104 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_320
timestamp 1621261055
transform 1 0 31872 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_328
timestamp 1621261055
transform 1 0 32640 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_642
timestamp 1621261055
transform 1 0 35520 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_336
timestamp 1621261055
transform 1 0 33408 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_344
timestamp 1621261055
transform 1 0 34176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_352
timestamp 1621261055
transform 1 0 34944 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_356
timestamp 1621261055
transform 1 0 35328 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_359
timestamp 1621261055
transform 1 0 35616 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_367
timestamp 1621261055
transform 1 0 36384 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_375
timestamp 1621261055
transform 1 0 37152 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_383
timestamp 1621261055
transform 1 0 37920 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_391
timestamp 1621261055
transform 1 0 38688 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_643
timestamp 1621261055
transform 1 0 40800 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_399
timestamp 1621261055
transform 1 0 39456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_407
timestamp 1621261055
transform 1 0 40224 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_411
timestamp 1621261055
transform 1 0 40608 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_414
timestamp 1621261055
transform 1 0 40896 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_422
timestamp 1621261055
transform 1 0 41664 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_430
timestamp 1621261055
transform 1 0 42432 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_438
timestamp 1621261055
transform 1 0 43200 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_446
timestamp 1621261055
transform 1 0 43968 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_454
timestamp 1621261055
transform 1 0 44736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_462
timestamp 1621261055
transform 1 0 45504 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_644
timestamp 1621261055
transform 1 0 46080 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_466
timestamp 1621261055
transform 1 0 45888 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_469
timestamp 1621261055
transform 1 0 46176 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_477
timestamp 1621261055
transform 1 0 46944 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_485
timestamp 1621261055
transform 1 0 47712 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_493
timestamp 1621261055
transform 1 0 48480 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_645
timestamp 1621261055
transform 1 0 51360 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_501
timestamp 1621261055
transform 1 0 49248 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_509
timestamp 1621261055
transform 1 0 50016 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_517
timestamp 1621261055
transform 1 0 50784 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_521
timestamp 1621261055
transform 1 0 51168 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_524
timestamp 1621261055
transform 1 0 51456 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_532
timestamp 1621261055
transform 1 0 52224 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_540
timestamp 1621261055
transform 1 0 52992 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_548
timestamp 1621261055
transform 1 0 53760 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_556
timestamp 1621261055
transform 1 0 54528 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_646
timestamp 1621261055
transform 1 0 56640 0 -1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_44_564
timestamp 1621261055
transform 1 0 55296 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_44_572
timestamp 1621261055
transform 1 0 56064 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_576
timestamp 1621261055
transform 1 0 56448 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_44_579
timestamp 1621261055
transform 1 0 56736 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_44_587
timestamp 1621261055
transform 1 0 57504 0 -1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_89
timestamp 1621261055
transform -1 0 58848 0 -1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_44_595
timestamp 1621261055
transform 1 0 58272 0 -1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_90
timestamp 1621261055
transform 1 0 1152 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_4
timestamp 1621261055
transform 1 0 1536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_12
timestamp 1621261055
transform 1 0 2304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_20
timestamp 1621261055
transform 1 0 3072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_28
timestamp 1621261055
transform 1 0 3840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_647
timestamp 1621261055
transform 1 0 6432 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_36
timestamp 1621261055
transform 1 0 4608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_44
timestamp 1621261055
transform 1 0 5376 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_52
timestamp 1621261055
transform 1 0 6144 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_54
timestamp 1621261055
transform 1 0 6336 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_56
timestamp 1621261055
transform 1 0 6528 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_64
timestamp 1621261055
transform 1 0 7296 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_72
timestamp 1621261055
transform 1 0 8064 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_80
timestamp 1621261055
transform 1 0 8832 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_88
timestamp 1621261055
transform 1 0 9600 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_96
timestamp 1621261055
transform 1 0 10368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_648
timestamp 1621261055
transform 1 0 11712 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_104
timestamp 1621261055
transform 1 0 11136 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_108
timestamp 1621261055
transform 1 0 11520 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_111
timestamp 1621261055
transform 1 0 11808 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_119
timestamp 1621261055
transform 1 0 12576 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_127
timestamp 1621261055
transform 1 0 13344 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_649
timestamp 1621261055
transform 1 0 16992 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_135
timestamp 1621261055
transform 1 0 14112 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_143
timestamp 1621261055
transform 1 0 14880 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_151
timestamp 1621261055
transform 1 0 15648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_159
timestamp 1621261055
transform 1 0 16416 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_163
timestamp 1621261055
transform 1 0 16800 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_166
timestamp 1621261055
transform 1 0 17088 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_174
timestamp 1621261055
transform 1 0 17856 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_182
timestamp 1621261055
transform 1 0 18624 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_190
timestamp 1621261055
transform 1 0 19392 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_198
timestamp 1621261055
transform 1 0 20160 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_650
timestamp 1621261055
transform 1 0 22272 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_206
timestamp 1621261055
transform 1 0 20928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_214
timestamp 1621261055
transform 1 0 21696 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_218
timestamp 1621261055
transform 1 0 22080 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_221
timestamp 1621261055
transform 1 0 22368 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_229
timestamp 1621261055
transform 1 0 23136 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_237
timestamp 1621261055
transform 1 0 23904 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_245
timestamp 1621261055
transform 1 0 24672 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_253
timestamp 1621261055
transform 1 0 25440 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_261
timestamp 1621261055
transform 1 0 26208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _076_
timestamp 1621261055
transform -1 0 29664 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_651
timestamp 1621261055
transform 1 0 27552 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_149
timestamp 1621261055
transform -1 0 29376 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_45_269
timestamp 1621261055
transform 1 0 26976 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_273
timestamp 1621261055
transform 1 0 27360 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_276
timestamp 1621261055
transform 1 0 27648 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_284
timestamp 1621261055
transform 1 0 28416 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_297
timestamp 1621261055
transform 1 0 29664 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_652
timestamp 1621261055
transform 1 0 32832 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_305
timestamp 1621261055
transform 1 0 30432 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_313
timestamp 1621261055
transform 1 0 31200 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_321
timestamp 1621261055
transform 1 0 31968 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_45_329
timestamp 1621261055
transform 1 0 32736 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_331
timestamp 1621261055
transform 1 0 32928 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_339
timestamp 1621261055
transform 1 0 33696 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_347
timestamp 1621261055
transform 1 0 34464 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_355
timestamp 1621261055
transform 1 0 35232 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_363
timestamp 1621261055
transform 1 0 36000 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _054_
timestamp 1621261055
transform 1 0 37440 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_653
timestamp 1621261055
transform 1 0 38112 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_371
timestamp 1621261055
transform 1 0 36768 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_375
timestamp 1621261055
transform 1 0 37152 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_45_377
timestamp 1621261055
transform 1 0 37344 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_381
timestamp 1621261055
transform 1 0 37728 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_45_386
timestamp 1621261055
transform 1 0 38208 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_394
timestamp 1621261055
transform 1 0 38976 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_402
timestamp 1621261055
transform 1 0 39744 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_410
timestamp 1621261055
transform 1 0 40512 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_418
timestamp 1621261055
transform 1 0 41280 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_426
timestamp 1621261055
transform 1 0 42048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _049_
timestamp 1621261055
transform 1 0 44736 0 1 32634
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_654
timestamp 1621261055
transform 1 0 43392 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_45_434
timestamp 1621261055
transform 1 0 42816 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_438
timestamp 1621261055
transform 1 0 43200 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_441
timestamp 1621261055
transform 1 0 43488 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_449
timestamp 1621261055
transform 1 0 44256 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_45_453
timestamp 1621261055
transform 1 0 44640 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_457
timestamp 1621261055
transform 1 0 45024 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_655
timestamp 1621261055
transform 1 0 48672 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_465
timestamp 1621261055
transform 1 0 45792 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_473
timestamp 1621261055
transform 1 0 46560 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_481
timestamp 1621261055
transform 1 0 47328 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_489
timestamp 1621261055
transform 1 0 48096 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_493
timestamp 1621261055
transform 1 0 48480 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_496
timestamp 1621261055
transform 1 0 48768 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_504
timestamp 1621261055
transform 1 0 49536 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_512
timestamp 1621261055
transform 1 0 50304 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_520
timestamp 1621261055
transform 1 0 51072 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_528
timestamp 1621261055
transform 1 0 51840 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_656
timestamp 1621261055
transform 1 0 53952 0 1 32634
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_45_536
timestamp 1621261055
transform 1 0 52608 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_544
timestamp 1621261055
transform 1 0 53376 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_548
timestamp 1621261055
transform 1 0 53760 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_45_551
timestamp 1621261055
transform 1 0 54048 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_559
timestamp 1621261055
transform 1 0 54816 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_567
timestamp 1621261055
transform 1 0 55584 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_575
timestamp 1621261055
transform 1 0 56352 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_45_583
timestamp 1621261055
transform 1 0 57120 0 1 32634
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_45_591
timestamp 1621261055
transform 1 0 57888 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_91
timestamp 1621261055
transform -1 0 58848 0 1 32634
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_45_595
timestamp 1621261055
transform 1 0 58272 0 1 32634
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_4
timestamp 1621261055
transform 1 0 1536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_4
timestamp 1621261055
transform 1 0 1536 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_94
timestamp 1621261055
transform 1 0 1152 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_92
timestamp 1621261055
transform 1 0 1152 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_12
timestamp 1621261055
transform 1 0 2304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_12
timestamp 1621261055
transform 1 0 2304 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_20
timestamp 1621261055
transform 1 0 3072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_20
timestamp 1621261055
transform 1 0 3072 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_28
timestamp 1621261055
transform 1 0 3840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_29
timestamp 1621261055
transform 1 0 3936 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_657
timestamp 1621261055
transform 1 0 3840 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_36
timestamp 1621261055
transform 1 0 4608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_37
timestamp 1621261055
transform 1 0 4704 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_44
timestamp 1621261055
transform 1 0 5376 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_45
timestamp 1621261055
transform 1 0 5472 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_56
timestamp 1621261055
transform 1 0 6528 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_54
timestamp 1621261055
transform 1 0 6336 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_52
timestamp 1621261055
transform 1 0 6144 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_53
timestamp 1621261055
transform 1 0 6240 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_668
timestamp 1621261055
transform 1 0 6432 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_64
timestamp 1621261055
transform 1 0 7296 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_61
timestamp 1621261055
transform 1 0 7008 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_72
timestamp 1621261055
transform 1 0 8064 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_69
timestamp 1621261055
transform 1 0 7776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_80
timestamp 1621261055
transform 1 0 8832 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_81
timestamp 1621261055
transform 1 0 8928 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_77
timestamp 1621261055
transform 1 0 8544 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_658
timestamp 1621261055
transform 1 0 9120 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_92
timestamp 1621261055
transform 1 0 9984 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_88
timestamp 1621261055
transform 1 0 9600 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_46_92
timestamp 1621261055
transform 1 0 9984 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_84
timestamp 1621261055
transform 1 0 9216 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _209_
timestamp 1621261055
transform 1 0 9696 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_100
timestamp 1621261055
transform 1 0 10752 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_100
timestamp 1621261055
transform 1 0 10752 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_111
timestamp 1621261055
transform 1 0 11808 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_108
timestamp 1621261055
transform 1 0 11520 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_116
timestamp 1621261055
transform 1 0 12288 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_108
timestamp 1621261055
transform 1 0 11520 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_669
timestamp 1621261055
transform 1 0 11712 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_119
timestamp 1621261055
transform 1 0 12576 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_124
timestamp 1621261055
transform 1 0 13056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_127
timestamp 1621261055
transform 1 0 13344 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_46_132
timestamp 1621261055
transform 1 0 13824 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_101
timestamp 1621261055
transform 1 0 13728 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_47_136
timestamp 1621261055
transform 1 0 14208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_139
timestamp 1621261055
transform 1 0 14496 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_136
timestamp 1621261055
transform 1 0 14208 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_659
timestamp 1621261055
transform 1 0 14400 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _154_
timestamp 1621261055
transform 1 0 13920 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_144
timestamp 1621261055
transform 1 0 14976 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_147
timestamp 1621261055
transform 1 0 15264 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_152
timestamp 1621261055
transform 1 0 15744 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_155
timestamp 1621261055
transform 1 0 16032 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_47_164
timestamp 1621261055
transform 1 0 16896 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_47_160
timestamp 1621261055
transform 1 0 16512 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_163
timestamp 1621261055
transform 1 0 16800 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_670
timestamp 1621261055
transform 1 0 16992 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_170
timestamp 1621261055
transform 1 0 17472 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_166
timestamp 1621261055
transform 1 0 17088 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_171
timestamp 1621261055
transform 1 0 17568 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _090_
timestamp 1621261055
transform 1 0 17664 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_175
timestamp 1621261055
transform 1 0 17952 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_179
timestamp 1621261055
transform 1 0 18336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_191
timestamp 1621261055
transform 1 0 19488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_183
timestamp 1621261055
transform 1 0 18720 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_191
timestamp 1621261055
transform 1 0 19488 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_187
timestamp 1621261055
transform 1 0 19104 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_194
timestamp 1621261055
transform 1 0 19776 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_660
timestamp 1621261055
transform 1 0 19680 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_199
timestamp 1621261055
transform 1 0 20256 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_202
timestamp 1621261055
transform 1 0 20544 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_212
timestamp 1621261055
transform 1 0 21504 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_210
timestamp 1621261055
transform 1 0 21312 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_222
timestamp 1621261055
transform 1 0 21024 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _147_
timestamp 1621261055
transform 1 0 21216 0 1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_221
timestamp 1621261055
transform 1 0 22368 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_218
timestamp 1621261055
transform 1 0 22080 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_671
timestamp 1621261055
transform 1 0 22272 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_229
timestamp 1621261055
transform 1 0 23136 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_226
timestamp 1621261055
transform 1 0 22848 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_237
timestamp 1621261055
transform 1 0 23904 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_234
timestamp 1621261055
transform 1 0 23616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_245
timestamp 1621261055
transform 1 0 24672 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_246
timestamp 1621261055
transform 1 0 24768 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_242
timestamp 1621261055
transform 1 0 24384 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_661
timestamp 1621261055
transform 1 0 24960 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_253
timestamp 1621261055
transform 1 0 25440 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_257
timestamp 1621261055
transform 1 0 25824 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_249
timestamp 1621261055
transform 1 0 25056 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_261
timestamp 1621261055
transform 1 0 26208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_269
timestamp 1621261055
transform 1 0 26976 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_265
timestamp 1621261055
transform 1 0 26592 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_276
timestamp 1621261055
transform 1 0 27648 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_273
timestamp 1621261055
transform 1 0 27360 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_281
timestamp 1621261055
transform 1 0 28128 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_273
timestamp 1621261055
transform 1 0 27360 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_672
timestamp 1621261055
transform 1 0 27552 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_284
timestamp 1621261055
transform 1 0 28416 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_289
timestamp 1621261055
transform 1 0 28896 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_292
timestamp 1621261055
transform 1 0 29184 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_167
timestamp 1621261055
transform -1 0 29472 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _089_
timestamp 1621261055
transform -1 0 29760 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_300
timestamp 1621261055
transform 1 0 29952 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_304
timestamp 1621261055
transform 1 0 30336 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_302
timestamp 1621261055
transform 1 0 30144 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_46_298
timestamp 1621261055
transform 1 0 29760 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_662
timestamp 1621261055
transform 1 0 30240 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_308
timestamp 1621261055
transform 1 0 30720 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_312
timestamp 1621261055
transform 1 0 31104 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_316
timestamp 1621261055
transform 1 0 31488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_320
timestamp 1621261055
transform 1 0 31872 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_328
timestamp 1621261055
transform 1 0 32640 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_324
timestamp 1621261055
transform 1 0 32256 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_328
timestamp 1621261055
transform 1 0 32640 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_673
timestamp 1621261055
transform 1 0 32832 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_331
timestamp 1621261055
transform 1 0 32928 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_336
timestamp 1621261055
transform 1 0 33408 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_347
timestamp 1621261055
transform 1 0 34464 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_339
timestamp 1621261055
transform 1 0 33696 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_346
timestamp 1621261055
transform 1 0 34368 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_344
timestamp 1621261055
transform 1 0 34176 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _190_
timestamp 1621261055
transform 1 0 34464 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_355
timestamp 1621261055
transform 1 0 35232 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_350
timestamp 1621261055
transform 1 0 34752 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_363
timestamp 1621261055
transform 1 0 36000 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_359
timestamp 1621261055
transform 1 0 35616 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_663
timestamp 1621261055
transform 1 0 35520 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_371
timestamp 1621261055
transform 1 0 36768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_367
timestamp 1621261055
transform 1 0 36384 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_379
timestamp 1621261055
transform 1 0 37536 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_379
timestamp 1621261055
transform 1 0 37536 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_375
timestamp 1621261055
transform 1 0 37152 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_386
timestamp 1621261055
transform 1 0 38208 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_383
timestamp 1621261055
transform 1 0 37920 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_387
timestamp 1621261055
transform 1 0 38304 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_381
timestamp 1621261055
transform 1 0 37728 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_206
timestamp 1621261055
transform 1 0 37824 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_674
timestamp 1621261055
transform 1 0 38112 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _136_
timestamp 1621261055
transform 1 0 38016 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_394
timestamp 1621261055
transform 1 0 38976 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_395
timestamp 1621261055
transform 1 0 39072 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_402
timestamp 1621261055
transform 1 0 39744 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_403
timestamp 1621261055
transform 1 0 39840 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_410
timestamp 1621261055
transform 1 0 40512 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_411
timestamp 1621261055
transform 1 0 40608 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_664
timestamp 1621261055
transform 1 0 40800 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_418
timestamp 1621261055
transform 1 0 41280 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_422
timestamp 1621261055
transform 1 0 41664 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_414
timestamp 1621261055
transform 1 0 40896 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_426
timestamp 1621261055
transform 1 0 42048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_46_426
timestamp 1621261055
transform 1 0 42048 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_181
timestamp 1621261055
transform -1 0 42336 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _101_
timestamp 1621261055
transform -1 0 42624 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_47_434
timestamp 1621261055
transform 1 0 42816 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_432
timestamp 1621261055
transform 1 0 42624 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_441
timestamp 1621261055
transform 1 0 43488 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_438
timestamp 1621261055
transform 1 0 43200 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_440
timestamp 1621261055
transform 1 0 43392 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_675
timestamp 1621261055
transform 1 0 43392 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_449
timestamp 1621261055
transform 1 0 44256 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_448
timestamp 1621261055
transform 1 0 44160 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_457
timestamp 1621261055
transform 1 0 45024 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_456
timestamp 1621261055
transform 1 0 44928 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_465
timestamp 1621261055
transform 1 0 45792 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_469
timestamp 1621261055
transform 1 0 46176 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_464
timestamp 1621261055
transform 1 0 45696 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_665
timestamp 1621261055
transform 1 0 46080 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_473
timestamp 1621261055
transform 1 0 46560 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_477
timestamp 1621261055
transform 1 0 46944 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_481
timestamp 1621261055
transform 1 0 47328 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_485
timestamp 1621261055
transform 1 0 47712 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_493
timestamp 1621261055
transform 1 0 48480 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_47_489
timestamp 1621261055
transform 1 0 48096 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_493
timestamp 1621261055
transform 1 0 48480 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_676
timestamp 1621261055
transform 1 0 48672 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_496
timestamp 1621261055
transform 1 0 48768 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_501
timestamp 1621261055
transform 1 0 49248 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_512
timestamp 1621261055
transform 1 0 50304 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_504
timestamp 1621261055
transform 1 0 49536 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_509
timestamp 1621261055
transform 1 0 50016 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_520
timestamp 1621261055
transform 1 0 51072 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_521
timestamp 1621261055
transform 1 0 51168 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_46_517
timestamp 1621261055
transform 1 0 50784 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_47_528
timestamp 1621261055
transform 1 0 51840 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_524
timestamp 1621261055
transform 1 0 51456 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_666
timestamp 1621261055
transform 1 0 51360 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_536
timestamp 1621261055
transform 1 0 52608 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_532
timestamp 1621261055
transform 1 0 52224 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_544
timestamp 1621261055
transform 1 0 53376 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_46_540
timestamp 1621261055
transform 1 0 52992 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_551
timestamp 1621261055
transform 1 0 54048 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_548
timestamp 1621261055
transform 1 0 53760 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_46_548
timestamp 1621261055
transform 1 0 53760 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_677
timestamp 1621261055
transform 1 0 53952 0 1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_47_559
timestamp 1621261055
transform 1 0 54816 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_556
timestamp 1621261055
transform 1 0 54528 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_47_567
timestamp 1621261055
transform 1 0 55584 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_567
timestamp 1621261055
transform 1 0 55584 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _112_
timestamp 1621261055
transform 1 0 55296 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_575
timestamp 1621261055
transform 1 0 56352 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_46_574
timestamp 1621261055
transform 1 0 56256 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_667
timestamp 1621261055
transform 1 0 56640 0 -1 33966
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _030_
timestamp 1621261055
transform 1 0 55968 0 -1 33966
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_47_583
timestamp 1621261055
transform 1 0 57120 0 1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_587
timestamp 1621261055
transform 1 0 57504 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_46_579
timestamp 1621261055
transform 1 0 56736 0 -1 33966
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_47_591
timestamp 1621261055
transform 1 0 57888 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_93
timestamp 1621261055
transform -1 0 58848 0 -1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_95
timestamp 1621261055
transform -1 0 58848 0 1 33966
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_46_595
timestamp 1621261055
transform 1 0 58272 0 -1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_47_595
timestamp 1621261055
transform 1 0 58272 0 1 33966
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_96
timestamp 1621261055
transform 1 0 1152 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_678
timestamp 1621261055
transform 1 0 3840 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_4
timestamp 1621261055
transform 1 0 1536 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_12
timestamp 1621261055
transform 1 0 2304 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_20
timestamp 1621261055
transform 1 0 3072 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_29
timestamp 1621261055
transform 1 0 3936 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_37
timestamp 1621261055
transform 1 0 4704 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_45
timestamp 1621261055
transform 1 0 5472 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_53
timestamp 1621261055
transform 1 0 6240 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_61
timestamp 1621261055
transform 1 0 7008 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_679
timestamp 1621261055
transform 1 0 9120 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_69
timestamp 1621261055
transform 1 0 7776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_77
timestamp 1621261055
transform 1 0 8544 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_81
timestamp 1621261055
transform 1 0 8928 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_84
timestamp 1621261055
transform 1 0 9216 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_92
timestamp 1621261055
transform 1 0 9984 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _109_
timestamp 1621261055
transform 1 0 12672 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_185
timestamp 1621261055
transform 1 0 12480 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_100
timestamp 1621261055
transform 1 0 10752 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_108
timestamp 1621261055
transform 1 0 11520 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_116
timestamp 1621261055
transform 1 0 12288 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_123
timestamp 1621261055
transform 1 0 12960 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_131
timestamp 1621261055
transform 1 0 13728 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_680
timestamp 1621261055
transform 1 0 14400 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_135
timestamp 1621261055
transform 1 0 14112 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_137
timestamp 1621261055
transform 1 0 14304 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_139
timestamp 1621261055
transform 1 0 14496 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_147
timestamp 1621261055
transform 1 0 15264 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_155
timestamp 1621261055
transform 1 0 16032 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_163
timestamp 1621261055
transform 1 0 16800 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_681
timestamp 1621261055
transform 1 0 19680 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_171
timestamp 1621261055
transform 1 0 17568 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_179
timestamp 1621261055
transform 1 0 18336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_187
timestamp 1621261055
transform 1 0 19104 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_191
timestamp 1621261055
transform 1 0 19488 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_194
timestamp 1621261055
transform 1 0 19776 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_202
timestamp 1621261055
transform 1 0 20544 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_210
timestamp 1621261055
transform 1 0 21312 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_218
timestamp 1621261055
transform 1 0 22080 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_226
timestamp 1621261055
transform 1 0 22848 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_682
timestamp 1621261055
transform 1 0 24960 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_234
timestamp 1621261055
transform 1 0 23616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_242
timestamp 1621261055
transform 1 0 24384 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_246
timestamp 1621261055
transform 1 0 24768 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_249
timestamp 1621261055
transform 1 0 25056 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_257
timestamp 1621261055
transform 1 0 25824 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_265
timestamp 1621261055
transform 1 0 26592 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_273
timestamp 1621261055
transform 1 0 27360 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_281
timestamp 1621261055
transform 1 0 28128 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_289
timestamp 1621261055
transform 1 0 28896 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_297
timestamp 1621261055
transform 1 0 29664 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_683
timestamp 1621261055
transform 1 0 30240 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_301
timestamp 1621261055
transform 1 0 30048 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_304
timestamp 1621261055
transform 1 0 30336 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_312
timestamp 1621261055
transform 1 0 31104 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_320
timestamp 1621261055
transform 1 0 31872 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_328
timestamp 1621261055
transform 1 0 32640 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_684
timestamp 1621261055
transform 1 0 35520 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_336
timestamp 1621261055
transform 1 0 33408 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_344
timestamp 1621261055
transform 1 0 34176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_352
timestamp 1621261055
transform 1 0 34944 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_356
timestamp 1621261055
transform 1 0 35328 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_359
timestamp 1621261055
transform 1 0 35616 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_367
timestamp 1621261055
transform 1 0 36384 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_375
timestamp 1621261055
transform 1 0 37152 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_383
timestamp 1621261055
transform 1 0 37920 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_391
timestamp 1621261055
transform 1 0 38688 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _207_
timestamp 1621261055
transform -1 0 41952 0 -1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_685
timestamp 1621261055
transform 1 0 40800 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_248
timestamp 1621261055
transform -1 0 41664 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_399
timestamp 1621261055
transform 1 0 39456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_407
timestamp 1621261055
transform 1 0 40224 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_411
timestamp 1621261055
transform 1 0 40608 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_48_414
timestamp 1621261055
transform 1 0 40896 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_418
timestamp 1621261055
transform 1 0 41280 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_425
timestamp 1621261055
transform 1 0 41952 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_433
timestamp 1621261055
transform 1 0 42720 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_441
timestamp 1621261055
transform 1 0 43488 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_449
timestamp 1621261055
transform 1 0 44256 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_457
timestamp 1621261055
transform 1 0 45024 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_686
timestamp 1621261055
transform 1 0 46080 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_465
timestamp 1621261055
transform 1 0 45792 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_48_467
timestamp 1621261055
transform 1 0 45984 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_469
timestamp 1621261055
transform 1 0 46176 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_477
timestamp 1621261055
transform 1 0 46944 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_485
timestamp 1621261055
transform 1 0 47712 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_493
timestamp 1621261055
transform 1 0 48480 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_687
timestamp 1621261055
transform 1 0 51360 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_501
timestamp 1621261055
transform 1 0 49248 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_509
timestamp 1621261055
transform 1 0 50016 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_517
timestamp 1621261055
transform 1 0 50784 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_521
timestamp 1621261055
transform 1 0 51168 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_524
timestamp 1621261055
transform 1 0 51456 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_532
timestamp 1621261055
transform 1 0 52224 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_540
timestamp 1621261055
transform 1 0 52992 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_548
timestamp 1621261055
transform 1 0 53760 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_556
timestamp 1621261055
transform 1 0 54528 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_688
timestamp 1621261055
transform 1 0 56640 0 -1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_48_564
timestamp 1621261055
transform 1 0 55296 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_48_572
timestamp 1621261055
transform 1 0 56064 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_576
timestamp 1621261055
transform 1 0 56448 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_48_579
timestamp 1621261055
transform 1 0 56736 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_48_587
timestamp 1621261055
transform 1 0 57504 0 -1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_97
timestamp 1621261055
transform -1 0 58848 0 -1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_48_595
timestamp 1621261055
transform 1 0 58272 0 -1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_98
timestamp 1621261055
transform 1 0 1152 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_49_4
timestamp 1621261055
transform 1 0 1536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_12
timestamp 1621261055
transform 1 0 2304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_20
timestamp 1621261055
transform 1 0 3072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_28
timestamp 1621261055
transform 1 0 3840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_689
timestamp 1621261055
transform 1 0 6432 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_36
timestamp 1621261055
transform 1 0 4608 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_44
timestamp 1621261055
transform 1 0 5376 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_52
timestamp 1621261055
transform 1 0 6144 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_49_54
timestamp 1621261055
transform 1 0 6336 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_56
timestamp 1621261055
transform 1 0 6528 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_64
timestamp 1621261055
transform 1 0 7296 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_72
timestamp 1621261055
transform 1 0 8064 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_80
timestamp 1621261055
transform 1 0 8832 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_88
timestamp 1621261055
transform 1 0 9600 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_96
timestamp 1621261055
transform 1 0 10368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_690
timestamp 1621261055
transform 1 0 11712 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_104
timestamp 1621261055
transform 1 0 11136 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_108
timestamp 1621261055
transform 1 0 11520 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_111
timestamp 1621261055
transform 1 0 11808 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_119
timestamp 1621261055
transform 1 0 12576 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_127
timestamp 1621261055
transform 1 0 13344 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_691
timestamp 1621261055
transform 1 0 16992 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_135
timestamp 1621261055
transform 1 0 14112 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_143
timestamp 1621261055
transform 1 0 14880 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_151
timestamp 1621261055
transform 1 0 15648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_159
timestamp 1621261055
transform 1 0 16416 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_163
timestamp 1621261055
transform 1 0 16800 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_166
timestamp 1621261055
transform 1 0 17088 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_174
timestamp 1621261055
transform 1 0 17856 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_182
timestamp 1621261055
transform 1 0 18624 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_190
timestamp 1621261055
transform 1 0 19392 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_198
timestamp 1621261055
transform 1 0 20160 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_692
timestamp 1621261055
transform 1 0 22272 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_206
timestamp 1621261055
transform 1 0 20928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_214
timestamp 1621261055
transform 1 0 21696 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_218
timestamp 1621261055
transform 1 0 22080 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_221
timestamp 1621261055
transform 1 0 22368 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_229
timestamp 1621261055
transform 1 0 23136 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_237
timestamp 1621261055
transform 1 0 23904 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_245
timestamp 1621261055
transform 1 0 24672 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_253
timestamp 1621261055
transform 1 0 25440 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_261
timestamp 1621261055
transform 1 0 26208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_693
timestamp 1621261055
transform 1 0 27552 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_49_269
timestamp 1621261055
transform 1 0 26976 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_273
timestamp 1621261055
transform 1 0 27360 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_276
timestamp 1621261055
transform 1 0 27648 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_284
timestamp 1621261055
transform 1 0 28416 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_292
timestamp 1621261055
transform 1 0 29184 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_694
timestamp 1621261055
transform 1 0 32832 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_300
timestamp 1621261055
transform 1 0 29952 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_308
timestamp 1621261055
transform 1 0 30720 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_316
timestamp 1621261055
transform 1 0 31488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_324
timestamp 1621261055
transform 1 0 32256 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_328
timestamp 1621261055
transform 1 0 32640 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_331
timestamp 1621261055
transform 1 0 32928 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_339
timestamp 1621261055
transform 1 0 33696 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_347
timestamp 1621261055
transform 1 0 34464 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_355
timestamp 1621261055
transform 1 0 35232 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_363
timestamp 1621261055
transform 1 0 36000 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_695
timestamp 1621261055
transform 1 0 38112 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_371
timestamp 1621261055
transform 1 0 36768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_379
timestamp 1621261055
transform 1 0 37536 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_383
timestamp 1621261055
transform 1 0 37920 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_386
timestamp 1621261055
transform 1 0 38208 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_394
timestamp 1621261055
transform 1 0 38976 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _013_
timestamp 1621261055
transform 1 0 41472 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_49_402
timestamp 1621261055
transform 1 0 39744 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_410
timestamp 1621261055
transform 1 0 40512 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_418
timestamp 1621261055
transform 1 0 41280 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_423
timestamp 1621261055
transform 1 0 41760 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_696
timestamp 1621261055
transform 1 0 43392 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_431
timestamp 1621261055
transform 1 0 42528 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_49_439
timestamp 1621261055
transform 1 0 43296 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_441
timestamp 1621261055
transform 1 0 43488 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_449
timestamp 1621261055
transform 1 0 44256 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_457
timestamp 1621261055
transform 1 0 45024 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _150_
timestamp 1621261055
transform 1 0 46464 0 1 35298
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_697
timestamp 1621261055
transform 1 0 48672 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_225
timestamp 1621261055
transform 1 0 46272 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_49_465
timestamp 1621261055
transform 1 0 45792 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_49_469
timestamp 1621261055
transform 1 0 46176 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_475
timestamp 1621261055
transform 1 0 46752 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_483
timestamp 1621261055
transform 1 0 47520 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_491
timestamp 1621261055
transform 1 0 48288 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_49_496
timestamp 1621261055
transform 1 0 48768 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_504
timestamp 1621261055
transform 1 0 49536 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_512
timestamp 1621261055
transform 1 0 50304 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_520
timestamp 1621261055
transform 1 0 51072 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_528
timestamp 1621261055
transform 1 0 51840 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_698
timestamp 1621261055
transform 1 0 53952 0 1 35298
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_49_536
timestamp 1621261055
transform 1 0 52608 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_544
timestamp 1621261055
transform 1 0 53376 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_548
timestamp 1621261055
transform 1 0 53760 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_49_551
timestamp 1621261055
transform 1 0 54048 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_559
timestamp 1621261055
transform 1 0 54816 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_567
timestamp 1621261055
transform 1 0 55584 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_575
timestamp 1621261055
transform 1 0 56352 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_49_583
timestamp 1621261055
transform 1 0 57120 0 1 35298
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_49_591
timestamp 1621261055
transform 1 0 57888 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_99
timestamp 1621261055
transform -1 0 58848 0 1 35298
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_49_595
timestamp 1621261055
transform 1 0 58272 0 1 35298
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_100
timestamp 1621261055
transform 1 0 1152 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_699
timestamp 1621261055
transform 1 0 3840 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_4
timestamp 1621261055
transform 1 0 1536 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_12
timestamp 1621261055
transform 1 0 2304 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_20
timestamp 1621261055
transform 1 0 3072 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_29
timestamp 1621261055
transform 1 0 3936 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_37
timestamp 1621261055
transform 1 0 4704 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_45
timestamp 1621261055
transform 1 0 5472 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_53
timestamp 1621261055
transform 1 0 6240 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_61
timestamp 1621261055
transform 1 0 7008 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_700
timestamp 1621261055
transform 1 0 9120 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_69
timestamp 1621261055
transform 1 0 7776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_77
timestamp 1621261055
transform 1 0 8544 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_81
timestamp 1621261055
transform 1 0 8928 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_84
timestamp 1621261055
transform 1 0 9216 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_92
timestamp 1621261055
transform 1 0 9984 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_100
timestamp 1621261055
transform 1 0 10752 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_108
timestamp 1621261055
transform 1 0 11520 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_116
timestamp 1621261055
transform 1 0 12288 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_124
timestamp 1621261055
transform 1 0 13056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_132
timestamp 1621261055
transform 1 0 13824 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_701
timestamp 1621261055
transform 1 0 14400 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_136
timestamp 1621261055
transform 1 0 14208 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_139
timestamp 1621261055
transform 1 0 14496 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_147
timestamp 1621261055
transform 1 0 15264 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_155
timestamp 1621261055
transform 1 0 16032 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_163
timestamp 1621261055
transform 1 0 16800 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_702
timestamp 1621261055
transform 1 0 19680 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_171
timestamp 1621261055
transform 1 0 17568 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_179
timestamp 1621261055
transform 1 0 18336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_187
timestamp 1621261055
transform 1 0 19104 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_191
timestamp 1621261055
transform 1 0 19488 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_194
timestamp 1621261055
transform 1 0 19776 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _017_
timestamp 1621261055
transform 1 0 21984 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _080_
timestamp 1621261055
transform 1 0 21312 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_153
timestamp 1621261055
transform 1 0 21120 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_202
timestamp 1621261055
transform 1 0 20544 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_206
timestamp 1621261055
transform 1 0 20928 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_50_213
timestamp 1621261055
transform 1 0 21600 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_220
timestamp 1621261055
transform 1 0 22272 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_228
timestamp 1621261055
transform 1 0 23040 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _141_
timestamp 1621261055
transform 1 0 25632 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_703
timestamp 1621261055
transform 1 0 24960 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_211
timestamp 1621261055
transform 1 0 25440 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_236
timestamp 1621261055
transform 1 0 23808 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_244
timestamp 1621261055
transform 1 0 24576 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_50_249
timestamp 1621261055
transform 1 0 25056 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_50_258
timestamp 1621261055
transform 1 0 25920 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_266
timestamp 1621261055
transform 1 0 26688 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_274
timestamp 1621261055
transform 1 0 27456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_282
timestamp 1621261055
transform 1 0 28224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_290
timestamp 1621261055
transform 1 0 28992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_704
timestamp 1621261055
transform 1 0 30240 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_50_298
timestamp 1621261055
transform 1 0 29760 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_50_302
timestamp 1621261055
transform 1 0 30144 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_304
timestamp 1621261055
transform 1 0 30336 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_312
timestamp 1621261055
transform 1 0 31104 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_320
timestamp 1621261055
transform 1 0 31872 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_328
timestamp 1621261055
transform 1 0 32640 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _059_
timestamp 1621261055
transform -1 0 33888 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_705
timestamp 1621261055
transform 1 0 35520 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_97
timestamp 1621261055
transform -1 0 33600 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_341
timestamp 1621261055
transform 1 0 33888 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_349
timestamp 1621261055
transform 1 0 34656 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_50_357
timestamp 1621261055
transform 1 0 35424 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_359
timestamp 1621261055
transform 1 0 35616 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _155_
timestamp 1621261055
transform 1 0 36768 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_104
timestamp 1621261055
transform 1 0 36576 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_367
timestamp 1621261055
transform 1 0 36384 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_374
timestamp 1621261055
transform 1 0 37056 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_382
timestamp 1621261055
transform 1 0 37824 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_390
timestamp 1621261055
transform 1 0 38592 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_706
timestamp 1621261055
transform 1 0 40800 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_398
timestamp 1621261055
transform 1 0 39360 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_406
timestamp 1621261055
transform 1 0 40128 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_410
timestamp 1621261055
transform 1 0 40512 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_412
timestamp 1621261055
transform 1 0 40704 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_414
timestamp 1621261055
transform 1 0 40896 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_422
timestamp 1621261055
transform 1 0 41664 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_430
timestamp 1621261055
transform 1 0 42432 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_438
timestamp 1621261055
transform 1 0 43200 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_446
timestamp 1621261055
transform 1 0 43968 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_454
timestamp 1621261055
transform 1 0 44736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_462
timestamp 1621261055
transform 1 0 45504 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_707
timestamp 1621261055
transform 1 0 46080 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_466
timestamp 1621261055
transform 1 0 45888 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_469
timestamp 1621261055
transform 1 0 46176 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_477
timestamp 1621261055
transform 1 0 46944 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_485
timestamp 1621261055
transform 1 0 47712 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_493
timestamp 1621261055
transform 1 0 48480 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _099_
timestamp 1621261055
transform 1 0 50400 0 -1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_708
timestamp 1621261055
transform 1 0 51360 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_501
timestamp 1621261055
transform 1 0 49248 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_509
timestamp 1621261055
transform 1 0 50016 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_50_516
timestamp 1621261055
transform 1 0 50688 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_520
timestamp 1621261055
transform 1 0 51072 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_50_522
timestamp 1621261055
transform 1 0 51264 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_524
timestamp 1621261055
transform 1 0 51456 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_532
timestamp 1621261055
transform 1 0 52224 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_540
timestamp 1621261055
transform 1 0 52992 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_548
timestamp 1621261055
transform 1 0 53760 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_556
timestamp 1621261055
transform 1 0 54528 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_709
timestamp 1621261055
transform 1 0 56640 0 -1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_50_564
timestamp 1621261055
transform 1 0 55296 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_50_572
timestamp 1621261055
transform 1 0 56064 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_576
timestamp 1621261055
transform 1 0 56448 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_50_579
timestamp 1621261055
transform 1 0 56736 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_50_587
timestamp 1621261055
transform 1 0 57504 0 -1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_101
timestamp 1621261055
transform -1 0 58848 0 -1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_50_595
timestamp 1621261055
transform 1 0 58272 0 -1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_102
timestamp 1621261055
transform 1 0 1152 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_4
timestamp 1621261055
transform 1 0 1536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_12
timestamp 1621261055
transform 1 0 2304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_20
timestamp 1621261055
transform 1 0 3072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_28
timestamp 1621261055
transform 1 0 3840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _016_
timestamp 1621261055
transform 1 0 6912 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_710
timestamp 1621261055
transform 1 0 6432 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_36
timestamp 1621261055
transform 1 0 4608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_44
timestamp 1621261055
transform 1 0 5376 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_52
timestamp 1621261055
transform 1 0 6144 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_54
timestamp 1621261055
transform 1 0 6336 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_56
timestamp 1621261055
transform 1 0 6528 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_63
timestamp 1621261055
transform 1 0 7200 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_71
timestamp 1621261055
transform 1 0 7968 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_79
timestamp 1621261055
transform 1 0 8736 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_87
timestamp 1621261055
transform 1 0 9504 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_95
timestamp 1621261055
transform 1 0 10272 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_711
timestamp 1621261055
transform 1 0 11712 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_103
timestamp 1621261055
transform 1 0 11040 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_107
timestamp 1621261055
transform 1 0 11424 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_109
timestamp 1621261055
transform 1 0 11616 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_111
timestamp 1621261055
transform 1 0 11808 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_119
timestamp 1621261055
transform 1 0 12576 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_127
timestamp 1621261055
transform 1 0 13344 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_712
timestamp 1621261055
transform 1 0 16992 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_135
timestamp 1621261055
transform 1 0 14112 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_143
timestamp 1621261055
transform 1 0 14880 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_151
timestamp 1621261055
transform 1 0 15648 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_159
timestamp 1621261055
transform 1 0 16416 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_163
timestamp 1621261055
transform 1 0 16800 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_166
timestamp 1621261055
transform 1 0 17088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_174
timestamp 1621261055
transform 1 0 17856 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_182
timestamp 1621261055
transform 1 0 18624 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_190
timestamp 1621261055
transform 1 0 19392 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_198
timestamp 1621261055
transform 1 0 20160 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_713
timestamp 1621261055
transform 1 0 22272 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_206
timestamp 1621261055
transform 1 0 20928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_214
timestamp 1621261055
transform 1 0 21696 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_218
timestamp 1621261055
transform 1 0 22080 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_221
timestamp 1621261055
transform 1 0 22368 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_229
timestamp 1621261055
transform 1 0 23136 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _010_
timestamp 1621261055
transform 1 0 24096 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _055_
timestamp 1621261055
transform 1 0 24768 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_237
timestamp 1621261055
transform 1 0 23904 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_51_242
timestamp 1621261055
transform 1 0 24384 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_51_249
timestamp 1621261055
transform 1 0 25056 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_257
timestamp 1621261055
transform 1 0 25824 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _144_
timestamp 1621261055
transform 1 0 28032 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_714
timestamp 1621261055
transform 1 0 27552 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_217
timestamp 1621261055
transform 1 0 27840 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_265
timestamp 1621261055
transform 1 0 26592 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_273
timestamp 1621261055
transform 1 0 27360 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_276
timestamp 1621261055
transform 1 0 27648 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_283
timestamp 1621261055
transform 1 0 28320 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_291
timestamp 1621261055
transform 1 0 29088 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_715
timestamp 1621261055
transform 1 0 32832 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_299
timestamp 1621261055
transform 1 0 29856 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_307
timestamp 1621261055
transform 1 0 30624 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_315
timestamp 1621261055
transform 1 0 31392 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_323
timestamp 1621261055
transform 1 0 32160 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_327
timestamp 1621261055
transform 1 0 32544 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_51_329
timestamp 1621261055
transform 1 0 32736 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_331
timestamp 1621261055
transform 1 0 32928 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_339
timestamp 1621261055
transform 1 0 33696 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_347
timestamp 1621261055
transform 1 0 34464 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_355
timestamp 1621261055
transform 1 0 35232 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_363
timestamp 1621261055
transform 1 0 36000 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_716
timestamp 1621261055
transform 1 0 38112 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_371
timestamp 1621261055
transform 1 0 36768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_379
timestamp 1621261055
transform 1 0 37536 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_383
timestamp 1621261055
transform 1 0 37920 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_386
timestamp 1621261055
transform 1 0 38208 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_394
timestamp 1621261055
transform 1 0 38976 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_402
timestamp 1621261055
transform 1 0 39744 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_410
timestamp 1621261055
transform 1 0 40512 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_418
timestamp 1621261055
transform 1 0 41280 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_426
timestamp 1621261055
transform 1 0 42048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_717
timestamp 1621261055
transform 1 0 43392 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_51_434
timestamp 1621261055
transform 1 0 42816 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_438
timestamp 1621261055
transform 1 0 43200 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_441
timestamp 1621261055
transform 1 0 43488 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_449
timestamp 1621261055
transform 1 0 44256 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_457
timestamp 1621261055
transform 1 0 45024 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_718
timestamp 1621261055
transform 1 0 48672 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_465
timestamp 1621261055
transform 1 0 45792 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_473
timestamp 1621261055
transform 1 0 46560 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_481
timestamp 1621261055
transform 1 0 47328 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_489
timestamp 1621261055
transform 1 0 48096 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_493
timestamp 1621261055
transform 1 0 48480 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_496
timestamp 1621261055
transform 1 0 48768 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_504
timestamp 1621261055
transform 1 0 49536 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_512
timestamp 1621261055
transform 1 0 50304 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_520
timestamp 1621261055
transform 1 0 51072 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_528
timestamp 1621261055
transform 1 0 51840 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_719
timestamp 1621261055
transform 1 0 53952 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_51_536
timestamp 1621261055
transform 1 0 52608 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_544
timestamp 1621261055
transform 1 0 53376 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_548
timestamp 1621261055
transform 1 0 53760 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_551
timestamp 1621261055
transform 1 0 54048 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_559
timestamp 1621261055
transform 1 0 54816 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _078_
timestamp 1621261055
transform 1 0 56160 0 1 36630
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_51_567
timestamp 1621261055
transform 1 0 55584 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_51_571
timestamp 1621261055
transform 1 0 55968 0 1 36630
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_51_576
timestamp 1621261055
transform 1 0 56448 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_51_584
timestamp 1621261055
transform 1 0 57216 0 1 36630
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_51_592
timestamp 1621261055
transform 1 0 57984 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_103
timestamp 1621261055
transform -1 0 58848 0 1 36630
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_51_596
timestamp 1621261055
transform 1 0 58368 0 1 36630
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _183_
timestamp 1621261055
transform 1 0 1632 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_104
timestamp 1621261055
transform 1 0 1152 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_720
timestamp 1621261055
transform 1 0 3840 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_240
timestamp 1621261055
transform 1 0 1920 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_4
timestamp 1621261055
transform 1 0 1536 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_10
timestamp 1621261055
transform 1 0 2112 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_18
timestamp 1621261055
transform 1 0 2880 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_26
timestamp 1621261055
transform 1 0 3648 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_29
timestamp 1621261055
transform 1 0 3936 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _215_
timestamp 1621261055
transform 1 0 5280 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_52_37
timestamp 1621261055
transform 1 0 4704 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_41
timestamp 1621261055
transform 1 0 5088 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_46
timestamp 1621261055
transform 1 0 5568 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_54
timestamp 1621261055
transform 1 0 6336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_62
timestamp 1621261055
transform 1 0 7104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_721
timestamp 1621261055
transform 1 0 9120 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_70
timestamp 1621261055
transform 1 0 7872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_78
timestamp 1621261055
transform 1 0 8640 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_52_82
timestamp 1621261055
transform 1 0 9024 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_84
timestamp 1621261055
transform 1 0 9216 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_92
timestamp 1621261055
transform 1 0 9984 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_100
timestamp 1621261055
transform 1 0 10752 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_108
timestamp 1621261055
transform 1 0 11520 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_116
timestamp 1621261055
transform 1 0 12288 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_124
timestamp 1621261055
transform 1 0 13056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_132
timestamp 1621261055
transform 1 0 13824 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_722
timestamp 1621261055
transform 1 0 14400 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_136
timestamp 1621261055
transform 1 0 14208 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_139
timestamp 1621261055
transform 1 0 14496 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_147
timestamp 1621261055
transform 1 0 15264 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_155
timestamp 1621261055
transform 1 0 16032 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_163
timestamp 1621261055
transform 1 0 16800 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_723
timestamp 1621261055
transform 1 0 19680 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_171
timestamp 1621261055
transform 1 0 17568 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_179
timestamp 1621261055
transform 1 0 18336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_187
timestamp 1621261055
transform 1 0 19104 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_191
timestamp 1621261055
transform 1 0 19488 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_194
timestamp 1621261055
transform 1 0 19776 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_202
timestamp 1621261055
transform 1 0 20544 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_210
timestamp 1621261055
transform 1 0 21312 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_218
timestamp 1621261055
transform 1 0 22080 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_226
timestamp 1621261055
transform 1 0 22848 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_724
timestamp 1621261055
transform 1 0 24960 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_234
timestamp 1621261055
transform 1 0 23616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_242
timestamp 1621261055
transform 1 0 24384 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_246
timestamp 1621261055
transform 1 0 24768 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_249
timestamp 1621261055
transform 1 0 25056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_257
timestamp 1621261055
transform 1 0 25824 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_265
timestamp 1621261055
transform 1 0 26592 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_273
timestamp 1621261055
transform 1 0 27360 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_281
timestamp 1621261055
transform 1 0 28128 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_289
timestamp 1621261055
transform 1 0 28896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_297
timestamp 1621261055
transform 1 0 29664 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_725
timestamp 1621261055
transform 1 0 30240 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_301
timestamp 1621261055
transform 1 0 30048 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_304
timestamp 1621261055
transform 1 0 30336 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_312
timestamp 1621261055
transform 1 0 31104 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_320
timestamp 1621261055
transform 1 0 31872 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_328
timestamp 1621261055
transform 1 0 32640 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_726
timestamp 1621261055
transform 1 0 35520 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_336
timestamp 1621261055
transform 1 0 33408 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_344
timestamp 1621261055
transform 1 0 34176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_352
timestamp 1621261055
transform 1 0 34944 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_356
timestamp 1621261055
transform 1 0 35328 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_359
timestamp 1621261055
transform 1 0 35616 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_367
timestamp 1621261055
transform 1 0 36384 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_375
timestamp 1621261055
transform 1 0 37152 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_383
timestamp 1621261055
transform 1 0 37920 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_391
timestamp 1621261055
transform 1 0 38688 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_727
timestamp 1621261055
transform 1 0 40800 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_399
timestamp 1621261055
transform 1 0 39456 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_407
timestamp 1621261055
transform 1 0 40224 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_411
timestamp 1621261055
transform 1 0 40608 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_414
timestamp 1621261055
transform 1 0 40896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_422
timestamp 1621261055
transform 1 0 41664 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_430
timestamp 1621261055
transform 1 0 42432 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_438
timestamp 1621261055
transform 1 0 43200 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_446
timestamp 1621261055
transform 1 0 43968 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_454
timestamp 1621261055
transform 1 0 44736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_462
timestamp 1621261055
transform 1 0 45504 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _145_
timestamp 1621261055
transform 1 0 47232 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_728
timestamp 1621261055
transform 1 0 46080 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_466
timestamp 1621261055
transform 1 0 45888 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_469
timestamp 1621261055
transform 1 0 46176 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_477
timestamp 1621261055
transform 1 0 46944 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_479
timestamp 1621261055
transform 1 0 47136 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_483
timestamp 1621261055
transform 1 0 47520 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_491
timestamp 1621261055
transform 1 0 48288 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _200_
timestamp 1621261055
transform -1 0 52128 0 -1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_729
timestamp 1621261055
transform 1 0 51360 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_236
timestamp 1621261055
transform -1 0 51840 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_499
timestamp 1621261055
transform 1 0 49056 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_507
timestamp 1621261055
transform 1 0 49824 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_515
timestamp 1621261055
transform 1 0 50592 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_524
timestamp 1621261055
transform 1 0 51456 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_52_531
timestamp 1621261055
transform 1 0 52128 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_539
timestamp 1621261055
transform 1 0 52896 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_547
timestamp 1621261055
transform 1 0 53664 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_555
timestamp 1621261055
transform 1 0 54432 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_730
timestamp 1621261055
transform 1 0 56640 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_563
timestamp 1621261055
transform 1 0 55200 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_52_571
timestamp 1621261055
transform 1 0 55968 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_575
timestamp 1621261055
transform 1 0 56352 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_52_577
timestamp 1621261055
transform 1 0 56544 0 -1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_52_579
timestamp 1621261055
transform 1 0 56736 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_52_587
timestamp 1621261055
transform 1 0 57504 0 -1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_105
timestamp 1621261055
transform -1 0 58848 0 -1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_52_595
timestamp 1621261055
transform 1 0 58272 0 -1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_106
timestamp 1621261055
transform 1 0 1152 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_4
timestamp 1621261055
transform 1 0 1536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_12
timestamp 1621261055
transform 1 0 2304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_20
timestamp 1621261055
transform 1 0 3072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_28
timestamp 1621261055
transform 1 0 3840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_731
timestamp 1621261055
transform 1 0 6432 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_36
timestamp 1621261055
transform 1 0 4608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_44
timestamp 1621261055
transform 1 0 5376 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_52
timestamp 1621261055
transform 1 0 6144 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_54
timestamp 1621261055
transform 1 0 6336 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_56
timestamp 1621261055
transform 1 0 6528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_64
timestamp 1621261055
transform 1 0 7296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_72
timestamp 1621261055
transform 1 0 8064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_80
timestamp 1621261055
transform 1 0 8832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_88
timestamp 1621261055
transform 1 0 9600 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_96
timestamp 1621261055
transform 1 0 10368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_732
timestamp 1621261055
transform 1 0 11712 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_104
timestamp 1621261055
transform 1 0 11136 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_108
timestamp 1621261055
transform 1 0 11520 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_111
timestamp 1621261055
transform 1 0 11808 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_119
timestamp 1621261055
transform 1 0 12576 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_127
timestamp 1621261055
transform 1 0 13344 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_733
timestamp 1621261055
transform 1 0 16992 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_135
timestamp 1621261055
transform 1 0 14112 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_143
timestamp 1621261055
transform 1 0 14880 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_151
timestamp 1621261055
transform 1 0 15648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_159
timestamp 1621261055
transform 1 0 16416 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_163
timestamp 1621261055
transform 1 0 16800 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _037_
timestamp 1621261055
transform 1 0 17472 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_53_166
timestamp 1621261055
transform 1 0 17088 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_173
timestamp 1621261055
transform 1 0 17760 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_181
timestamp 1621261055
transform 1 0 18528 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_189
timestamp 1621261055
transform 1 0 19296 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_197
timestamp 1621261055
transform 1 0 20064 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_734
timestamp 1621261055
transform 1 0 22272 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_205
timestamp 1621261055
transform 1 0 20832 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_213
timestamp 1621261055
transform 1 0 21600 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_217
timestamp 1621261055
transform 1 0 21984 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_219
timestamp 1621261055
transform 1 0 22176 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_221
timestamp 1621261055
transform 1 0 22368 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_229
timestamp 1621261055
transform 1 0 23136 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_237
timestamp 1621261055
transform 1 0 23904 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_245
timestamp 1621261055
transform 1 0 24672 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_253
timestamp 1621261055
transform 1 0 25440 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_261
timestamp 1621261055
transform 1 0 26208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_735
timestamp 1621261055
transform 1 0 27552 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_269
timestamp 1621261055
transform 1 0 26976 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_273
timestamp 1621261055
transform 1 0 27360 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_276
timestamp 1621261055
transform 1 0 27648 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_284
timestamp 1621261055
transform 1 0 28416 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_292
timestamp 1621261055
transform 1 0 29184 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_736
timestamp 1621261055
transform 1 0 32832 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_300
timestamp 1621261055
transform 1 0 29952 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_308
timestamp 1621261055
transform 1 0 30720 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_316
timestamp 1621261055
transform 1 0 31488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_324
timestamp 1621261055
transform 1 0 32256 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_328
timestamp 1621261055
transform 1 0 32640 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_331
timestamp 1621261055
transform 1 0 32928 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_339
timestamp 1621261055
transform 1 0 33696 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_347
timestamp 1621261055
transform 1 0 34464 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_355
timestamp 1621261055
transform 1 0 35232 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_363
timestamp 1621261055
transform 1 0 36000 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _044_
timestamp 1621261055
transform 1 0 36672 0 1 37962
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_737
timestamp 1621261055
transform 1 0 38112 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_367
timestamp 1621261055
transform 1 0 36384 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_53_369
timestamp 1621261055
transform 1 0 36576 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_373
timestamp 1621261055
transform 1 0 36960 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_381
timestamp 1621261055
transform 1 0 37728 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_53_386
timestamp 1621261055
transform 1 0 38208 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_394
timestamp 1621261055
transform 1 0 38976 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_402
timestamp 1621261055
transform 1 0 39744 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_410
timestamp 1621261055
transform 1 0 40512 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_418
timestamp 1621261055
transform 1 0 41280 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_426
timestamp 1621261055
transform 1 0 42048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_738
timestamp 1621261055
transform 1 0 43392 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_53_434
timestamp 1621261055
transform 1 0 42816 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_438
timestamp 1621261055
transform 1 0 43200 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_441
timestamp 1621261055
transform 1 0 43488 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_449
timestamp 1621261055
transform 1 0 44256 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_457
timestamp 1621261055
transform 1 0 45024 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_739
timestamp 1621261055
transform 1 0 48672 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_465
timestamp 1621261055
transform 1 0 45792 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_473
timestamp 1621261055
transform 1 0 46560 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_481
timestamp 1621261055
transform 1 0 47328 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_489
timestamp 1621261055
transform 1 0 48096 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_493
timestamp 1621261055
transform 1 0 48480 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_496
timestamp 1621261055
transform 1 0 48768 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_504
timestamp 1621261055
transform 1 0 49536 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_512
timestamp 1621261055
transform 1 0 50304 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_520
timestamp 1621261055
transform 1 0 51072 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_528
timestamp 1621261055
transform 1 0 51840 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_740
timestamp 1621261055
transform 1 0 53952 0 1 37962
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_53_536
timestamp 1621261055
transform 1 0 52608 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_544
timestamp 1621261055
transform 1 0 53376 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_548
timestamp 1621261055
transform 1 0 53760 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_53_551
timestamp 1621261055
transform 1 0 54048 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_559
timestamp 1621261055
transform 1 0 54816 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_567
timestamp 1621261055
transform 1 0 55584 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_575
timestamp 1621261055
transform 1 0 56352 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_53_583
timestamp 1621261055
transform 1 0 57120 0 1 37962
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_53_591
timestamp 1621261055
transform 1 0 57888 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_107
timestamp 1621261055
transform -1 0 58848 0 1 37962
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_53_595
timestamp 1621261055
transform 1 0 58272 0 1 37962
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_4
timestamp 1621261055
transform 1 0 1536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_4
timestamp 1621261055
transform 1 0 1536 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_110
timestamp 1621261055
transform 1 0 1152 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_108
timestamp 1621261055
transform 1 0 1152 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_12
timestamp 1621261055
transform 1 0 2304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_12
timestamp 1621261055
transform 1 0 2304 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_20
timestamp 1621261055
transform 1 0 3072 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_20
timestamp 1621261055
transform 1 0 3072 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_28
timestamp 1621261055
transform 1 0 3840 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_29
timestamp 1621261055
transform 1 0 3936 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_741
timestamp 1621261055
transform 1 0 3840 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_36
timestamp 1621261055
transform 1 0 4608 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_37
timestamp 1621261055
transform 1 0 4704 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_44
timestamp 1621261055
transform 1 0 5376 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_45
timestamp 1621261055
transform 1 0 5472 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_56
timestamp 1621261055
transform 1 0 6528 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_55_54
timestamp 1621261055
transform 1 0 6336 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_52
timestamp 1621261055
transform 1 0 6144 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_53
timestamp 1621261055
transform 1 0 6240 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_752
timestamp 1621261055
transform 1 0 6432 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_64
timestamp 1621261055
transform 1 0 7296 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_61
timestamp 1621261055
transform 1 0 7008 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_72
timestamp 1621261055
transform 1 0 8064 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_69
timestamp 1621261055
transform 1 0 7776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_80
timestamp 1621261055
transform 1 0 8832 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_81
timestamp 1621261055
transform 1 0 8928 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_77
timestamp 1621261055
transform 1 0 8544 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_742
timestamp 1621261055
transform 1 0 9120 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_88
timestamp 1621261055
transform 1 0 9600 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_92
timestamp 1621261055
transform 1 0 9984 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_84
timestamp 1621261055
transform 1 0 9216 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_96
timestamp 1621261055
transform 1 0 10368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_104
timestamp 1621261055
transform 1 0 11136 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_100
timestamp 1621261055
transform 1 0 10752 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_111
timestamp 1621261055
transform 1 0 11808 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_108
timestamp 1621261055
transform 1 0 11520 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_116
timestamp 1621261055
transform 1 0 12288 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_108
timestamp 1621261055
transform 1 0 11520 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_753
timestamp 1621261055
transform 1 0 11712 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_119
timestamp 1621261055
transform 1 0 12576 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_124
timestamp 1621261055
transform 1 0 13056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_127
timestamp 1621261055
transform 1 0 13344 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_132
timestamp 1621261055
transform 1 0 13824 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_135
timestamp 1621261055
transform 1 0 14112 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_139
timestamp 1621261055
transform 1 0 14496 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_136
timestamp 1621261055
transform 1 0 14208 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_743
timestamp 1621261055
transform 1 0 14400 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_143
timestamp 1621261055
transform 1 0 14880 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_147
timestamp 1621261055
transform 1 0 15264 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_151
timestamp 1621261055
transform 1 0 15648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_155
timestamp 1621261055
transform 1 0 16032 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_163
timestamp 1621261055
transform 1 0 16800 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_159
timestamp 1621261055
transform 1 0 16416 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_163
timestamp 1621261055
transform 1 0 16800 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_754
timestamp 1621261055
transform 1 0 16992 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_166
timestamp 1621261055
transform 1 0 17088 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_171
timestamp 1621261055
transform 1 0 17568 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_182
timestamp 1621261055
transform 1 0 18624 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_174
timestamp 1621261055
transform 1 0 17856 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_179
timestamp 1621261055
transform 1 0 18336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_190
timestamp 1621261055
transform 1 0 19392 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_191
timestamp 1621261055
transform 1 0 19488 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_187
timestamp 1621261055
transform 1 0 19104 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_198
timestamp 1621261055
transform 1 0 20160 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_194
timestamp 1621261055
transform 1 0 19776 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_744
timestamp 1621261055
transform 1 0 19680 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_206
timestamp 1621261055
transform 1 0 20928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_202
timestamp 1621261055
transform 1 0 20544 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_214
timestamp 1621261055
transform 1 0 21696 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_210
timestamp 1621261055
transform 1 0 21312 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_221
timestamp 1621261055
transform 1 0 22368 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_218
timestamp 1621261055
transform 1 0 22080 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_218
timestamp 1621261055
transform 1 0 22080 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_755
timestamp 1621261055
transform 1 0 22272 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_229
timestamp 1621261055
transform 1 0 23136 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_226
timestamp 1621261055
transform 1 0 22848 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_237
timestamp 1621261055
transform 1 0 23904 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_234
timestamp 1621261055
transform 1 0 23616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_245
timestamp 1621261055
transform 1 0 24672 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_246
timestamp 1621261055
transform 1 0 24768 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_242
timestamp 1621261055
transform 1 0 24384 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_745
timestamp 1621261055
transform 1 0 24960 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_253
timestamp 1621261055
transform 1 0 25440 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_257
timestamp 1621261055
transform 1 0 25824 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_249
timestamp 1621261055
transform 1 0 25056 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_261
timestamp 1621261055
transform 1 0 26208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_269
timestamp 1621261055
transform 1 0 26976 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_265
timestamp 1621261055
transform 1 0 26592 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_276
timestamp 1621261055
transform 1 0 27648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_273
timestamp 1621261055
transform 1 0 27360 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_281
timestamp 1621261055
transform 1 0 28128 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_273
timestamp 1621261055
transform 1 0 27360 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_756
timestamp 1621261055
transform 1 0 27552 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_284
timestamp 1621261055
transform 1 0 28416 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_289
timestamp 1621261055
transform 1 0 28896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_292
timestamp 1621261055
transform 1 0 29184 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_297
timestamp 1621261055
transform 1 0 29664 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_300
timestamp 1621261055
transform 1 0 29952 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_304
timestamp 1621261055
transform 1 0 30336 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_301
timestamp 1621261055
transform 1 0 30048 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_746
timestamp 1621261055
transform 1 0 30240 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_308
timestamp 1621261055
transform 1 0 30720 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_312
timestamp 1621261055
transform 1 0 31104 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_316
timestamp 1621261055
transform 1 0 31488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_323
timestamp 1621261055
transform 1 0 32160 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _024_
timestamp 1621261055
transform 1 0 31872 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_328
timestamp 1621261055
transform 1 0 32640 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_55_324
timestamp 1621261055
transform 1 0 32256 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_757
timestamp 1621261055
transform 1 0 32832 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_331
timestamp 1621261055
transform 1 0 32928 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_331
timestamp 1621261055
transform 1 0 32928 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_347
timestamp 1621261055
transform 1 0 34464 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_339
timestamp 1621261055
transform 1 0 33696 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_343
timestamp 1621261055
transform 1 0 34080 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_54_339
timestamp 1621261055
transform 1 0 33696 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_194
timestamp 1621261055
transform 1 0 34176 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _121_
timestamp 1621261055
transform 1 0 34368 0 -1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_55_355
timestamp 1621261055
transform 1 0 35232 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_349
timestamp 1621261055
transform 1 0 34656 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_363
timestamp 1621261055
transform 1 0 36000 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_359
timestamp 1621261055
transform 1 0 35616 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_54_357
timestamp 1621261055
transform 1 0 35424 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_747
timestamp 1621261055
transform 1 0 35520 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_371
timestamp 1621261055
transform 1 0 36768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_367
timestamp 1621261055
transform 1 0 36384 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_379
timestamp 1621261055
transform 1 0 37536 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_375
timestamp 1621261055
transform 1 0 37152 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_386
timestamp 1621261055
transform 1 0 38208 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_383
timestamp 1621261055
transform 1 0 37920 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_383
timestamp 1621261055
transform 1 0 37920 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_758
timestamp 1621261055
transform 1 0 38112 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_394
timestamp 1621261055
transform 1 0 38976 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_391
timestamp 1621261055
transform 1 0 38688 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_402
timestamp 1621261055
transform 1 0 39744 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_399
timestamp 1621261055
transform 1 0 39456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_410
timestamp 1621261055
transform 1 0 40512 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_411
timestamp 1621261055
transform 1 0 40608 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_407
timestamp 1621261055
transform 1 0 40224 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_748
timestamp 1621261055
transform 1 0 40800 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_418
timestamp 1621261055
transform 1 0 41280 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_422
timestamp 1621261055
transform 1 0 41664 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_414
timestamp 1621261055
transform 1 0 40896 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_426
timestamp 1621261055
transform 1 0 42048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_434
timestamp 1621261055
transform 1 0 42816 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_430
timestamp 1621261055
transform 1 0 42432 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_441
timestamp 1621261055
transform 1 0 43488 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_438
timestamp 1621261055
transform 1 0 43200 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_54_446
timestamp 1621261055
transform 1 0 43968 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_438
timestamp 1621261055
transform 1 0 43200 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_759
timestamp 1621261055
transform 1 0 43392 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_449
timestamp 1621261055
transform 1 0 44256 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_454
timestamp 1621261055
transform 1 0 44736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_457
timestamp 1621261055
transform 1 0 45024 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_54_462
timestamp 1621261055
transform 1 0 45504 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_55_465
timestamp 1621261055
transform 1 0 45792 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_469
timestamp 1621261055
transform 1 0 46176 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_466
timestamp 1621261055
transform 1 0 45888 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_749
timestamp 1621261055
transform 1 0 46080 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_473
timestamp 1621261055
transform 1 0 46560 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_477
timestamp 1621261055
transform 1 0 46944 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_55_485
timestamp 1621261055
transform 1 0 47712 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_55_481
timestamp 1621261055
transform 1 0 47328 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_485
timestamp 1621261055
transform 1 0 47712 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_140
timestamp 1621261055
transform 1 0 47808 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _179_
timestamp 1621261055
transform 1 0 48000 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_55_491
timestamp 1621261055
transform 1 0 48288 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_54_493
timestamp 1621261055
transform 1 0 48480 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_760
timestamp 1621261055
transform 1 0 48672 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_496
timestamp 1621261055
transform 1 0 48768 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_501
timestamp 1621261055
transform 1 0 49248 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_512
timestamp 1621261055
transform 1 0 50304 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_504
timestamp 1621261055
transform 1 0 49536 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_509
timestamp 1621261055
transform 1 0 50016 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_55_520
timestamp 1621261055
transform 1 0 51072 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_521
timestamp 1621261055
transform 1 0 51168 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_517
timestamp 1621261055
transform 1 0 50784 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_111
timestamp 1621261055
transform 1 0 51168 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_55_526
timestamp 1621261055
transform 1 0 51648 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_524
timestamp 1621261055
transform 1 0 51456 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_750
timestamp 1621261055
transform 1 0 51360 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _162_
timestamp 1621261055
transform 1 0 51360 0 1 39294
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_761
timestamp 1621261055
transform 1 0 53952 0 1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_54_532
timestamp 1621261055
transform 1 0 52224 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_540
timestamp 1621261055
transform 1 0 52992 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_548
timestamp 1621261055
transform 1 0 53760 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_556
timestamp 1621261055
transform 1 0 54528 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_534
timestamp 1621261055
transform 1 0 52416 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_542
timestamp 1621261055
transform 1 0 53184 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_551
timestamp 1621261055
transform 1 0 54048 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_559
timestamp 1621261055
transform 1 0 54816 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_567
timestamp 1621261055
transform 1 0 55584 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_564
timestamp 1621261055
transform 1 0 55296 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_55_575
timestamp 1621261055
transform 1 0 56352 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_576
timestamp 1621261055
transform 1 0 56448 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_54_572
timestamp 1621261055
transform 1 0 56064 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_751
timestamp 1621261055
transform 1 0 56640 0 -1 39294
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_55_583
timestamp 1621261055
transform 1 0 57120 0 1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_587
timestamp 1621261055
transform 1 0 57504 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_54_579
timestamp 1621261055
transform 1 0 56736 0 -1 39294
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_55_591
timestamp 1621261055
transform 1 0 57888 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_109
timestamp 1621261055
transform -1 0 58848 0 -1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_111
timestamp 1621261055
transform -1 0 58848 0 1 39294
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_54_595
timestamp 1621261055
transform 1 0 58272 0 -1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_55_595
timestamp 1621261055
transform 1 0 58272 0 1 39294
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_112
timestamp 1621261055
transform 1 0 1152 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_762
timestamp 1621261055
transform 1 0 3840 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_4
timestamp 1621261055
transform 1 0 1536 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_12
timestamp 1621261055
transform 1 0 2304 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_20
timestamp 1621261055
transform 1 0 3072 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_29
timestamp 1621261055
transform 1 0 3936 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_37
timestamp 1621261055
transform 1 0 4704 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_45
timestamp 1621261055
transform 1 0 5472 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_53
timestamp 1621261055
transform 1 0 6240 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_61
timestamp 1621261055
transform 1 0 7008 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_763
timestamp 1621261055
transform 1 0 9120 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_69
timestamp 1621261055
transform 1 0 7776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_77
timestamp 1621261055
transform 1 0 8544 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_81
timestamp 1621261055
transform 1 0 8928 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_84
timestamp 1621261055
transform 1 0 9216 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_92
timestamp 1621261055
transform 1 0 9984 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_100
timestamp 1621261055
transform 1 0 10752 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_108
timestamp 1621261055
transform 1 0 11520 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_116
timestamp 1621261055
transform 1 0 12288 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_124
timestamp 1621261055
transform 1 0 13056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_132
timestamp 1621261055
transform 1 0 13824 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _021_
timestamp 1621261055
transform 1 0 16512 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_764
timestamp 1621261055
transform 1 0 14400 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_213
timestamp 1621261055
transform -1 0 17184 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_136
timestamp 1621261055
transform 1 0 14208 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_139
timestamp 1621261055
transform 1 0 14496 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_147
timestamp 1621261055
transform 1 0 15264 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_155
timestamp 1621261055
transform 1 0 16032 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_56_159
timestamp 1621261055
transform 1 0 16416 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_163
timestamp 1621261055
transform 1 0 16800 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _065_
timestamp 1621261055
transform -1 0 17472 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_765
timestamp 1621261055
transform 1 0 19680 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_170
timestamp 1621261055
transform 1 0 17472 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_178
timestamp 1621261055
transform 1 0 18240 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_186
timestamp 1621261055
transform 1 0 19008 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_190
timestamp 1621261055
transform 1 0 19392 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_192
timestamp 1621261055
transform 1 0 19584 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_194
timestamp 1621261055
transform 1 0 19776 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_258
timestamp 1621261055
transform -1 0 23520 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_202
timestamp 1621261055
transform 1 0 20544 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_210
timestamp 1621261055
transform 1 0 21312 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_218
timestamp 1621261055
transform 1 0 22080 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_226
timestamp 1621261055
transform 1 0 22848 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_56_230
timestamp 1621261055
transform 1 0 23232 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _188_
timestamp 1621261055
transform -1 0 23808 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_766
timestamp 1621261055
transform 1 0 24960 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_236
timestamp 1621261055
transform 1 0 23808 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_244
timestamp 1621261055
transform 1 0 24576 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_56_249
timestamp 1621261055
transform 1 0 25056 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_257
timestamp 1621261055
transform 1 0 25824 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_265
timestamp 1621261055
transform 1 0 26592 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_273
timestamp 1621261055
transform 1 0 27360 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_281
timestamp 1621261055
transform 1 0 28128 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_289
timestamp 1621261055
transform 1 0 28896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_297
timestamp 1621261055
transform 1 0 29664 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_767
timestamp 1621261055
transform 1 0 30240 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_301
timestamp 1621261055
transform 1 0 30048 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_304
timestamp 1621261055
transform 1 0 30336 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_312
timestamp 1621261055
transform 1 0 31104 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_320
timestamp 1621261055
transform 1 0 31872 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_328
timestamp 1621261055
transform 1 0 32640 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_768
timestamp 1621261055
transform 1 0 35520 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_336
timestamp 1621261055
transform 1 0 33408 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_344
timestamp 1621261055
transform 1 0 34176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_352
timestamp 1621261055
transform 1 0 34944 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_356
timestamp 1621261055
transform 1 0 35328 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_359
timestamp 1621261055
transform 1 0 35616 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_367
timestamp 1621261055
transform 1 0 36384 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_375
timestamp 1621261055
transform 1 0 37152 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_383
timestamp 1621261055
transform 1 0 37920 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_391
timestamp 1621261055
transform 1 0 38688 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_769
timestamp 1621261055
transform 1 0 40800 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_399
timestamp 1621261055
transform 1 0 39456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_407
timestamp 1621261055
transform 1 0 40224 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_411
timestamp 1621261055
transform 1 0 40608 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_414
timestamp 1621261055
transform 1 0 40896 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_422
timestamp 1621261055
transform 1 0 41664 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_430
timestamp 1621261055
transform 1 0 42432 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_438
timestamp 1621261055
transform 1 0 43200 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_446
timestamp 1621261055
transform 1 0 43968 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_454
timestamp 1621261055
transform 1 0 44736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_462
timestamp 1621261055
transform 1 0 45504 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _064_
timestamp 1621261055
transform -1 0 47712 0 -1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_770
timestamp 1621261055
transform 1 0 46080 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_202
timestamp 1621261055
transform -1 0 47424 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_466
timestamp 1621261055
transform 1 0 45888 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_469
timestamp 1621261055
transform 1 0 46176 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_477
timestamp 1621261055
transform 1 0 46944 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_56_479
timestamp 1621261055
transform 1 0 47136 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_485
timestamp 1621261055
transform 1 0 47712 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_493
timestamp 1621261055
transform 1 0 48480 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_771
timestamp 1621261055
transform 1 0 51360 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_501
timestamp 1621261055
transform 1 0 49248 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_509
timestamp 1621261055
transform 1 0 50016 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_517
timestamp 1621261055
transform 1 0 50784 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_521
timestamp 1621261055
transform 1 0 51168 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_524
timestamp 1621261055
transform 1 0 51456 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_532
timestamp 1621261055
transform 1 0 52224 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_540
timestamp 1621261055
transform 1 0 52992 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_548
timestamp 1621261055
transform 1 0 53760 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_556
timestamp 1621261055
transform 1 0 54528 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_772
timestamp 1621261055
transform 1 0 56640 0 -1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_56_564
timestamp 1621261055
transform 1 0 55296 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_56_572
timestamp 1621261055
transform 1 0 56064 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_576
timestamp 1621261055
transform 1 0 56448 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_56_579
timestamp 1621261055
transform 1 0 56736 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_56_587
timestamp 1621261055
transform 1 0 57504 0 -1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_113
timestamp 1621261055
transform -1 0 58848 0 -1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_56_595
timestamp 1621261055
transform 1 0 58272 0 -1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_114
timestamp 1621261055
transform 1 0 1152 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_57_4
timestamp 1621261055
transform 1 0 1536 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_12
timestamp 1621261055
transform 1 0 2304 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_20
timestamp 1621261055
transform 1 0 3072 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_28
timestamp 1621261055
transform 1 0 3840 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_773
timestamp 1621261055
transform 1 0 6432 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_36
timestamp 1621261055
transform 1 0 4608 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_44
timestamp 1621261055
transform 1 0 5376 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_52
timestamp 1621261055
transform 1 0 6144 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_54
timestamp 1621261055
transform 1 0 6336 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_56
timestamp 1621261055
transform 1 0 6528 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_64
timestamp 1621261055
transform 1 0 7296 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_72
timestamp 1621261055
transform 1 0 8064 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_80
timestamp 1621261055
transform 1 0 8832 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_88
timestamp 1621261055
transform 1 0 9600 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_96
timestamp 1621261055
transform 1 0 10368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_774
timestamp 1621261055
transform 1 0 11712 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_104
timestamp 1621261055
transform 1 0 11136 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_108
timestamp 1621261055
transform 1 0 11520 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_111
timestamp 1621261055
transform 1 0 11808 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_119
timestamp 1621261055
transform 1 0 12576 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_127
timestamp 1621261055
transform 1 0 13344 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_775
timestamp 1621261055
transform 1 0 16992 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_135
timestamp 1621261055
transform 1 0 14112 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_143
timestamp 1621261055
transform 1 0 14880 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_151
timestamp 1621261055
transform 1 0 15648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_159
timestamp 1621261055
transform 1 0 16416 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_163
timestamp 1621261055
transform 1 0 16800 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_166
timestamp 1621261055
transform 1 0 17088 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_174
timestamp 1621261055
transform 1 0 17856 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_182
timestamp 1621261055
transform 1 0 18624 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_190
timestamp 1621261055
transform 1 0 19392 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_198
timestamp 1621261055
transform 1 0 20160 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_776
timestamp 1621261055
transform 1 0 22272 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_206
timestamp 1621261055
transform 1 0 20928 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_214
timestamp 1621261055
transform 1 0 21696 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_218
timestamp 1621261055
transform 1 0 22080 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_221
timestamp 1621261055
transform 1 0 22368 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_229
timestamp 1621261055
transform 1 0 23136 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_237
timestamp 1621261055
transform 1 0 23904 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_245
timestamp 1621261055
transform 1 0 24672 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_253
timestamp 1621261055
transform 1 0 25440 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_261
timestamp 1621261055
transform 1 0 26208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_777
timestamp 1621261055
transform 1 0 27552 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_269
timestamp 1621261055
transform 1 0 26976 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_273
timestamp 1621261055
transform 1 0 27360 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_276
timestamp 1621261055
transform 1 0 27648 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_284
timestamp 1621261055
transform 1 0 28416 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_292
timestamp 1621261055
transform 1 0 29184 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_778
timestamp 1621261055
transform 1 0 32832 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_300
timestamp 1621261055
transform 1 0 29952 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_308
timestamp 1621261055
transform 1 0 30720 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_316
timestamp 1621261055
transform 1 0 31488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_324
timestamp 1621261055
transform 1 0 32256 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_328
timestamp 1621261055
transform 1 0 32640 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _208_
timestamp 1621261055
transform -1 0 34080 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_250
timestamp 1621261055
transform -1 0 33792 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_57_331
timestamp 1621261055
transform 1 0 32928 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_335
timestamp 1621261055
transform 1 0 33312 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_337
timestamp 1621261055
transform 1 0 33504 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_343
timestamp 1621261055
transform 1 0 34080 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_351
timestamp 1621261055
transform 1 0 34848 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_359
timestamp 1621261055
transform 1 0 35616 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_779
timestamp 1621261055
transform 1 0 38112 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_367
timestamp 1621261055
transform 1 0 36384 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_375
timestamp 1621261055
transform 1 0 37152 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_383
timestamp 1621261055
transform 1 0 37920 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_386
timestamp 1621261055
transform 1 0 38208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_394
timestamp 1621261055
transform 1 0 38976 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_402
timestamp 1621261055
transform 1 0 39744 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_410
timestamp 1621261055
transform 1 0 40512 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_418
timestamp 1621261055
transform 1 0 41280 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_426
timestamp 1621261055
transform 1 0 42048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_780
timestamp 1621261055
transform 1 0 43392 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_57_434
timestamp 1621261055
transform 1 0 42816 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_438
timestamp 1621261055
transform 1 0 43200 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_441
timestamp 1621261055
transform 1 0 43488 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_449
timestamp 1621261055
transform 1 0 44256 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_457
timestamp 1621261055
transform 1 0 45024 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_781
timestamp 1621261055
transform 1 0 48672 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_465
timestamp 1621261055
transform 1 0 45792 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_473
timestamp 1621261055
transform 1 0 46560 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_481
timestamp 1621261055
transform 1 0 47328 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_489
timestamp 1621261055
transform 1 0 48096 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_493
timestamp 1621261055
transform 1 0 48480 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _070_
timestamp 1621261055
transform -1 0 50208 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_143
timestamp 1621261055
transform -1 0 49920 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_496
timestamp 1621261055
transform 1 0 48768 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_504
timestamp 1621261055
transform 1 0 49536 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_57_511
timestamp 1621261055
transform 1 0 50208 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_519
timestamp 1621261055
transform 1 0 50976 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_527
timestamp 1621261055
transform 1 0 51744 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_782
timestamp 1621261055
transform 1 0 53952 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_535
timestamp 1621261055
transform 1 0 52512 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_543
timestamp 1621261055
transform 1 0 53280 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_547
timestamp 1621261055
transform 1 0 53664 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_57_549
timestamp 1621261055
transform 1 0 53856 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_57_551
timestamp 1621261055
transform 1 0 54048 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_559
timestamp 1621261055
transform 1 0 54816 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _007_
timestamp 1621261055
transform 1 0 57696 0 1 40626
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_57_567
timestamp 1621261055
transform 1 0 55584 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_57_575
timestamp 1621261055
transform 1 0 56352 0 1 40626
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_57_583
timestamp 1621261055
transform 1 0 57120 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_57_587
timestamp 1621261055
transform 1 0 57504 0 1 40626
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_57_592
timestamp 1621261055
transform 1 0 57984 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_115
timestamp 1621261055
transform -1 0 58848 0 1 40626
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_57_596
timestamp 1621261055
transform 1 0 58368 0 1 40626
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  PHY_116
timestamp 1621261055
transform 1 0 1152 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_783
timestamp 1621261055
transform 1 0 3840 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_4
timestamp 1621261055
transform 1 0 1536 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_12
timestamp 1621261055
transform 1 0 2304 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_20
timestamp 1621261055
transform 1 0 3072 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_29
timestamp 1621261055
transform 1 0 3936 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_37
timestamp 1621261055
transform 1 0 4704 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_45
timestamp 1621261055
transform 1 0 5472 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_53
timestamp 1621261055
transform 1 0 6240 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_61
timestamp 1621261055
transform 1 0 7008 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_784
timestamp 1621261055
transform 1 0 9120 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_69
timestamp 1621261055
transform 1 0 7776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_77
timestamp 1621261055
transform 1 0 8544 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_81
timestamp 1621261055
transform 1 0 8928 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_84
timestamp 1621261055
transform 1 0 9216 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_92
timestamp 1621261055
transform 1 0 9984 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_100
timestamp 1621261055
transform 1 0 10752 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_108
timestamp 1621261055
transform 1 0 11520 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_116
timestamp 1621261055
transform 1 0 12288 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_124
timestamp 1621261055
transform 1 0 13056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_132
timestamp 1621261055
transform 1 0 13824 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_785
timestamp 1621261055
transform 1 0 14400 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_136
timestamp 1621261055
transform 1 0 14208 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_139
timestamp 1621261055
transform 1 0 14496 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_147
timestamp 1621261055
transform 1 0 15264 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_155
timestamp 1621261055
transform 1 0 16032 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_163
timestamp 1621261055
transform 1 0 16800 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_786
timestamp 1621261055
transform 1 0 19680 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_171
timestamp 1621261055
transform 1 0 17568 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_179
timestamp 1621261055
transform 1 0 18336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_187
timestamp 1621261055
transform 1 0 19104 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_191
timestamp 1621261055
transform 1 0 19488 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_194
timestamp 1621261055
transform 1 0 19776 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_202
timestamp 1621261055
transform 1 0 20544 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_210
timestamp 1621261055
transform 1 0 21312 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_218
timestamp 1621261055
transform 1 0 22080 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_226
timestamp 1621261055
transform 1 0 22848 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_787
timestamp 1621261055
transform 1 0 24960 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_234
timestamp 1621261055
transform 1 0 23616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_242
timestamp 1621261055
transform 1 0 24384 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_246
timestamp 1621261055
transform 1 0 24768 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_249
timestamp 1621261055
transform 1 0 25056 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_257
timestamp 1621261055
transform 1 0 25824 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_265
timestamp 1621261055
transform 1 0 26592 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_273
timestamp 1621261055
transform 1 0 27360 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_281
timestamp 1621261055
transform 1 0 28128 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_289
timestamp 1621261055
transform 1 0 28896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_297
timestamp 1621261055
transform 1 0 29664 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_788
timestamp 1621261055
transform 1 0 30240 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_301
timestamp 1621261055
transform 1 0 30048 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_304
timestamp 1621261055
transform 1 0 30336 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_312
timestamp 1621261055
transform 1 0 31104 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_320
timestamp 1621261055
transform 1 0 31872 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_328
timestamp 1621261055
transform 1 0 32640 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_789
timestamp 1621261055
transform 1 0 35520 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_336
timestamp 1621261055
transform 1 0 33408 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_344
timestamp 1621261055
transform 1 0 34176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_352
timestamp 1621261055
transform 1 0 34944 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_356
timestamp 1621261055
transform 1 0 35328 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_359
timestamp 1621261055
transform 1 0 35616 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_367
timestamp 1621261055
transform 1 0 36384 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_375
timestamp 1621261055
transform 1 0 37152 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_383
timestamp 1621261055
transform 1 0 37920 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_391
timestamp 1621261055
transform 1 0 38688 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_790
timestamp 1621261055
transform 1 0 40800 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_399
timestamp 1621261055
transform 1 0 39456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_407
timestamp 1621261055
transform 1 0 40224 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_411
timestamp 1621261055
transform 1 0 40608 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_414
timestamp 1621261055
transform 1 0 40896 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_422
timestamp 1621261055
transform 1 0 41664 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_430
timestamp 1621261055
transform 1 0 42432 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_438
timestamp 1621261055
transform 1 0 43200 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_446
timestamp 1621261055
transform 1 0 43968 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_454
timestamp 1621261055
transform 1 0 44736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_462
timestamp 1621261055
transform 1 0 45504 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_791
timestamp 1621261055
transform 1 0 46080 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_466
timestamp 1621261055
transform 1 0 45888 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_469
timestamp 1621261055
transform 1 0 46176 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_477
timestamp 1621261055
transform 1 0 46944 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_485
timestamp 1621261055
transform 1 0 47712 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_493
timestamp 1621261055
transform 1 0 48480 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_792
timestamp 1621261055
transform 1 0 51360 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_501
timestamp 1621261055
transform 1 0 49248 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_509
timestamp 1621261055
transform 1 0 50016 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_517
timestamp 1621261055
transform 1 0 50784 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_521
timestamp 1621261055
transform 1 0 51168 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_524
timestamp 1621261055
transform 1 0 51456 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_532
timestamp 1621261055
transform 1 0 52224 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_540
timestamp 1621261055
transform 1 0 52992 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_548
timestamp 1621261055
transform 1 0 53760 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_556
timestamp 1621261055
transform 1 0 54528 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_793
timestamp 1621261055
transform 1 0 56640 0 -1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_58_564
timestamp 1621261055
transform 1 0 55296 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_58_572
timestamp 1621261055
transform 1 0 56064 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_576
timestamp 1621261055
transform 1 0 56448 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_58_579
timestamp 1621261055
transform 1 0 56736 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_58_587
timestamp 1621261055
transform 1 0 57504 0 -1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_117
timestamp 1621261055
transform -1 0 58848 0 -1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_58_595
timestamp 1621261055
transform 1 0 58272 0 -1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _069_
timestamp 1621261055
transform 1 0 3360 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_118
timestamp 1621261055
transform 1 0 1152 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_59_4
timestamp 1621261055
transform 1 0 1536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_12
timestamp 1621261055
transform 1 0 2304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_20
timestamp 1621261055
transform 1 0 3072 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_22
timestamp 1621261055
transform 1 0 3264 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_26
timestamp 1621261055
transform 1 0 3648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_794
timestamp 1621261055
transform 1 0 6432 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_34
timestamp 1621261055
transform 1 0 4416 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_42
timestamp 1621261055
transform 1 0 5184 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_50
timestamp 1621261055
transform 1 0 5952 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_59_54
timestamp 1621261055
transform 1 0 6336 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_56
timestamp 1621261055
transform 1 0 6528 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_64
timestamp 1621261055
transform 1 0 7296 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_72
timestamp 1621261055
transform 1 0 8064 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_80
timestamp 1621261055
transform 1 0 8832 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_88
timestamp 1621261055
transform 1 0 9600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_96
timestamp 1621261055
transform 1 0 10368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_795
timestamp 1621261055
transform 1 0 11712 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_104
timestamp 1621261055
transform 1 0 11136 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_108
timestamp 1621261055
transform 1 0 11520 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_111
timestamp 1621261055
transform 1 0 11808 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_119
timestamp 1621261055
transform 1 0 12576 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_127
timestamp 1621261055
transform 1 0 13344 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_796
timestamp 1621261055
transform 1 0 16992 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_135
timestamp 1621261055
transform 1 0 14112 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_143
timestamp 1621261055
transform 1 0 14880 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_151
timestamp 1621261055
transform 1 0 15648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_159
timestamp 1621261055
transform 1 0 16416 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_163
timestamp 1621261055
transform 1 0 16800 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_166
timestamp 1621261055
transform 1 0 17088 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_174
timestamp 1621261055
transform 1 0 17856 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_182
timestamp 1621261055
transform 1 0 18624 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_190
timestamp 1621261055
transform 1 0 19392 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_198
timestamp 1621261055
transform 1 0 20160 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_797
timestamp 1621261055
transform 1 0 22272 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_206
timestamp 1621261055
transform 1 0 20928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_214
timestamp 1621261055
transform 1 0 21696 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_218
timestamp 1621261055
transform 1 0 22080 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_221
timestamp 1621261055
transform 1 0 22368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_229
timestamp 1621261055
transform 1 0 23136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_237
timestamp 1621261055
transform 1 0 23904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_245
timestamp 1621261055
transform 1 0 24672 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_253
timestamp 1621261055
transform 1 0 25440 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_261
timestamp 1621261055
transform 1 0 26208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_798
timestamp 1621261055
transform 1 0 27552 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_59_269
timestamp 1621261055
transform 1 0 26976 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_273
timestamp 1621261055
transform 1 0 27360 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_276
timestamp 1621261055
transform 1 0 27648 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_284
timestamp 1621261055
transform 1 0 28416 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_292
timestamp 1621261055
transform 1 0 29184 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_296
timestamp 1621261055
transform 1 0 29568 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _187_
timestamp 1621261055
transform -1 0 30240 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_799
timestamp 1621261055
transform 1 0 32832 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_256
timestamp 1621261055
transform -1 0 29952 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_303
timestamp 1621261055
transform 1 0 30240 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_311
timestamp 1621261055
transform 1 0 31008 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_319
timestamp 1621261055
transform 1 0 31776 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_327
timestamp 1621261055
transform 1 0 32544 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_59_329
timestamp 1621261055
transform 1 0 32736 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_331
timestamp 1621261055
transform 1 0 32928 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_339
timestamp 1621261055
transform 1 0 33696 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_347
timestamp 1621261055
transform 1 0 34464 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_355
timestamp 1621261055
transform 1 0 35232 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_363
timestamp 1621261055
transform 1 0 36000 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_800
timestamp 1621261055
transform 1 0 38112 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_371
timestamp 1621261055
transform 1 0 36768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_379
timestamp 1621261055
transform 1 0 37536 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_383
timestamp 1621261055
transform 1 0 37920 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_386
timestamp 1621261055
transform 1 0 38208 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_394
timestamp 1621261055
transform 1 0 38976 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_402
timestamp 1621261055
transform 1 0 39744 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_410
timestamp 1621261055
transform 1 0 40512 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_418
timestamp 1621261055
transform 1 0 41280 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_426
timestamp 1621261055
transform 1 0 42048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _137_
timestamp 1621261055
transform -1 0 45600 0 1 41958
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_801
timestamp 1621261055
transform 1 0 43392 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_208
timestamp 1621261055
transform -1 0 45312 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_59_434
timestamp 1621261055
transform 1 0 42816 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_438
timestamp 1621261055
transform 1 0 43200 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_441
timestamp 1621261055
transform 1 0 43488 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_449
timestamp 1621261055
transform 1 0 44256 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_59_457
timestamp 1621261055
transform 1 0 45024 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_802
timestamp 1621261055
transform 1 0 48672 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_463
timestamp 1621261055
transform 1 0 45600 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_471
timestamp 1621261055
transform 1 0 46368 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_479
timestamp 1621261055
transform 1 0 47136 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_487
timestamp 1621261055
transform 1 0 47904 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_496
timestamp 1621261055
transform 1 0 48768 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_504
timestamp 1621261055
transform 1 0 49536 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_512
timestamp 1621261055
transform 1 0 50304 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_520
timestamp 1621261055
transform 1 0 51072 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_528
timestamp 1621261055
transform 1 0 51840 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_803
timestamp 1621261055
transform 1 0 53952 0 1 41958
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_59_536
timestamp 1621261055
transform 1 0 52608 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_544
timestamp 1621261055
transform 1 0 53376 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_548
timestamp 1621261055
transform 1 0 53760 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_59_551
timestamp 1621261055
transform 1 0 54048 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_559
timestamp 1621261055
transform 1 0 54816 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_567
timestamp 1621261055
transform 1 0 55584 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_575
timestamp 1621261055
transform 1 0 56352 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_59_583
timestamp 1621261055
transform 1 0 57120 0 1 41958
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_59_591
timestamp 1621261055
transform 1 0 57888 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_119
timestamp 1621261055
transform -1 0 58848 0 1 41958
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_59_595
timestamp 1621261055
transform 1 0 58272 0 1 41958
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_120
timestamp 1621261055
transform 1 0 1152 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_804
timestamp 1621261055
transform 1 0 3840 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_4
timestamp 1621261055
transform 1 0 1536 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_12
timestamp 1621261055
transform 1 0 2304 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_20
timestamp 1621261055
transform 1 0 3072 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_29
timestamp 1621261055
transform 1 0 3936 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_37
timestamp 1621261055
transform 1 0 4704 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_45
timestamp 1621261055
transform 1 0 5472 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_53
timestamp 1621261055
transform 1 0 6240 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_61
timestamp 1621261055
transform 1 0 7008 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_805
timestamp 1621261055
transform 1 0 9120 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_69
timestamp 1621261055
transform 1 0 7776 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_77
timestamp 1621261055
transform 1 0 8544 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_81
timestamp 1621261055
transform 1 0 8928 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_84
timestamp 1621261055
transform 1 0 9216 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_92
timestamp 1621261055
transform 1 0 9984 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_100
timestamp 1621261055
transform 1 0 10752 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_108
timestamp 1621261055
transform 1 0 11520 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_116
timestamp 1621261055
transform 1 0 12288 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_124
timestamp 1621261055
transform 1 0 13056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_132
timestamp 1621261055
transform 1 0 13824 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _094_
timestamp 1621261055
transform 1 0 16224 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_806
timestamp 1621261055
transform 1 0 14400 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_171
timestamp 1621261055
transform 1 0 16032 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_136
timestamp 1621261055
transform 1 0 14208 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_139
timestamp 1621261055
transform 1 0 14496 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_147
timestamp 1621261055
transform 1 0 15264 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_160
timestamp 1621261055
transform 1 0 16512 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _204_
timestamp 1621261055
transform -1 0 20448 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_807
timestamp 1621261055
transform 1 0 19680 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_242
timestamp 1621261055
transform -1 0 20160 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_168
timestamp 1621261055
transform 1 0 17280 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_176
timestamp 1621261055
transform 1 0 18048 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_184
timestamp 1621261055
transform 1 0 18816 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_60_192
timestamp 1621261055
transform 1 0 19584 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_194
timestamp 1621261055
transform 1 0 19776 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _074_
timestamp 1621261055
transform -1 0 23136 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_147
timestamp 1621261055
transform -1 0 22848 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_201
timestamp 1621261055
transform 1 0 20448 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_209
timestamp 1621261055
transform 1 0 21216 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_217
timestamp 1621261055
transform 1 0 21984 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_221
timestamp 1621261055
transform 1 0 22368 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_223
timestamp 1621261055
transform 1 0 22560 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_229
timestamp 1621261055
transform 1 0 23136 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_808
timestamp 1621261055
transform 1 0 24960 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_237
timestamp 1621261055
transform 1 0 23904 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_245
timestamp 1621261055
transform 1 0 24672 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_247
timestamp 1621261055
transform 1 0 24864 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_249
timestamp 1621261055
transform 1 0 25056 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_257
timestamp 1621261055
transform 1 0 25824 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_265
timestamp 1621261055
transform 1 0 26592 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_273
timestamp 1621261055
transform 1 0 27360 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_281
timestamp 1621261055
transform 1 0 28128 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_289
timestamp 1621261055
transform 1 0 28896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_297
timestamp 1621261055
transform 1 0 29664 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_809
timestamp 1621261055
transform 1 0 30240 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_301
timestamp 1621261055
transform 1 0 30048 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_304
timestamp 1621261055
transform 1 0 30336 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_312
timestamp 1621261055
transform 1 0 31104 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_320
timestamp 1621261055
transform 1 0 31872 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_328
timestamp 1621261055
transform 1 0 32640 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_810
timestamp 1621261055
transform 1 0 35520 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_336
timestamp 1621261055
transform 1 0 33408 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_344
timestamp 1621261055
transform 1 0 34176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_352
timestamp 1621261055
transform 1 0 34944 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_356
timestamp 1621261055
transform 1 0 35328 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_359
timestamp 1621261055
transform 1 0 35616 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_367
timestamp 1621261055
transform 1 0 36384 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_375
timestamp 1621261055
transform 1 0 37152 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_383
timestamp 1621261055
transform 1 0 37920 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_391
timestamp 1621261055
transform 1 0 38688 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_811
timestamp 1621261055
transform 1 0 40800 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_399
timestamp 1621261055
transform 1 0 39456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_407
timestamp 1621261055
transform 1 0 40224 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_411
timestamp 1621261055
transform 1 0 40608 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_414
timestamp 1621261055
transform 1 0 40896 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_422
timestamp 1621261055
transform 1 0 41664 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_430
timestamp 1621261055
transform 1 0 42432 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_438
timestamp 1621261055
transform 1 0 43200 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_446
timestamp 1621261055
transform 1 0 43968 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_454
timestamp 1621261055
transform 1 0 44736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_462
timestamp 1621261055
transform 1 0 45504 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_812
timestamp 1621261055
transform 1 0 46080 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_466
timestamp 1621261055
transform 1 0 45888 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_469
timestamp 1621261055
transform 1 0 46176 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_477
timestamp 1621261055
transform 1 0 46944 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_485
timestamp 1621261055
transform 1 0 47712 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_493
timestamp 1621261055
transform 1 0 48480 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_813
timestamp 1621261055
transform 1 0 51360 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_501
timestamp 1621261055
transform 1 0 49248 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_509
timestamp 1621261055
transform 1 0 50016 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_517
timestamp 1621261055
transform 1 0 50784 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_521
timestamp 1621261055
transform 1 0 51168 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_524
timestamp 1621261055
transform 1 0 51456 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _143_
timestamp 1621261055
transform -1 0 52992 0 -1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_215
timestamp 1621261055
transform -1 0 52704 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_532
timestamp 1621261055
transform 1 0 52224 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_60_534
timestamp 1621261055
transform 1 0 52416 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_540
timestamp 1621261055
transform 1 0 52992 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_548
timestamp 1621261055
transform 1 0 53760 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_556
timestamp 1621261055
transform 1 0 54528 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_814
timestamp 1621261055
transform 1 0 56640 0 -1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_60_564
timestamp 1621261055
transform 1 0 55296 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_60_572
timestamp 1621261055
transform 1 0 56064 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_576
timestamp 1621261055
transform 1 0 56448 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_60_579
timestamp 1621261055
transform 1 0 56736 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_60_587
timestamp 1621261055
transform 1 0 57504 0 -1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_121
timestamp 1621261055
transform -1 0 58848 0 -1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_60_595
timestamp 1621261055
transform 1 0 58272 0 -1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_62_4
timestamp 1621261055
transform 1 0 1536 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_4
timestamp 1621261055
transform 1 0 1536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_124
timestamp 1621261055
transform 1 0 1152 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_122
timestamp 1621261055
transform 1 0 1152 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_12
timestamp 1621261055
transform 1 0 2304 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_12
timestamp 1621261055
transform 1 0 2304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_20
timestamp 1621261055
transform 1 0 3072 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_20
timestamp 1621261055
transform 1 0 3072 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_29
timestamp 1621261055
transform 1 0 3936 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_28
timestamp 1621261055
transform 1 0 3840 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_198
timestamp 1621261055
transform 1 0 4128 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_825
timestamp 1621261055
transform 1 0 3840 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _126_
timestamp 1621261055
transform 1 0 4320 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_36
timestamp 1621261055
transform 1 0 4608 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_36
timestamp 1621261055
transform 1 0 4608 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_44
timestamp 1621261055
transform 1 0 5376 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_44
timestamp 1621261055
transform 1 0 5376 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_52
timestamp 1621261055
transform 1 0 6144 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_56
timestamp 1621261055
transform 1 0 6528 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_54
timestamp 1621261055
transform 1 0 6336 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_52
timestamp 1621261055
transform 1 0 6144 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_815
timestamp 1621261055
transform 1 0 6432 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_60
timestamp 1621261055
transform 1 0 6912 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_64
timestamp 1621261055
transform 1 0 7296 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_68
timestamp 1621261055
transform 1 0 7680 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_72
timestamp 1621261055
transform 1 0 8064 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_62_82
timestamp 1621261055
transform 1 0 9024 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_80
timestamp 1621261055
transform 1 0 8832 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_76
timestamp 1621261055
transform 1 0 8448 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_80
timestamp 1621261055
transform 1 0 8832 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_826
timestamp 1621261055
transform 1 0 9120 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_92
timestamp 1621261055
transform 1 0 9984 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_84
timestamp 1621261055
transform 1 0 9216 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_88
timestamp 1621261055
transform 1 0 9600 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_96
timestamp 1621261055
transform 1 0 10368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_100
timestamp 1621261055
transform 1 0 10752 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_104
timestamp 1621261055
transform 1 0 11136 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_116
timestamp 1621261055
transform 1 0 12288 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_108
timestamp 1621261055
transform 1 0 11520 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_111
timestamp 1621261055
transform 1 0 11808 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_108
timestamp 1621261055
transform 1 0 11520 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_816
timestamp 1621261055
transform 1 0 11712 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_124
timestamp 1621261055
transform 1 0 13056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_119
timestamp 1621261055
transform 1 0 12576 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_132
timestamp 1621261055
transform 1 0 13824 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_127
timestamp 1621261055
transform 1 0 13344 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_139
timestamp 1621261055
transform 1 0 14496 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_136
timestamp 1621261055
transform 1 0 14208 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_135
timestamp 1621261055
transform 1 0 14112 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_827
timestamp 1621261055
transform 1 0 14400 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_147
timestamp 1621261055
transform 1 0 15264 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_143
timestamp 1621261055
transform 1 0 14880 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_155
timestamp 1621261055
transform 1 0 16032 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_151
timestamp 1621261055
transform 1 0 15648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_163
timestamp 1621261055
transform 1 0 16800 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_163
timestamp 1621261055
transform 1 0 16800 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_159
timestamp 1621261055
transform 1 0 16416 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_817
timestamp 1621261055
transform 1 0 16992 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_171
timestamp 1621261055
transform 1 0 17568 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_173
timestamp 1621261055
transform 1 0 17760 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_166
timestamp 1621261055
transform 1 0 17088 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_122
timestamp 1621261055
transform 1 0 17280 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _169_
timestamp 1621261055
transform 1 0 17472 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_179
timestamp 1621261055
transform 1 0 18336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_181
timestamp 1621261055
transform 1 0 18528 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_191
timestamp 1621261055
transform 1 0 19488 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_187
timestamp 1621261055
transform 1 0 19104 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_189
timestamp 1621261055
transform 1 0 19296 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_194
timestamp 1621261055
transform 1 0 19776 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_197
timestamp 1621261055
transform 1 0 20064 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_828
timestamp 1621261055
transform 1 0 19680 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_202
timestamp 1621261055
transform 1 0 20544 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_205
timestamp 1621261055
transform 1 0 20832 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_210
timestamp 1621261055
transform 1 0 21312 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_213
timestamp 1621261055
transform 1 0 21600 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_218
timestamp 1621261055
transform 1 0 22080 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_221
timestamp 1621261055
transform 1 0 22368 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_219
timestamp 1621261055
transform 1 0 22176 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_217
timestamp 1621261055
transform 1 0 21984 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_818
timestamp 1621261055
transform 1 0 22272 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_226
timestamp 1621261055
transform 1 0 22848 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_229
timestamp 1621261055
transform 1 0 23136 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_234
timestamp 1621261055
transform 1 0 23616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_237
timestamp 1621261055
transform 1 0 23904 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_246
timestamp 1621261055
transform 1 0 24768 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_242
timestamp 1621261055
transform 1 0 24384 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_245
timestamp 1621261055
transform 1 0 24672 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_829
timestamp 1621261055
transform 1 0 24960 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_257
timestamp 1621261055
transform 1 0 25824 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_249
timestamp 1621261055
transform 1 0 25056 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_253
timestamp 1621261055
transform 1 0 25440 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_261
timestamp 1621261055
transform 1 0 26208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_265
timestamp 1621261055
transform 1 0 26592 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_269
timestamp 1621261055
transform 1 0 26976 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_281
timestamp 1621261055
transform 1 0 28128 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_273
timestamp 1621261055
transform 1 0 27360 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_276
timestamp 1621261055
transform 1 0 27648 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_273
timestamp 1621261055
transform 1 0 27360 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_819
timestamp 1621261055
transform 1 0 27552 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_289
timestamp 1621261055
transform 1 0 28896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_284
timestamp 1621261055
transform 1 0 28416 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_297
timestamp 1621261055
transform 1 0 29664 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_292
timestamp 1621261055
transform 1 0 29184 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_304
timestamp 1621261055
transform 1 0 30336 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_301
timestamp 1621261055
transform 1 0 30048 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_61_300
timestamp 1621261055
transform 1 0 29952 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_830
timestamp 1621261055
transform 1 0 30240 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_312
timestamp 1621261055
transform 1 0 31104 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_308
timestamp 1621261055
transform 1 0 30720 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_320
timestamp 1621261055
transform 1 0 31872 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_316
timestamp 1621261055
transform 1 0 31488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_328
timestamp 1621261055
transform 1 0 32640 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_328
timestamp 1621261055
transform 1 0 32640 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_324
timestamp 1621261055
transform 1 0 32256 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_820
timestamp 1621261055
transform 1 0 32832 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_336
timestamp 1621261055
transform 1 0 33408 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_331
timestamp 1621261055
transform 1 0 32928 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_344
timestamp 1621261055
transform 1 0 34176 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_347
timestamp 1621261055
transform 1 0 34464 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_339
timestamp 1621261055
transform 1 0 33696 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_356
timestamp 1621261055
transform 1 0 35328 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_352
timestamp 1621261055
transform 1 0 34944 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_355
timestamp 1621261055
transform 1 0 35232 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_359
timestamp 1621261055
transform 1 0 35616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_363
timestamp 1621261055
transform 1 0 36000 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_831
timestamp 1621261055
transform 1 0 35520 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_367
timestamp 1621261055
transform 1 0 36384 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_371
timestamp 1621261055
transform 1 0 36768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_375
timestamp 1621261055
transform 1 0 37152 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_379
timestamp 1621261055
transform 1 0 37536 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_383
timestamp 1621261055
transform 1 0 37920 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_386
timestamp 1621261055
transform 1 0 38208 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_383
timestamp 1621261055
transform 1 0 37920 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_821
timestamp 1621261055
transform 1 0 38112 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_391
timestamp 1621261055
transform 1 0 38688 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_394
timestamp 1621261055
transform 1 0 38976 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_399
timestamp 1621261055
transform 1 0 39456 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_402
timestamp 1621261055
transform 1 0 39744 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_411
timestamp 1621261055
transform 1 0 40608 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_407
timestamp 1621261055
transform 1 0 40224 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_410
timestamp 1621261055
transform 1 0 40512 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_832
timestamp 1621261055
transform 1 0 40800 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_422
timestamp 1621261055
transform 1 0 41664 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_414
timestamp 1621261055
transform 1 0 40896 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_418
timestamp 1621261055
transform 1 0 41280 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_426
timestamp 1621261055
transform 1 0 42048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_430
timestamp 1621261055
transform 1 0 42432 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_434
timestamp 1621261055
transform 1 0 42816 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_446
timestamp 1621261055
transform 1 0 43968 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_438
timestamp 1621261055
transform 1 0 43200 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_441
timestamp 1621261055
transform 1 0 43488 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_438
timestamp 1621261055
transform 1 0 43200 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_822
timestamp 1621261055
transform 1 0 43392 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_454
timestamp 1621261055
transform 1 0 44736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_449
timestamp 1621261055
transform 1 0 44256 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_462
timestamp 1621261055
transform 1 0 45504 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_61_457
timestamp 1621261055
transform 1 0 45024 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_469
timestamp 1621261055
transform 1 0 46176 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_466
timestamp 1621261055
transform 1 0 45888 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_465
timestamp 1621261055
transform 1 0 45792 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_99
timestamp 1621261055
transform 1 0 46176 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_833
timestamp 1621261055
transform 1 0 46080 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_476
timestamp 1621261055
transform 1 0 46848 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_474
timestamp 1621261055
transform 1 0 46656 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_204
timestamp 1621261055
transform -1 0 46560 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _153_
timestamp 1621261055
transform 1 0 46368 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__conb_1  _133_
timestamp 1621261055
transform -1 0 46848 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_484
timestamp 1621261055
transform 1 0 47616 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_482
timestamp 1621261055
transform 1 0 47424 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_187
timestamp 1621261055
transform -1 0 47808 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _111_
timestamp 1621261055
transform -1 0 48096 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_492
timestamp 1621261055
transform 1 0 48384 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_493
timestamp 1621261055
transform 1 0 48480 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_61_489
timestamp 1621261055
transform 1 0 48096 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_823
timestamp 1621261055
transform 1 0 48672 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_500
timestamp 1621261055
transform 1 0 49152 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_496
timestamp 1621261055
transform 1 0 48768 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_508
timestamp 1621261055
transform 1 0 49920 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_512
timestamp 1621261055
transform 1 0 50304 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_504
timestamp 1621261055
transform 1 0 49536 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_520
timestamp 1621261055
transform 1 0 51072 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_62_516
timestamp 1621261055
transform 1 0 50688 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_157
timestamp 1621261055
transform -1 0 51264 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_62_528
timestamp 1621261055
transform 1 0 51840 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_62_524
timestamp 1621261055
transform 1 0 51456 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_62_522
timestamp 1621261055
transform 1 0 51264 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_525
timestamp 1621261055
transform 1 0 51552 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_834
timestamp 1621261055
transform 1 0 51360 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _082_
timestamp 1621261055
transform -1 0 51552 0 1 43290
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_534
timestamp 1621261055
transform 1 0 52416 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_533
timestamp 1621261055
transform 1 0 52320 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_260
timestamp 1621261055
transform -1 0 52128 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _191_
timestamp 1621261055
transform -1 0 52416 0 -1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_62_542
timestamp 1621261055
transform 1 0 53184 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_541
timestamp 1621261055
transform 1 0 53088 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_550
timestamp 1621261055
transform 1 0 53952 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_551
timestamp 1621261055
transform 1 0 54048 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_61_549
timestamp 1621261055
transform 1 0 53856 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_824
timestamp 1621261055
transform 1 0 53952 0 1 43290
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_62_558
timestamp 1621261055
transform 1 0 54720 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_559
timestamp 1621261055
transform 1 0 54816 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_835
timestamp 1621261055
transform 1 0 56640 0 -1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_61_567
timestamp 1621261055
transform 1 0 55584 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_575
timestamp 1621261055
transform 1 0 56352 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_61_583
timestamp 1621261055
transform 1 0 57120 0 1 43290
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_61_591
timestamp 1621261055
transform 1 0 57888 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_566
timestamp 1621261055
transform 1 0 55488 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_62_574
timestamp 1621261055
transform 1 0 56256 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_62_579
timestamp 1621261055
transform 1 0 56736 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_62_587
timestamp 1621261055
transform 1 0 57504 0 -1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_123
timestamp 1621261055
transform -1 0 58848 0 1 43290
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_125
timestamp 1621261055
transform -1 0 58848 0 -1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_61_595
timestamp 1621261055
transform 1 0 58272 0 1 43290
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_62_595
timestamp 1621261055
transform 1 0 58272 0 -1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_126
timestamp 1621261055
transform 1 0 1152 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_63_4
timestamp 1621261055
transform 1 0 1536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_12
timestamp 1621261055
transform 1 0 2304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_20
timestamp 1621261055
transform 1 0 3072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_28
timestamp 1621261055
transform 1 0 3840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_836
timestamp 1621261055
transform 1 0 6432 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_36
timestamp 1621261055
transform 1 0 4608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_44
timestamp 1621261055
transform 1 0 5376 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_52
timestamp 1621261055
transform 1 0 6144 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_54
timestamp 1621261055
transform 1 0 6336 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_56
timestamp 1621261055
transform 1 0 6528 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_64
timestamp 1621261055
transform 1 0 7296 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_72
timestamp 1621261055
transform 1 0 8064 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_80
timestamp 1621261055
transform 1 0 8832 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_88
timestamp 1621261055
transform 1 0 9600 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_96
timestamp 1621261055
transform 1 0 10368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _097_
timestamp 1621261055
transform 1 0 12192 0 1 44622
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_837
timestamp 1621261055
transform 1 0 11712 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_175
timestamp 1621261055
transform 1 0 12000 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_63_104
timestamp 1621261055
transform 1 0 11136 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_108
timestamp 1621261055
transform 1 0 11520 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_111
timestamp 1621261055
transform 1 0 11808 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_118
timestamp 1621261055
transform 1 0 12480 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_126
timestamp 1621261055
transform 1 0 13248 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_838
timestamp 1621261055
transform 1 0 16992 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_134
timestamp 1621261055
transform 1 0 14016 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_142
timestamp 1621261055
transform 1 0 14784 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_150
timestamp 1621261055
transform 1 0 15552 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_158
timestamp 1621261055
transform 1 0 16320 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_162
timestamp 1621261055
transform 1 0 16704 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_63_164
timestamp 1621261055
transform 1 0 16896 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_166
timestamp 1621261055
transform 1 0 17088 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_174
timestamp 1621261055
transform 1 0 17856 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_182
timestamp 1621261055
transform 1 0 18624 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_190
timestamp 1621261055
transform 1 0 19392 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_198
timestamp 1621261055
transform 1 0 20160 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_839
timestamp 1621261055
transform 1 0 22272 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_206
timestamp 1621261055
transform 1 0 20928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_214
timestamp 1621261055
transform 1 0 21696 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_218
timestamp 1621261055
transform 1 0 22080 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_221
timestamp 1621261055
transform 1 0 22368 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_229
timestamp 1621261055
transform 1 0 23136 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_237
timestamp 1621261055
transform 1 0 23904 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_245
timestamp 1621261055
transform 1 0 24672 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_253
timestamp 1621261055
transform 1 0 25440 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_261
timestamp 1621261055
transform 1 0 26208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_840
timestamp 1621261055
transform 1 0 27552 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_269
timestamp 1621261055
transform 1 0 26976 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_273
timestamp 1621261055
transform 1 0 27360 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_276
timestamp 1621261055
transform 1 0 27648 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_284
timestamp 1621261055
transform 1 0 28416 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_292
timestamp 1621261055
transform 1 0 29184 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_841
timestamp 1621261055
transform 1 0 32832 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_300
timestamp 1621261055
transform 1 0 29952 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_308
timestamp 1621261055
transform 1 0 30720 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_316
timestamp 1621261055
transform 1 0 31488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_324
timestamp 1621261055
transform 1 0 32256 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_328
timestamp 1621261055
transform 1 0 32640 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_331
timestamp 1621261055
transform 1 0 32928 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_339
timestamp 1621261055
transform 1 0 33696 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_347
timestamp 1621261055
transform 1 0 34464 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_355
timestamp 1621261055
transform 1 0 35232 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_363
timestamp 1621261055
transform 1 0 36000 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_842
timestamp 1621261055
transform 1 0 38112 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_371
timestamp 1621261055
transform 1 0 36768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_379
timestamp 1621261055
transform 1 0 37536 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_383
timestamp 1621261055
transform 1 0 37920 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_386
timestamp 1621261055
transform 1 0 38208 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_394
timestamp 1621261055
transform 1 0 38976 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_402
timestamp 1621261055
transform 1 0 39744 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_410
timestamp 1621261055
transform 1 0 40512 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_418
timestamp 1621261055
transform 1 0 41280 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_426
timestamp 1621261055
transform 1 0 42048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_843
timestamp 1621261055
transform 1 0 43392 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_63_434
timestamp 1621261055
transform 1 0 42816 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_438
timestamp 1621261055
transform 1 0 43200 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_441
timestamp 1621261055
transform 1 0 43488 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_449
timestamp 1621261055
transform 1 0 44256 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_457
timestamp 1621261055
transform 1 0 45024 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_844
timestamp 1621261055
transform 1 0 48672 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_465
timestamp 1621261055
transform 1 0 45792 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_473
timestamp 1621261055
transform 1 0 46560 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_481
timestamp 1621261055
transform 1 0 47328 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_489
timestamp 1621261055
transform 1 0 48096 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_493
timestamp 1621261055
transform 1 0 48480 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_496
timestamp 1621261055
transform 1 0 48768 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_504
timestamp 1621261055
transform 1 0 49536 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_512
timestamp 1621261055
transform 1 0 50304 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_520
timestamp 1621261055
transform 1 0 51072 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_528
timestamp 1621261055
transform 1 0 51840 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_845
timestamp 1621261055
transform 1 0 53952 0 1 44622
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_63_536
timestamp 1621261055
transform 1 0 52608 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_544
timestamp 1621261055
transform 1 0 53376 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_548
timestamp 1621261055
transform 1 0 53760 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_63_551
timestamp 1621261055
transform 1 0 54048 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_559
timestamp 1621261055
transform 1 0 54816 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_567
timestamp 1621261055
transform 1 0 55584 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_575
timestamp 1621261055
transform 1 0 56352 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_63_583
timestamp 1621261055
transform 1 0 57120 0 1 44622
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_63_591
timestamp 1621261055
transform 1 0 57888 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_127
timestamp 1621261055
transform -1 0 58848 0 1 44622
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_63_595
timestamp 1621261055
transform 1 0 58272 0 1 44622
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_128
timestamp 1621261055
transform 1 0 1152 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_846
timestamp 1621261055
transform 1 0 3840 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_4
timestamp 1621261055
transform 1 0 1536 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_12
timestamp 1621261055
transform 1 0 2304 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_20
timestamp 1621261055
transform 1 0 3072 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_29
timestamp 1621261055
transform 1 0 3936 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_37
timestamp 1621261055
transform 1 0 4704 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_45
timestamp 1621261055
transform 1 0 5472 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_53
timestamp 1621261055
transform 1 0 6240 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_61
timestamp 1621261055
transform 1 0 7008 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_847
timestamp 1621261055
transform 1 0 9120 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_69
timestamp 1621261055
transform 1 0 7776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_77
timestamp 1621261055
transform 1 0 8544 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_81
timestamp 1621261055
transform 1 0 8928 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_84
timestamp 1621261055
transform 1 0 9216 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_92
timestamp 1621261055
transform 1 0 9984 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _205_
timestamp 1621261055
transform -1 0 12864 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_244
timestamp 1621261055
transform -1 0 12576 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_100
timestamp 1621261055
transform 1 0 10752 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_108
timestamp 1621261055
transform 1 0 11520 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_64_116
timestamp 1621261055
transform 1 0 12288 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_122
timestamp 1621261055
transform 1 0 12864 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_130
timestamp 1621261055
transform 1 0 13632 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_848
timestamp 1621261055
transform 1 0 14400 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_139
timestamp 1621261055
transform 1 0 14496 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_147
timestamp 1621261055
transform 1 0 15264 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_155
timestamp 1621261055
transform 1 0 16032 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_163
timestamp 1621261055
transform 1 0 16800 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_849
timestamp 1621261055
transform 1 0 19680 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_171
timestamp 1621261055
transform 1 0 17568 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_179
timestamp 1621261055
transform 1 0 18336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_187
timestamp 1621261055
transform 1 0 19104 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_191
timestamp 1621261055
transform 1 0 19488 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_194
timestamp 1621261055
transform 1 0 19776 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_202
timestamp 1621261055
transform 1 0 20544 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_210
timestamp 1621261055
transform 1 0 21312 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_218
timestamp 1621261055
transform 1 0 22080 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_226
timestamp 1621261055
transform 1 0 22848 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_850
timestamp 1621261055
transform 1 0 24960 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_234
timestamp 1621261055
transform 1 0 23616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_242
timestamp 1621261055
transform 1 0 24384 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_246
timestamp 1621261055
transform 1 0 24768 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_249
timestamp 1621261055
transform 1 0 25056 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_257
timestamp 1621261055
transform 1 0 25824 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_265
timestamp 1621261055
transform 1 0 26592 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_273
timestamp 1621261055
transform 1 0 27360 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_281
timestamp 1621261055
transform 1 0 28128 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_289
timestamp 1621261055
transform 1 0 28896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_297
timestamp 1621261055
transform 1 0 29664 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_851
timestamp 1621261055
transform 1 0 30240 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_301
timestamp 1621261055
transform 1 0 30048 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_304
timestamp 1621261055
transform 1 0 30336 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_312
timestamp 1621261055
transform 1 0 31104 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_320
timestamp 1621261055
transform 1 0 31872 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_328
timestamp 1621261055
transform 1 0 32640 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_852
timestamp 1621261055
transform 1 0 35520 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_336
timestamp 1621261055
transform 1 0 33408 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_344
timestamp 1621261055
transform 1 0 34176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_352
timestamp 1621261055
transform 1 0 34944 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_356
timestamp 1621261055
transform 1 0 35328 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_359
timestamp 1621261055
transform 1 0 35616 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_367
timestamp 1621261055
transform 1 0 36384 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_375
timestamp 1621261055
transform 1 0 37152 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_383
timestamp 1621261055
transform 1 0 37920 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_391
timestamp 1621261055
transform 1 0 38688 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_853
timestamp 1621261055
transform 1 0 40800 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_64_399
timestamp 1621261055
transform 1 0 39456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_407
timestamp 1621261055
transform 1 0 40224 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_411
timestamp 1621261055
transform 1 0 40608 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_414
timestamp 1621261055
transform 1 0 40896 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_422
timestamp 1621261055
transform 1 0 41664 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_430
timestamp 1621261055
transform 1 0 42432 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_438
timestamp 1621261055
transform 1 0 43200 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_446
timestamp 1621261055
transform 1 0 43968 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_454
timestamp 1621261055
transform 1 0 44736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_462
timestamp 1621261055
transform 1 0 45504 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _038_
timestamp 1621261055
transform 1 0 47808 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_854
timestamp 1621261055
transform 1 0 46080 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_466
timestamp 1621261055
transform 1 0 45888 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_469
timestamp 1621261055
transform 1 0 46176 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_477
timestamp 1621261055
transform 1 0 46944 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_64_485
timestamp 1621261055
transform 1 0 47712 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_489
timestamp 1621261055
transform 1 0 48096 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_493
timestamp 1621261055
transform 1 0 48480 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_64_495
timestamp 1621261055
transform 1 0 48672 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _100_
timestamp 1621261055
transform -1 0 49248 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_855
timestamp 1621261055
transform 1 0 51360 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_179
timestamp 1621261055
transform -1 0 48960 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_501
timestamp 1621261055
transform 1 0 49248 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_509
timestamp 1621261055
transform 1 0 50016 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_64_517
timestamp 1621261055
transform 1 0 50784 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_521
timestamp 1621261055
transform 1 0 51168 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_64_524
timestamp 1621261055
transform 1 0 51456 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_532
timestamp 1621261055
transform 1 0 52224 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_540
timestamp 1621261055
transform 1 0 52992 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_548
timestamp 1621261055
transform 1 0 53760 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_556
timestamp 1621261055
transform 1 0 54528 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _168_
timestamp 1621261055
transform -1 0 56256 0 -1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_856
timestamp 1621261055
transform 1 0 56640 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_120
timestamp 1621261055
transform -1 0 55968 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_64_564
timestamp 1621261055
transform 1 0 55296 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_64_568
timestamp 1621261055
transform 1 0 55680 0 -1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_64_574
timestamp 1621261055
transform 1 0 56256 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_64_579
timestamp 1621261055
transform 1 0 56736 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_64_587
timestamp 1621261055
transform 1 0 57504 0 -1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_129
timestamp 1621261055
transform -1 0 58848 0 -1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_64_595
timestamp 1621261055
transform 1 0 58272 0 -1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_130
timestamp 1621261055
transform 1 0 1152 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_4
timestamp 1621261055
transform 1 0 1536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_12
timestamp 1621261055
transform 1 0 2304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_20
timestamp 1621261055
transform 1 0 3072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_28
timestamp 1621261055
transform 1 0 3840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_857
timestamp 1621261055
transform 1 0 6432 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_36
timestamp 1621261055
transform 1 0 4608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_44
timestamp 1621261055
transform 1 0 5376 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_52
timestamp 1621261055
transform 1 0 6144 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_65_54
timestamp 1621261055
transform 1 0 6336 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_56
timestamp 1621261055
transform 1 0 6528 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_64
timestamp 1621261055
transform 1 0 7296 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_72
timestamp 1621261055
transform 1 0 8064 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_80
timestamp 1621261055
transform 1 0 8832 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_88
timestamp 1621261055
transform 1 0 9600 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_96
timestamp 1621261055
transform 1 0 10368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_858
timestamp 1621261055
transform 1 0 11712 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_104
timestamp 1621261055
transform 1 0 11136 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_108
timestamp 1621261055
transform 1 0 11520 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_111
timestamp 1621261055
transform 1 0 11808 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_119
timestamp 1621261055
transform 1 0 12576 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_127
timestamp 1621261055
transform 1 0 13344 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_859
timestamp 1621261055
transform 1 0 16992 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_135
timestamp 1621261055
transform 1 0 14112 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_143
timestamp 1621261055
transform 1 0 14880 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_151
timestamp 1621261055
transform 1 0 15648 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_159
timestamp 1621261055
transform 1 0 16416 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_163
timestamp 1621261055
transform 1 0 16800 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _165_
timestamp 1621261055
transform 1 0 17760 0 1 45954
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_114
timestamp 1621261055
transform 1 0 17568 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_65_166
timestamp 1621261055
transform 1 0 17088 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_65_170
timestamp 1621261055
transform 1 0 17472 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_176
timestamp 1621261055
transform 1 0 18048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_184
timestamp 1621261055
transform 1 0 18816 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_192
timestamp 1621261055
transform 1 0 19584 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_860
timestamp 1621261055
transform 1 0 22272 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_200
timestamp 1621261055
transform 1 0 20352 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_208
timestamp 1621261055
transform 1 0 21120 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_216
timestamp 1621261055
transform 1 0 21888 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_65_221
timestamp 1621261055
transform 1 0 22368 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_229
timestamp 1621261055
transform 1 0 23136 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_237
timestamp 1621261055
transform 1 0 23904 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_245
timestamp 1621261055
transform 1 0 24672 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_253
timestamp 1621261055
transform 1 0 25440 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_261
timestamp 1621261055
transform 1 0 26208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_861
timestamp 1621261055
transform 1 0 27552 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_269
timestamp 1621261055
transform 1 0 26976 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_273
timestamp 1621261055
transform 1 0 27360 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_276
timestamp 1621261055
transform 1 0 27648 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_284
timestamp 1621261055
transform 1 0 28416 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_292
timestamp 1621261055
transform 1 0 29184 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_862
timestamp 1621261055
transform 1 0 32832 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_300
timestamp 1621261055
transform 1 0 29952 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_308
timestamp 1621261055
transform 1 0 30720 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_316
timestamp 1621261055
transform 1 0 31488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_324
timestamp 1621261055
transform 1 0 32256 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_328
timestamp 1621261055
transform 1 0 32640 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_331
timestamp 1621261055
transform 1 0 32928 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_339
timestamp 1621261055
transform 1 0 33696 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_347
timestamp 1621261055
transform 1 0 34464 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_355
timestamp 1621261055
transform 1 0 35232 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_363
timestamp 1621261055
transform 1 0 36000 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_863
timestamp 1621261055
transform 1 0 38112 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_371
timestamp 1621261055
transform 1 0 36768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_379
timestamp 1621261055
transform 1 0 37536 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_383
timestamp 1621261055
transform 1 0 37920 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_386
timestamp 1621261055
transform 1 0 38208 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_394
timestamp 1621261055
transform 1 0 38976 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_402
timestamp 1621261055
transform 1 0 39744 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_410
timestamp 1621261055
transform 1 0 40512 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_418
timestamp 1621261055
transform 1 0 41280 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_426
timestamp 1621261055
transform 1 0 42048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_864
timestamp 1621261055
transform 1 0 43392 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_65_434
timestamp 1621261055
transform 1 0 42816 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_438
timestamp 1621261055
transform 1 0 43200 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_441
timestamp 1621261055
transform 1 0 43488 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_449
timestamp 1621261055
transform 1 0 44256 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_457
timestamp 1621261055
transform 1 0 45024 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_865
timestamp 1621261055
transform 1 0 48672 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_465
timestamp 1621261055
transform 1 0 45792 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_473
timestamp 1621261055
transform 1 0 46560 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_481
timestamp 1621261055
transform 1 0 47328 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_489
timestamp 1621261055
transform 1 0 48096 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_493
timestamp 1621261055
transform 1 0 48480 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_496
timestamp 1621261055
transform 1 0 48768 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_504
timestamp 1621261055
transform 1 0 49536 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_512
timestamp 1621261055
transform 1 0 50304 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_520
timestamp 1621261055
transform 1 0 51072 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_528
timestamp 1621261055
transform 1 0 51840 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_866
timestamp 1621261055
transform 1 0 53952 0 1 45954
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_65_536
timestamp 1621261055
transform 1 0 52608 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_544
timestamp 1621261055
transform 1 0 53376 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_548
timestamp 1621261055
transform 1 0 53760 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_65_551
timestamp 1621261055
transform 1 0 54048 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_559
timestamp 1621261055
transform 1 0 54816 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_567
timestamp 1621261055
transform 1 0 55584 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_575
timestamp 1621261055
transform 1 0 56352 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_65_583
timestamp 1621261055
transform 1 0 57120 0 1 45954
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_65_591
timestamp 1621261055
transform 1 0 57888 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_131
timestamp 1621261055
transform -1 0 58848 0 1 45954
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_65_595
timestamp 1621261055
transform 1 0 58272 0 1 45954
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_132
timestamp 1621261055
transform 1 0 1152 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_867
timestamp 1621261055
transform 1 0 3840 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_4
timestamp 1621261055
transform 1 0 1536 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_12
timestamp 1621261055
transform 1 0 2304 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_20
timestamp 1621261055
transform 1 0 3072 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_29
timestamp 1621261055
transform 1 0 3936 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_37
timestamp 1621261055
transform 1 0 4704 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_45
timestamp 1621261055
transform 1 0 5472 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_53
timestamp 1621261055
transform 1 0 6240 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_61
timestamp 1621261055
transform 1 0 7008 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_868
timestamp 1621261055
transform 1 0 9120 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_69
timestamp 1621261055
transform 1 0 7776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_77
timestamp 1621261055
transform 1 0 8544 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_81
timestamp 1621261055
transform 1 0 8928 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_84
timestamp 1621261055
transform 1 0 9216 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_92
timestamp 1621261055
transform 1 0 9984 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_100
timestamp 1621261055
transform 1 0 10752 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_108
timestamp 1621261055
transform 1 0 11520 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_116
timestamp 1621261055
transform 1 0 12288 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_124
timestamp 1621261055
transform 1 0 13056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_132
timestamp 1621261055
transform 1 0 13824 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_869
timestamp 1621261055
transform 1 0 14400 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_136
timestamp 1621261055
transform 1 0 14208 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_139
timestamp 1621261055
transform 1 0 14496 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_147
timestamp 1621261055
transform 1 0 15264 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_155
timestamp 1621261055
transform 1 0 16032 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_163
timestamp 1621261055
transform 1 0 16800 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_870
timestamp 1621261055
transform 1 0 19680 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_171
timestamp 1621261055
transform 1 0 17568 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_179
timestamp 1621261055
transform 1 0 18336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_187
timestamp 1621261055
transform 1 0 19104 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_191
timestamp 1621261055
transform 1 0 19488 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_194
timestamp 1621261055
transform 1 0 19776 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_202
timestamp 1621261055
transform 1 0 20544 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_210
timestamp 1621261055
transform 1 0 21312 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_218
timestamp 1621261055
transform 1 0 22080 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_226
timestamp 1621261055
transform 1 0 22848 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_871
timestamp 1621261055
transform 1 0 24960 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_234
timestamp 1621261055
transform 1 0 23616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_242
timestamp 1621261055
transform 1 0 24384 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_246
timestamp 1621261055
transform 1 0 24768 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_249
timestamp 1621261055
transform 1 0 25056 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_257
timestamp 1621261055
transform 1 0 25824 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_265
timestamp 1621261055
transform 1 0 26592 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_273
timestamp 1621261055
transform 1 0 27360 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_281
timestamp 1621261055
transform 1 0 28128 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_289
timestamp 1621261055
transform 1 0 28896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_297
timestamp 1621261055
transform 1 0 29664 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_872
timestamp 1621261055
transform 1 0 30240 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_301
timestamp 1621261055
transform 1 0 30048 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_304
timestamp 1621261055
transform 1 0 30336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_312
timestamp 1621261055
transform 1 0 31104 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_320
timestamp 1621261055
transform 1 0 31872 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_328
timestamp 1621261055
transform 1 0 32640 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_873
timestamp 1621261055
transform 1 0 35520 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_336
timestamp 1621261055
transform 1 0 33408 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_344
timestamp 1621261055
transform 1 0 34176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_352
timestamp 1621261055
transform 1 0 34944 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_356
timestamp 1621261055
transform 1 0 35328 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_359
timestamp 1621261055
transform 1 0 35616 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _120_
timestamp 1621261055
transform 1 0 36576 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_192
timestamp 1621261055
transform 1 0 36384 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_372
timestamp 1621261055
transform 1 0 36864 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_380
timestamp 1621261055
transform 1 0 37632 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_388
timestamp 1621261055
transform 1 0 38400 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_396
timestamp 1621261055
transform 1 0 39168 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_874
timestamp 1621261055
transform 1 0 40800 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_404
timestamp 1621261055
transform 1 0 39936 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_66_412
timestamp 1621261055
transform 1 0 40704 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_414
timestamp 1621261055
transform 1 0 40896 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_422
timestamp 1621261055
transform 1 0 41664 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_430
timestamp 1621261055
transform 1 0 42432 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_438
timestamp 1621261055
transform 1 0 43200 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_446
timestamp 1621261055
transform 1 0 43968 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_454
timestamp 1621261055
transform 1 0 44736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_462
timestamp 1621261055
transform 1 0 45504 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_875
timestamp 1621261055
transform 1 0 46080 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_466
timestamp 1621261055
transform 1 0 45888 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_469
timestamp 1621261055
transform 1 0 46176 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_477
timestamp 1621261055
transform 1 0 46944 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_485
timestamp 1621261055
transform 1 0 47712 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_493
timestamp 1621261055
transform 1 0 48480 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_876
timestamp 1621261055
transform 1 0 51360 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_501
timestamp 1621261055
transform 1 0 49248 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_509
timestamp 1621261055
transform 1 0 50016 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_66_517
timestamp 1621261055
transform 1 0 50784 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_521
timestamp 1621261055
transform 1 0 51168 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_66_524
timestamp 1621261055
transform 1 0 51456 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _032_
timestamp 1621261055
transform 1 0 52512 0 -1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_532
timestamp 1621261055
transform 1 0 52224 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_66_534
timestamp 1621261055
transform 1 0 52416 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_538
timestamp 1621261055
transform 1 0 52800 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_546
timestamp 1621261055
transform 1 0 53568 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_554
timestamp 1621261055
transform 1 0 54336 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_877
timestamp 1621261055
transform 1 0 56640 0 -1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_66_562
timestamp 1621261055
transform 1 0 55104 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_570
timestamp 1621261055
transform 1 0 55872 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_579
timestamp 1621261055
transform 1 0 56736 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_66_587
timestamp 1621261055
transform 1 0 57504 0 -1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_133
timestamp 1621261055
transform -1 0 58848 0 -1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_66_595
timestamp 1621261055
transform 1 0 58272 0 -1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_134
timestamp 1621261055
transform 1 0 1152 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_4
timestamp 1621261055
transform 1 0 1536 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_12
timestamp 1621261055
transform 1 0 2304 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_20
timestamp 1621261055
transform 1 0 3072 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_28
timestamp 1621261055
transform 1 0 3840 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_878
timestamp 1621261055
transform 1 0 6432 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_36
timestamp 1621261055
transform 1 0 4608 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_44
timestamp 1621261055
transform 1 0 5376 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_52
timestamp 1621261055
transform 1 0 6144 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_54
timestamp 1621261055
transform 1 0 6336 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_56
timestamp 1621261055
transform 1 0 6528 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_64
timestamp 1621261055
transform 1 0 7296 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _093_
timestamp 1621261055
transform 1 0 8160 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_169
timestamp 1621261055
transform 1 0 7968 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_68
timestamp 1621261055
transform 1 0 7680 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_70
timestamp 1621261055
transform 1 0 7872 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_76
timestamp 1621261055
transform 1 0 8448 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_84
timestamp 1621261055
transform 1 0 9216 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_92
timestamp 1621261055
transform 1 0 9984 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_879
timestamp 1621261055
transform 1 0 11712 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_100
timestamp 1621261055
transform 1 0 10752 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_108
timestamp 1621261055
transform 1 0 11520 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_111
timestamp 1621261055
transform 1 0 11808 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_119
timestamp 1621261055
transform 1 0 12576 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_127
timestamp 1621261055
transform 1 0 13344 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_880
timestamp 1621261055
transform 1 0 16992 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_135
timestamp 1621261055
transform 1 0 14112 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_143
timestamp 1621261055
transform 1 0 14880 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_151
timestamp 1621261055
transform 1 0 15648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_159
timestamp 1621261055
transform 1 0 16416 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_163
timestamp 1621261055
transform 1 0 16800 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_166
timestamp 1621261055
transform 1 0 17088 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_174
timestamp 1621261055
transform 1 0 17856 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_182
timestamp 1621261055
transform 1 0 18624 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_190
timestamp 1621261055
transform 1 0 19392 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_198
timestamp 1621261055
transform 1 0 20160 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_881
timestamp 1621261055
transform 1 0 22272 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_206
timestamp 1621261055
transform 1 0 20928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_214
timestamp 1621261055
transform 1 0 21696 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_218
timestamp 1621261055
transform 1 0 22080 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_221
timestamp 1621261055
transform 1 0 22368 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_229
timestamp 1621261055
transform 1 0 23136 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_237
timestamp 1621261055
transform 1 0 23904 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_245
timestamp 1621261055
transform 1 0 24672 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_253
timestamp 1621261055
transform 1 0 25440 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_261
timestamp 1621261055
transform 1 0 26208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_882
timestamp 1621261055
transform 1 0 27552 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_269
timestamp 1621261055
transform 1 0 26976 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_273
timestamp 1621261055
transform 1 0 27360 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_276
timestamp 1621261055
transform 1 0 27648 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_284
timestamp 1621261055
transform 1 0 28416 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_292
timestamp 1621261055
transform 1 0 29184 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_883
timestamp 1621261055
transform 1 0 32832 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_300
timestamp 1621261055
transform 1 0 29952 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_308
timestamp 1621261055
transform 1 0 30720 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_316
timestamp 1621261055
transform 1 0 31488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_324
timestamp 1621261055
transform 1 0 32256 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_328
timestamp 1621261055
transform 1 0 32640 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_331
timestamp 1621261055
transform 1 0 32928 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_339
timestamp 1621261055
transform 1 0 33696 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_347
timestamp 1621261055
transform 1 0 34464 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_355
timestamp 1621261055
transform 1 0 35232 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_363
timestamp 1621261055
transform 1 0 36000 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_884
timestamp 1621261055
transform 1 0 38112 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_371
timestamp 1621261055
transform 1 0 36768 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_379
timestamp 1621261055
transform 1 0 37536 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_383
timestamp 1621261055
transform 1 0 37920 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_386
timestamp 1621261055
transform 1 0 38208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_394
timestamp 1621261055
transform 1 0 38976 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_402
timestamp 1621261055
transform 1 0 39744 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_410
timestamp 1621261055
transform 1 0 40512 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_418
timestamp 1621261055
transform 1 0 41280 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_426
timestamp 1621261055
transform 1 0 42048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_885
timestamp 1621261055
transform 1 0 43392 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_67_434
timestamp 1621261055
transform 1 0 42816 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_438
timestamp 1621261055
transform 1 0 43200 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_67_441
timestamp 1621261055
transform 1 0 43488 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_449
timestamp 1621261055
transform 1 0 44256 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_457
timestamp 1621261055
transform 1 0 45024 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_886
timestamp 1621261055
transform 1 0 48672 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_465
timestamp 1621261055
transform 1 0 45792 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_473
timestamp 1621261055
transform 1 0 46560 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_481
timestamp 1621261055
transform 1 0 47328 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_489
timestamp 1621261055
transform 1 0 48096 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_493
timestamp 1621261055
transform 1 0 48480 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _011_
timestamp 1621261055
transform 1 0 49152 0 1 47286
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_67_496
timestamp 1621261055
transform 1 0 48768 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_67_503
timestamp 1621261055
transform 1 0 49440 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_511
timestamp 1621261055
transform 1 0 50208 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_519
timestamp 1621261055
transform 1 0 50976 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_527
timestamp 1621261055
transform 1 0 51744 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_887
timestamp 1621261055
transform 1 0 53952 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_535
timestamp 1621261055
transform 1 0 52512 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_543
timestamp 1621261055
transform 1 0 53280 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_547
timestamp 1621261055
transform 1 0 53664 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_67_549
timestamp 1621261055
transform 1 0 53856 0 1 47286
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_67_551
timestamp 1621261055
transform 1 0 54048 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_559
timestamp 1621261055
transform 1 0 54816 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_567
timestamp 1621261055
transform 1 0 55584 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_575
timestamp 1621261055
transform 1 0 56352 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_67_583
timestamp 1621261055
transform 1 0 57120 0 1 47286
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_67_591
timestamp 1621261055
transform 1 0 57888 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_135
timestamp 1621261055
transform -1 0 58848 0 1 47286
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_67_595
timestamp 1621261055
transform 1 0 58272 0 1 47286
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _172_
timestamp 1621261055
transform 1 0 2496 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  PHY_136
timestamp 1621261055
transform 1 0 1152 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_888
timestamp 1621261055
transform 1 0 3840 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_127
timestamp 1621261055
transform 1 0 2304 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_4
timestamp 1621261055
transform 1 0 1536 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_17
timestamp 1621261055
transform 1 0 2784 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_25
timestamp 1621261055
transform 1 0 3552 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_68_27
timestamp 1621261055
transform 1 0 3744 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_29
timestamp 1621261055
transform 1 0 3936 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_37
timestamp 1621261055
transform 1 0 4704 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_45
timestamp 1621261055
transform 1 0 5472 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_53
timestamp 1621261055
transform 1 0 6240 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_61
timestamp 1621261055
transform 1 0 7008 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_889
timestamp 1621261055
transform 1 0 9120 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_69
timestamp 1621261055
transform 1 0 7776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_77
timestamp 1621261055
transform 1 0 8544 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_81
timestamp 1621261055
transform 1 0 8928 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_84
timestamp 1621261055
transform 1 0 9216 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_92
timestamp 1621261055
transform 1 0 9984 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_100
timestamp 1621261055
transform 1 0 10752 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_108
timestamp 1621261055
transform 1 0 11520 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_116
timestamp 1621261055
transform 1 0 12288 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_124
timestamp 1621261055
transform 1 0 13056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_132
timestamp 1621261055
transform 1 0 13824 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_890
timestamp 1621261055
transform 1 0 14400 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_136
timestamp 1621261055
transform 1 0 14208 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_139
timestamp 1621261055
transform 1 0 14496 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_147
timestamp 1621261055
transform 1 0 15264 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_155
timestamp 1621261055
transform 1 0 16032 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_163
timestamp 1621261055
transform 1 0 16800 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_891
timestamp 1621261055
transform 1 0 19680 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_171
timestamp 1621261055
transform 1 0 17568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_179
timestamp 1621261055
transform 1 0 18336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_187
timestamp 1621261055
transform 1 0 19104 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_191
timestamp 1621261055
transform 1 0 19488 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_194
timestamp 1621261055
transform 1 0 19776 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_202
timestamp 1621261055
transform 1 0 20544 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_210
timestamp 1621261055
transform 1 0 21312 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_218
timestamp 1621261055
transform 1 0 22080 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_226
timestamp 1621261055
transform 1 0 22848 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_892
timestamp 1621261055
transform 1 0 24960 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_234
timestamp 1621261055
transform 1 0 23616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_242
timestamp 1621261055
transform 1 0 24384 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_246
timestamp 1621261055
transform 1 0 24768 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_249
timestamp 1621261055
transform 1 0 25056 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_257
timestamp 1621261055
transform 1 0 25824 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_265
timestamp 1621261055
transform 1 0 26592 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_273
timestamp 1621261055
transform 1 0 27360 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_281
timestamp 1621261055
transform 1 0 28128 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_289
timestamp 1621261055
transform 1 0 28896 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_297
timestamp 1621261055
transform 1 0 29664 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_893
timestamp 1621261055
transform 1 0 30240 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_301
timestamp 1621261055
transform 1 0 30048 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_304
timestamp 1621261055
transform 1 0 30336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_312
timestamp 1621261055
transform 1 0 31104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_320
timestamp 1621261055
transform 1 0 31872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_328
timestamp 1621261055
transform 1 0 32640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_894
timestamp 1621261055
transform 1 0 35520 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_336
timestamp 1621261055
transform 1 0 33408 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_344
timestamp 1621261055
transform 1 0 34176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_352
timestamp 1621261055
transform 1 0 34944 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_356
timestamp 1621261055
transform 1 0 35328 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_359
timestamp 1621261055
transform 1 0 35616 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_367
timestamp 1621261055
transform 1 0 36384 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_375
timestamp 1621261055
transform 1 0 37152 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_383
timestamp 1621261055
transform 1 0 37920 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_391
timestamp 1621261055
transform 1 0 38688 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _118_
timestamp 1621261055
transform -1 0 41568 0 -1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_895
timestamp 1621261055
transform 1 0 40800 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_190
timestamp 1621261055
transform -1 0 41280 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_399
timestamp 1621261055
transform 1 0 39456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_407
timestamp 1621261055
transform 1 0 40224 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_411
timestamp 1621261055
transform 1 0 40608 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_414
timestamp 1621261055
transform 1 0 40896 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_421
timestamp 1621261055
transform 1 0 41568 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_429
timestamp 1621261055
transform 1 0 42336 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_437
timestamp 1621261055
transform 1 0 43104 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_445
timestamp 1621261055
transform 1 0 43872 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_453
timestamp 1621261055
transform 1 0 44640 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_461
timestamp 1621261055
transform 1 0 45408 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_896
timestamp 1621261055
transform 1 0 46080 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_465
timestamp 1621261055
transform 1 0 45792 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_68_467
timestamp 1621261055
transform 1 0 45984 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_469
timestamp 1621261055
transform 1 0 46176 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_477
timestamp 1621261055
transform 1 0 46944 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_485
timestamp 1621261055
transform 1 0 47712 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_493
timestamp 1621261055
transform 1 0 48480 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_897
timestamp 1621261055
transform 1 0 51360 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_501
timestamp 1621261055
transform 1 0 49248 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_509
timestamp 1621261055
transform 1 0 50016 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_517
timestamp 1621261055
transform 1 0 50784 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_521
timestamp 1621261055
transform 1 0 51168 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_524
timestamp 1621261055
transform 1 0 51456 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_532
timestamp 1621261055
transform 1 0 52224 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_540
timestamp 1621261055
transform 1 0 52992 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_548
timestamp 1621261055
transform 1 0 53760 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_556
timestamp 1621261055
transform 1 0 54528 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_898
timestamp 1621261055
transform 1 0 56640 0 -1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_68_564
timestamp 1621261055
transform 1 0 55296 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_68_572
timestamp 1621261055
transform 1 0 56064 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_576
timestamp 1621261055
transform 1 0 56448 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_68_579
timestamp 1621261055
transform 1 0 56736 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_68_587
timestamp 1621261055
transform 1 0 57504 0 -1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_137
timestamp 1621261055
transform -1 0 58848 0 -1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_68_595
timestamp 1621261055
transform 1 0 58272 0 -1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_4
timestamp 1621261055
transform 1 0 1536 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_4
timestamp 1621261055
transform 1 0 1536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_140
timestamp 1621261055
transform 1 0 1152 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_138
timestamp 1621261055
transform 1 0 1152 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_12
timestamp 1621261055
transform 1 0 2304 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_12
timestamp 1621261055
transform 1 0 2304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_20
timestamp 1621261055
transform 1 0 3072 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_20
timestamp 1621261055
transform 1 0 3072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_29
timestamp 1621261055
transform 1 0 3936 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_28
timestamp 1621261055
transform 1 0 3840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_219
timestamp 1621261055
transform 1 0 4128 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_909
timestamp 1621261055
transform 1 0 3840 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _146_
timestamp 1621261055
transform 1 0 4320 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_36
timestamp 1621261055
transform 1 0 4608 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_36
timestamp 1621261055
transform 1 0 4608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_44
timestamp 1621261055
transform 1 0 5376 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_44
timestamp 1621261055
transform 1 0 5376 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_52
timestamp 1621261055
transform 1 0 6144 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_56
timestamp 1621261055
transform 1 0 6528 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_69_54
timestamp 1621261055
transform 1 0 6336 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_52
timestamp 1621261055
transform 1 0 6144 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_899
timestamp 1621261055
transform 1 0 6432 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_60
timestamp 1621261055
transform 1 0 6912 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_64
timestamp 1621261055
transform 1 0 7296 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_68
timestamp 1621261055
transform 1 0 7680 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_72
timestamp 1621261055
transform 1 0 8064 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_70_82
timestamp 1621261055
transform 1 0 9024 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_80
timestamp 1621261055
transform 1 0 8832 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_76
timestamp 1621261055
transform 1 0 8448 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_80
timestamp 1621261055
transform 1 0 8832 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_910
timestamp 1621261055
transform 1 0 9120 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_92
timestamp 1621261055
transform 1 0 9984 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_84
timestamp 1621261055
transform 1 0 9216 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_88
timestamp 1621261055
transform 1 0 9600 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_96
timestamp 1621261055
transform 1 0 10368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_100
timestamp 1621261055
transform 1 0 10752 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_104
timestamp 1621261055
transform 1 0 11136 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_116
timestamp 1621261055
transform 1 0 12288 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_108
timestamp 1621261055
transform 1 0 11520 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_111
timestamp 1621261055
transform 1 0 11808 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_108
timestamp 1621261055
transform 1 0 11520 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_900
timestamp 1621261055
transform 1 0 11712 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_124
timestamp 1621261055
transform 1 0 13056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_119
timestamp 1621261055
transform 1 0 12576 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_132
timestamp 1621261055
transform 1 0 13824 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_127
timestamp 1621261055
transform 1 0 13344 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_139
timestamp 1621261055
transform 1 0 14496 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_136
timestamp 1621261055
transform 1 0 14208 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_135
timestamp 1621261055
transform 1 0 14112 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_911
timestamp 1621261055
transform 1 0 14400 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_147
timestamp 1621261055
transform 1 0 15264 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_143
timestamp 1621261055
transform 1 0 14880 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_155
timestamp 1621261055
transform 1 0 16032 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_151
timestamp 1621261055
transform 1 0 15648 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_163
timestamp 1621261055
transform 1 0 16800 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_163
timestamp 1621261055
transform 1 0 16800 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_159
timestamp 1621261055
transform 1 0 16416 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_901
timestamp 1621261055
transform 1 0 16992 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_171
timestamp 1621261055
transform 1 0 17568 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_166
timestamp 1621261055
transform 1 0 17088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_179
timestamp 1621261055
transform 1 0 18336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_182
timestamp 1621261055
transform 1 0 18624 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_174
timestamp 1621261055
transform 1 0 17856 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_191
timestamp 1621261055
transform 1 0 19488 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_187
timestamp 1621261055
transform 1 0 19104 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_190
timestamp 1621261055
transform 1 0 19392 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_194
timestamp 1621261055
transform 1 0 19776 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_198
timestamp 1621261055
transform 1 0 20160 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_912
timestamp 1621261055
transform 1 0 19680 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_202
timestamp 1621261055
transform 1 0 20544 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_206
timestamp 1621261055
transform 1 0 20928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_210
timestamp 1621261055
transform 1 0 21312 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_214
timestamp 1621261055
transform 1 0 21696 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_218
timestamp 1621261055
transform 1 0 22080 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_221
timestamp 1621261055
transform 1 0 22368 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_218
timestamp 1621261055
transform 1 0 22080 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_902
timestamp 1621261055
transform 1 0 22272 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_226
timestamp 1621261055
transform 1 0 22848 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_229
timestamp 1621261055
transform 1 0 23136 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_234
timestamp 1621261055
transform 1 0 23616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_237
timestamp 1621261055
transform 1 0 23904 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_246
timestamp 1621261055
transform 1 0 24768 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_242
timestamp 1621261055
transform 1 0 24384 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_245
timestamp 1621261055
transform 1 0 24672 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_913
timestamp 1621261055
transform 1 0 24960 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_257
timestamp 1621261055
transform 1 0 25824 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_249
timestamp 1621261055
transform 1 0 25056 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_253
timestamp 1621261055
transform 1 0 25440 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_261
timestamp 1621261055
transform 1 0 26208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_265
timestamp 1621261055
transform 1 0 26592 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_269
timestamp 1621261055
transform 1 0 26976 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_281
timestamp 1621261055
transform 1 0 28128 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_273
timestamp 1621261055
transform 1 0 27360 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_276
timestamp 1621261055
transform 1 0 27648 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_273
timestamp 1621261055
transform 1 0 27360 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_196
timestamp 1621261055
transform 1 0 27840 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_903
timestamp 1621261055
transform 1 0 27552 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _123_
timestamp 1621261055
transform 1 0 28032 0 1 48618
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_289
timestamp 1621261055
transform 1 0 28896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_283
timestamp 1621261055
transform 1 0 28320 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_297
timestamp 1621261055
transform 1 0 29664 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_291
timestamp 1621261055
transform 1 0 29088 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_304
timestamp 1621261055
transform 1 0 30336 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_301
timestamp 1621261055
transform 1 0 30048 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_299
timestamp 1621261055
transform 1 0 29856 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_914
timestamp 1621261055
transform 1 0 30240 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_312
timestamp 1621261055
transform 1 0 31104 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_307
timestamp 1621261055
transform 1 0 30624 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_320
timestamp 1621261055
transform 1 0 31872 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_323
timestamp 1621261055
transform 1 0 32160 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_315
timestamp 1621261055
transform 1 0 31392 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_70_328
timestamp 1621261055
transform 1 0 32640 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_69_329
timestamp 1621261055
transform 1 0 32736 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_327
timestamp 1621261055
transform 1 0 32544 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_904
timestamp 1621261055
transform 1 0 32832 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_332
timestamp 1621261055
transform 1 0 33024 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_331
timestamp 1621261055
transform 1 0 32928 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_165
timestamp 1621261055
transform -1 0 33408 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _088_
timestamp 1621261055
transform -1 0 33696 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_70_347
timestamp 1621261055
transform 1 0 34464 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_339
timestamp 1621261055
transform 1 0 33696 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_347
timestamp 1621261055
transform 1 0 34464 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_339
timestamp 1621261055
transform 1 0 33696 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_355
timestamp 1621261055
transform 1 0 35232 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_355
timestamp 1621261055
transform 1 0 35232 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_359
timestamp 1621261055
transform 1 0 35616 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_70_357
timestamp 1621261055
transform 1 0 35424 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_69_363
timestamp 1621261055
transform 1 0 36000 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_915
timestamp 1621261055
transform 1 0 35520 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_367
timestamp 1621261055
transform 1 0 36384 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_371
timestamp 1621261055
transform 1 0 36768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_375
timestamp 1621261055
transform 1 0 37152 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_379
timestamp 1621261055
transform 1 0 37536 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_383
timestamp 1621261055
transform 1 0 37920 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_386
timestamp 1621261055
transform 1 0 38208 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_383
timestamp 1621261055
transform 1 0 37920 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_905
timestamp 1621261055
transform 1 0 38112 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_391
timestamp 1621261055
transform 1 0 38688 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_394
timestamp 1621261055
transform 1 0 38976 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_399
timestamp 1621261055
transform 1 0 39456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_402
timestamp 1621261055
transform 1 0 39744 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_411
timestamp 1621261055
transform 1 0 40608 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_407
timestamp 1621261055
transform 1 0 40224 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_410
timestamp 1621261055
transform 1 0 40512 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_916
timestamp 1621261055
transform 1 0 40800 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_422
timestamp 1621261055
transform 1 0 41664 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_414
timestamp 1621261055
transform 1 0 40896 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_418
timestamp 1621261055
transform 1 0 41280 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_426
timestamp 1621261055
transform 1 0 42048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_430
timestamp 1621261055
transform 1 0 42432 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_434
timestamp 1621261055
transform 1 0 42816 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_446
timestamp 1621261055
transform 1 0 43968 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_70_438
timestamp 1621261055
transform 1 0 43200 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_441
timestamp 1621261055
transform 1 0 43488 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_438
timestamp 1621261055
transform 1 0 43200 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_906
timestamp 1621261055
transform 1 0 43392 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_453
timestamp 1621261055
transform 1 0 44640 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_449
timestamp 1621261055
transform 1 0 44256 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_238
timestamp 1621261055
transform -1 0 44352 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _201_
timestamp 1621261055
transform -1 0 44640 0 -1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_70_461
timestamp 1621261055
transform 1 0 45408 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_457
timestamp 1621261055
transform 1 0 45024 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_469
timestamp 1621261055
transform 1 0 46176 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_70_467
timestamp 1621261055
transform 1 0 45984 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_465
timestamp 1621261055
transform 1 0 45792 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_69_465
timestamp 1621261055
transform 1 0 45792 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_917
timestamp 1621261055
transform 1 0 46080 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_477
timestamp 1621261055
transform 1 0 46944 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_473
timestamp 1621261055
transform 1 0 46560 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_485
timestamp 1621261055
transform 1 0 47712 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_481
timestamp 1621261055
transform 1 0 47328 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_493
timestamp 1621261055
transform 1 0 48480 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_493
timestamp 1621261055
transform 1 0 48480 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_69_489
timestamp 1621261055
transform 1 0 48096 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_907
timestamp 1621261055
transform 1 0 48672 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_501
timestamp 1621261055
transform 1 0 49248 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_496
timestamp 1621261055
transform 1 0 48768 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_509
timestamp 1621261055
transform 1 0 50016 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_512
timestamp 1621261055
transform 1 0 50304 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_504
timestamp 1621261055
transform 1 0 49536 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_521
timestamp 1621261055
transform 1 0 51168 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_517
timestamp 1621261055
transform 1 0 50784 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_520
timestamp 1621261055
transform 1 0 51072 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_524
timestamp 1621261055
transform 1 0 51456 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_528
timestamp 1621261055
transform 1 0 51840 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_918
timestamp 1621261055
transform 1 0 51360 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_532
timestamp 1621261055
transform 1 0 52224 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_536
timestamp 1621261055
transform 1 0 52608 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_540
timestamp 1621261055
transform 1 0 52992 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_544
timestamp 1621261055
transform 1 0 53376 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_70_548
timestamp 1621261055
transform 1 0 53760 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_551
timestamp 1621261055
transform 1 0 54048 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_548
timestamp 1621261055
transform 1 0 53760 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_908
timestamp 1621261055
transform 1 0 53952 0 1 48618
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_556
timestamp 1621261055
transform 1 0 54528 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_559
timestamp 1621261055
transform 1 0 54816 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_564
timestamp 1621261055
transform 1 0 55296 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_567
timestamp 1621261055
transform 1 0 55584 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_576
timestamp 1621261055
transform 1 0 56448 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_70_572
timestamp 1621261055
transform 1 0 56064 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_69_575
timestamp 1621261055
transform 1 0 56352 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_919
timestamp 1621261055
transform 1 0 56640 0 -1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_70_587
timestamp 1621261055
transform 1 0 57504 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_70_579
timestamp 1621261055
transform 1 0 56736 0 -1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_69_583
timestamp 1621261055
transform 1 0 57120 0 1 48618
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_69_591
timestamp 1621261055
transform 1 0 57888 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_139
timestamp 1621261055
transform -1 0 58848 0 1 48618
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_141
timestamp 1621261055
transform -1 0 58848 0 -1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_69_595
timestamp 1621261055
transform 1 0 58272 0 1 48618
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_70_595
timestamp 1621261055
transform 1 0 58272 0 -1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_142
timestamp 1621261055
transform 1 0 1152 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_71_4
timestamp 1621261055
transform 1 0 1536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_12
timestamp 1621261055
transform 1 0 2304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_20
timestamp 1621261055
transform 1 0 3072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_28
timestamp 1621261055
transform 1 0 3840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_920
timestamp 1621261055
transform 1 0 6432 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_36
timestamp 1621261055
transform 1 0 4608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_44
timestamp 1621261055
transform 1 0 5376 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_52
timestamp 1621261055
transform 1 0 6144 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_54
timestamp 1621261055
transform 1 0 6336 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_56
timestamp 1621261055
transform 1 0 6528 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_64
timestamp 1621261055
transform 1 0 7296 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _095_
timestamp 1621261055
transform 1 0 10080 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_173
timestamp 1621261055
transform 1 0 9888 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_72
timestamp 1621261055
transform 1 0 8064 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_80
timestamp 1621261055
transform 1 0 8832 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_88
timestamp 1621261055
transform 1 0 9600 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_90
timestamp 1621261055
transform 1 0 9792 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_96
timestamp 1621261055
transform 1 0 10368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_921
timestamp 1621261055
transform 1 0 11712 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_104
timestamp 1621261055
transform 1 0 11136 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_108
timestamp 1621261055
transform 1 0 11520 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_111
timestamp 1621261055
transform 1 0 11808 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_119
timestamp 1621261055
transform 1 0 12576 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_127
timestamp 1621261055
transform 1 0 13344 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_922
timestamp 1621261055
transform 1 0 16992 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_135
timestamp 1621261055
transform 1 0 14112 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_143
timestamp 1621261055
transform 1 0 14880 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_151
timestamp 1621261055
transform 1 0 15648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_159
timestamp 1621261055
transform 1 0 16416 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_163
timestamp 1621261055
transform 1 0 16800 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_166
timestamp 1621261055
transform 1 0 17088 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_174
timestamp 1621261055
transform 1 0 17856 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_182
timestamp 1621261055
transform 1 0 18624 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_190
timestamp 1621261055
transform 1 0 19392 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_198
timestamp 1621261055
transform 1 0 20160 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_923
timestamp 1621261055
transform 1 0 22272 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_206
timestamp 1621261055
transform 1 0 20928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_214
timestamp 1621261055
transform 1 0 21696 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_218
timestamp 1621261055
transform 1 0 22080 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_221
timestamp 1621261055
transform 1 0 22368 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_229
timestamp 1621261055
transform 1 0 23136 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_237
timestamp 1621261055
transform 1 0 23904 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_245
timestamp 1621261055
transform 1 0 24672 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_253
timestamp 1621261055
transform 1 0 25440 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_261
timestamp 1621261055
transform 1 0 26208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_924
timestamp 1621261055
transform 1 0 27552 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_269
timestamp 1621261055
transform 1 0 26976 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_273
timestamp 1621261055
transform 1 0 27360 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_276
timestamp 1621261055
transform 1 0 27648 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_284
timestamp 1621261055
transform 1 0 28416 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_292
timestamp 1621261055
transform 1 0 29184 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_925
timestamp 1621261055
transform 1 0 32832 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_300
timestamp 1621261055
transform 1 0 29952 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_308
timestamp 1621261055
transform 1 0 30720 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_316
timestamp 1621261055
transform 1 0 31488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_324
timestamp 1621261055
transform 1 0 32256 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_328
timestamp 1621261055
transform 1 0 32640 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_331
timestamp 1621261055
transform 1 0 32928 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_339
timestamp 1621261055
transform 1 0 33696 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_347
timestamp 1621261055
transform 1 0 34464 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_355
timestamp 1621261055
transform 1 0 35232 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_363
timestamp 1621261055
transform 1 0 36000 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_926
timestamp 1621261055
transform 1 0 38112 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_371
timestamp 1621261055
transform 1 0 36768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_379
timestamp 1621261055
transform 1 0 37536 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_383
timestamp 1621261055
transform 1 0 37920 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_386
timestamp 1621261055
transform 1 0 38208 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_394
timestamp 1621261055
transform 1 0 38976 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_402
timestamp 1621261055
transform 1 0 39744 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_410
timestamp 1621261055
transform 1 0 40512 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_418
timestamp 1621261055
transform 1 0 41280 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_426
timestamp 1621261055
transform 1 0 42048 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_927
timestamp 1621261055
transform 1 0 43392 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_71_434
timestamp 1621261055
transform 1 0 42816 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_438
timestamp 1621261055
transform 1 0 43200 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_441
timestamp 1621261055
transform 1 0 43488 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_449
timestamp 1621261055
transform 1 0 44256 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_457
timestamp 1621261055
transform 1 0 45024 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_928
timestamp 1621261055
transform 1 0 48672 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_465
timestamp 1621261055
transform 1 0 45792 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_473
timestamp 1621261055
transform 1 0 46560 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_481
timestamp 1621261055
transform 1 0 47328 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_489
timestamp 1621261055
transform 1 0 48096 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_493
timestamp 1621261055
transform 1 0 48480 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_71_496
timestamp 1621261055
transform 1 0 48768 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_504
timestamp 1621261055
transform 1 0 49536 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_512
timestamp 1621261055
transform 1 0 50304 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_520
timestamp 1621261055
transform 1 0 51072 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_528
timestamp 1621261055
transform 1 0 51840 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _052_
timestamp 1621261055
transform 1 0 54720 0 1 49950
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_929
timestamp 1621261055
transform 1 0 53952 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_536
timestamp 1621261055
transform 1 0 52608 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_544
timestamp 1621261055
transform 1 0 53376 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_548
timestamp 1621261055
transform 1 0 53760 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_71_551
timestamp 1621261055
transform 1 0 54048 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_71_555
timestamp 1621261055
transform 1 0 54432 0 1 49950
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_71_557
timestamp 1621261055
transform 1 0 54624 0 1 49950
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_71_561
timestamp 1621261055
transform 1 0 55008 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_569
timestamp 1621261055
transform 1 0 55776 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_577
timestamp 1621261055
transform 1 0 56544 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_71_585
timestamp 1621261055
transform 1 0 57312 0 1 49950
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_71_593
timestamp 1621261055
transform 1 0 58080 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_143
timestamp 1621261055
transform -1 0 58848 0 1 49950
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_144
timestamp 1621261055
transform 1 0 1152 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_930
timestamp 1621261055
transform 1 0 3840 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_4
timestamp 1621261055
transform 1 0 1536 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_12
timestamp 1621261055
transform 1 0 2304 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_20
timestamp 1621261055
transform 1 0 3072 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_29
timestamp 1621261055
transform 1 0 3936 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_37
timestamp 1621261055
transform 1 0 4704 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_45
timestamp 1621261055
transform 1 0 5472 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_53
timestamp 1621261055
transform 1 0 6240 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_61
timestamp 1621261055
transform 1 0 7008 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_69
timestamp 1621261055
transform 1 0 7776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_81
timestamp 1621261055
transform 1 0 8928 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_72_77
timestamp 1621261055
transform 1 0 8544 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_931
timestamp 1621261055
transform 1 0 9120 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_72_91
timestamp 1621261055
transform 1 0 9888 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_84
timestamp 1621261055
transform 1 0 9216 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_252
timestamp 1621261055
transform 1 0 9408 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _211_
timestamp 1621261055
transform 1 0 9600 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__fill_1  FILLER_72_97
timestamp 1621261055
transform 1 0 10464 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_95
timestamp 1621261055
transform 1 0 10272 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_137
timestamp 1621261055
transform 1 0 10560 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _178_
timestamp 1621261055
transform 1 0 10752 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_72_103
timestamp 1621261055
transform 1 0 11040 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_111
timestamp 1621261055
transform 1 0 11808 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_119
timestamp 1621261055
transform 1 0 12576 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_127
timestamp 1621261055
transform 1 0 13344 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_932
timestamp 1621261055
transform 1 0 14400 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_135
timestamp 1621261055
transform 1 0 14112 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_72_137
timestamp 1621261055
transform 1 0 14304 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_139
timestamp 1621261055
transform 1 0 14496 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_147
timestamp 1621261055
transform 1 0 15264 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_155
timestamp 1621261055
transform 1 0 16032 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_163
timestamp 1621261055
transform 1 0 16800 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_933
timestamp 1621261055
transform 1 0 19680 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_171
timestamp 1621261055
transform 1 0 17568 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_179
timestamp 1621261055
transform 1 0 18336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_187
timestamp 1621261055
transform 1 0 19104 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_191
timestamp 1621261055
transform 1 0 19488 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_194
timestamp 1621261055
transform 1 0 19776 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_202
timestamp 1621261055
transform 1 0 20544 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_210
timestamp 1621261055
transform 1 0 21312 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_218
timestamp 1621261055
transform 1 0 22080 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_226
timestamp 1621261055
transform 1 0 22848 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_934
timestamp 1621261055
transform 1 0 24960 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_234
timestamp 1621261055
transform 1 0 23616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_242
timestamp 1621261055
transform 1 0 24384 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_246
timestamp 1621261055
transform 1 0 24768 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_249
timestamp 1621261055
transform 1 0 25056 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_257
timestamp 1621261055
transform 1 0 25824 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_265
timestamp 1621261055
transform 1 0 26592 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_273
timestamp 1621261055
transform 1 0 27360 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_281
timestamp 1621261055
transform 1 0 28128 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_289
timestamp 1621261055
transform 1 0 28896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_297
timestamp 1621261055
transform 1 0 29664 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_935
timestamp 1621261055
transform 1 0 30240 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_301
timestamp 1621261055
transform 1 0 30048 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_304
timestamp 1621261055
transform 1 0 30336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_312
timestamp 1621261055
transform 1 0 31104 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_320
timestamp 1621261055
transform 1 0 31872 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_328
timestamp 1621261055
transform 1 0 32640 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_936
timestamp 1621261055
transform 1 0 35520 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_336
timestamp 1621261055
transform 1 0 33408 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_344
timestamp 1621261055
transform 1 0 34176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_352
timestamp 1621261055
transform 1 0 34944 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_356
timestamp 1621261055
transform 1 0 35328 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_359
timestamp 1621261055
transform 1 0 35616 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_367
timestamp 1621261055
transform 1 0 36384 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_375
timestamp 1621261055
transform 1 0 37152 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_383
timestamp 1621261055
transform 1 0 37920 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_391
timestamp 1621261055
transform 1 0 38688 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_937
timestamp 1621261055
transform 1 0 40800 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_399
timestamp 1621261055
transform 1 0 39456 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_407
timestamp 1621261055
transform 1 0 40224 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_411
timestamp 1621261055
transform 1 0 40608 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_414
timestamp 1621261055
transform 1 0 40896 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_422
timestamp 1621261055
transform 1 0 41664 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_430
timestamp 1621261055
transform 1 0 42432 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_438
timestamp 1621261055
transform 1 0 43200 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_446
timestamp 1621261055
transform 1 0 43968 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_454
timestamp 1621261055
transform 1 0 44736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_462
timestamp 1621261055
transform 1 0 45504 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_938
timestamp 1621261055
transform 1 0 46080 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_466
timestamp 1621261055
transform 1 0 45888 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_72_469
timestamp 1621261055
transform 1 0 46176 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_477
timestamp 1621261055
transform 1 0 46944 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_485
timestamp 1621261055
transform 1 0 47712 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_493
timestamp 1621261055
transform 1 0 48480 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _015_
timestamp 1621261055
transform 1 0 51840 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_939
timestamp 1621261055
transform 1 0 51360 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_501
timestamp 1621261055
transform 1 0 49248 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_509
timestamp 1621261055
transform 1 0 50016 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_72_517
timestamp 1621261055
transform 1 0 50784 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_521
timestamp 1621261055
transform 1 0 51168 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_72_524
timestamp 1621261055
transform 1 0 51456 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _034_
timestamp 1621261055
transform 1 0 52512 0 -1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_72_531
timestamp 1621261055
transform 1 0 52128 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_72_538
timestamp 1621261055
transform 1 0 52800 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_546
timestamp 1621261055
transform 1 0 53568 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_554
timestamp 1621261055
transform 1 0 54336 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_940
timestamp 1621261055
transform 1 0 56640 0 -1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_72_562
timestamp 1621261055
transform 1 0 55104 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_570
timestamp 1621261055
transform 1 0 55872 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_579
timestamp 1621261055
transform 1 0 56736 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_72_587
timestamp 1621261055
transform 1 0 57504 0 -1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_145
timestamp 1621261055
transform -1 0 58848 0 -1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_72_595
timestamp 1621261055
transform 1 0 58272 0 -1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_146
timestamp 1621261055
transform 1 0 1152 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_73_4
timestamp 1621261055
transform 1 0 1536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_12
timestamp 1621261055
transform 1 0 2304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_20
timestamp 1621261055
transform 1 0 3072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_28
timestamp 1621261055
transform 1 0 3840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_941
timestamp 1621261055
transform 1 0 6432 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_36
timestamp 1621261055
transform 1 0 4608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_44
timestamp 1621261055
transform 1 0 5376 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_52
timestamp 1621261055
transform 1 0 6144 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_54
timestamp 1621261055
transform 1 0 6336 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_56
timestamp 1621261055
transform 1 0 6528 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_64
timestamp 1621261055
transform 1 0 7296 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_72
timestamp 1621261055
transform 1 0 8064 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_80
timestamp 1621261055
transform 1 0 8832 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_88
timestamp 1621261055
transform 1 0 9600 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_96
timestamp 1621261055
transform 1 0 10368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_942
timestamp 1621261055
transform 1 0 11712 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_104
timestamp 1621261055
transform 1 0 11136 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_108
timestamp 1621261055
transform 1 0 11520 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_111
timestamp 1621261055
transform 1 0 11808 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_119
timestamp 1621261055
transform 1 0 12576 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_127
timestamp 1621261055
transform 1 0 13344 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_943
timestamp 1621261055
transform 1 0 16992 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_135
timestamp 1621261055
transform 1 0 14112 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_143
timestamp 1621261055
transform 1 0 14880 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_151
timestamp 1621261055
transform 1 0 15648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_159
timestamp 1621261055
transform 1 0 16416 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_163
timestamp 1621261055
transform 1 0 16800 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_166
timestamp 1621261055
transform 1 0 17088 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_174
timestamp 1621261055
transform 1 0 17856 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_182
timestamp 1621261055
transform 1 0 18624 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_190
timestamp 1621261055
transform 1 0 19392 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_198
timestamp 1621261055
transform 1 0 20160 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_944
timestamp 1621261055
transform 1 0 22272 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_206
timestamp 1621261055
transform 1 0 20928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_214
timestamp 1621261055
transform 1 0 21696 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_218
timestamp 1621261055
transform 1 0 22080 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_221
timestamp 1621261055
transform 1 0 22368 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_229
timestamp 1621261055
transform 1 0 23136 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_237
timestamp 1621261055
transform 1 0 23904 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_245
timestamp 1621261055
transform 1 0 24672 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_253
timestamp 1621261055
transform 1 0 25440 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_261
timestamp 1621261055
transform 1 0 26208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_945
timestamp 1621261055
transform 1 0 27552 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_73_269
timestamp 1621261055
transform 1 0 26976 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_273
timestamp 1621261055
transform 1 0 27360 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_276
timestamp 1621261055
transform 1 0 27648 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_284
timestamp 1621261055
transform 1 0 28416 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_292
timestamp 1621261055
transform 1 0 29184 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_946
timestamp 1621261055
transform 1 0 32832 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_300
timestamp 1621261055
transform 1 0 29952 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_308
timestamp 1621261055
transform 1 0 30720 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_316
timestamp 1621261055
transform 1 0 31488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_324
timestamp 1621261055
transform 1 0 32256 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_328
timestamp 1621261055
transform 1 0 32640 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_331
timestamp 1621261055
transform 1 0 32928 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_339
timestamp 1621261055
transform 1 0 33696 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_347
timestamp 1621261055
transform 1 0 34464 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_355
timestamp 1621261055
transform 1 0 35232 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_363
timestamp 1621261055
transform 1 0 36000 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_947
timestamp 1621261055
transform 1 0 38112 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_371
timestamp 1621261055
transform 1 0 36768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_379
timestamp 1621261055
transform 1 0 37536 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_383
timestamp 1621261055
transform 1 0 37920 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_386
timestamp 1621261055
transform 1 0 38208 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_394
timestamp 1621261055
transform 1 0 38976 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _079_
timestamp 1621261055
transform -1 0 41568 0 1 51282
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_151
timestamp 1621261055
transform -1 0 41280 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_402
timestamp 1621261055
transform 1 0 39744 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_410
timestamp 1621261055
transform 1 0 40512 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_414
timestamp 1621261055
transform 1 0 40896 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_421
timestamp 1621261055
transform 1 0 41568 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_429
timestamp 1621261055
transform 1 0 42336 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_948
timestamp 1621261055
transform 1 0 43392 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_437
timestamp 1621261055
transform 1 0 43104 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_73_439
timestamp 1621261055
transform 1 0 43296 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_441
timestamp 1621261055
transform 1 0 43488 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_449
timestamp 1621261055
transform 1 0 44256 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_457
timestamp 1621261055
transform 1 0 45024 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_949
timestamp 1621261055
transform 1 0 48672 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_465
timestamp 1621261055
transform 1 0 45792 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_473
timestamp 1621261055
transform 1 0 46560 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_481
timestamp 1621261055
transform 1 0 47328 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_489
timestamp 1621261055
transform 1 0 48096 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_493
timestamp 1621261055
transform 1 0 48480 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_496
timestamp 1621261055
transform 1 0 48768 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_504
timestamp 1621261055
transform 1 0 49536 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_512
timestamp 1621261055
transform 1 0 50304 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_520
timestamp 1621261055
transform 1 0 51072 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_528
timestamp 1621261055
transform 1 0 51840 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_950
timestamp 1621261055
transform 1 0 53952 0 1 51282
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_73_536
timestamp 1621261055
transform 1 0 52608 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_544
timestamp 1621261055
transform 1 0 53376 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_548
timestamp 1621261055
transform 1 0 53760 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_73_551
timestamp 1621261055
transform 1 0 54048 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_559
timestamp 1621261055
transform 1 0 54816 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_567
timestamp 1621261055
transform 1 0 55584 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_575
timestamp 1621261055
transform 1 0 56352 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_73_583
timestamp 1621261055
transform 1 0 57120 0 1 51282
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_73_591
timestamp 1621261055
transform 1 0 57888 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_147
timestamp 1621261055
transform -1 0 58848 0 1 51282
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_73_595
timestamp 1621261055
transform 1 0 58272 0 1 51282
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_148
timestamp 1621261055
transform 1 0 1152 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_951
timestamp 1621261055
transform 1 0 3840 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_4
timestamp 1621261055
transform 1 0 1536 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_12
timestamp 1621261055
transform 1 0 2304 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_20
timestamp 1621261055
transform 1 0 3072 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_29
timestamp 1621261055
transform 1 0 3936 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_37
timestamp 1621261055
transform 1 0 4704 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_45
timestamp 1621261055
transform 1 0 5472 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_53
timestamp 1621261055
transform 1 0 6240 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_61
timestamp 1621261055
transform 1 0 7008 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_952
timestamp 1621261055
transform 1 0 9120 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_69
timestamp 1621261055
transform 1 0 7776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_77
timestamp 1621261055
transform 1 0 8544 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_81
timestamp 1621261055
transform 1 0 8928 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_84
timestamp 1621261055
transform 1 0 9216 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_92
timestamp 1621261055
transform 1 0 9984 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_100
timestamp 1621261055
transform 1 0 10752 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_108
timestamp 1621261055
transform 1 0 11520 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_116
timestamp 1621261055
transform 1 0 12288 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_124
timestamp 1621261055
transform 1 0 13056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_132
timestamp 1621261055
transform 1 0 13824 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_953
timestamp 1621261055
transform 1 0 14400 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_136
timestamp 1621261055
transform 1 0 14208 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_139
timestamp 1621261055
transform 1 0 14496 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_147
timestamp 1621261055
transform 1 0 15264 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_155
timestamp 1621261055
transform 1 0 16032 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_163
timestamp 1621261055
transform 1 0 16800 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_954
timestamp 1621261055
transform 1 0 19680 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_171
timestamp 1621261055
transform 1 0 17568 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_179
timestamp 1621261055
transform 1 0 18336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_187
timestamp 1621261055
transform 1 0 19104 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_191
timestamp 1621261055
transform 1 0 19488 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_194
timestamp 1621261055
transform 1 0 19776 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_202
timestamp 1621261055
transform 1 0 20544 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_210
timestamp 1621261055
transform 1 0 21312 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_218
timestamp 1621261055
transform 1 0 22080 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_226
timestamp 1621261055
transform 1 0 22848 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_955
timestamp 1621261055
transform 1 0 24960 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_234
timestamp 1621261055
transform 1 0 23616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_242
timestamp 1621261055
transform 1 0 24384 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_246
timestamp 1621261055
transform 1 0 24768 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_249
timestamp 1621261055
transform 1 0 25056 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_257
timestamp 1621261055
transform 1 0 25824 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_265
timestamp 1621261055
transform 1 0 26592 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_273
timestamp 1621261055
transform 1 0 27360 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_281
timestamp 1621261055
transform 1 0 28128 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_289
timestamp 1621261055
transform 1 0 28896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_297
timestamp 1621261055
transform 1 0 29664 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _020_
timestamp 1621261055
transform 1 0 32256 0 -1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_956
timestamp 1621261055
transform 1 0 30240 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_301
timestamp 1621261055
transform 1 0 30048 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_304
timestamp 1621261055
transform 1 0 30336 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_312
timestamp 1621261055
transform 1 0 31104 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_320
timestamp 1621261055
transform 1 0 31872 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_74_327
timestamp 1621261055
transform 1 0 32544 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_957
timestamp 1621261055
transform 1 0 35520 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_335
timestamp 1621261055
transform 1 0 33312 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_343
timestamp 1621261055
transform 1 0 34080 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_351
timestamp 1621261055
transform 1 0 34848 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_355
timestamp 1621261055
transform 1 0 35232 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_74_357
timestamp 1621261055
transform 1 0 35424 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_359
timestamp 1621261055
transform 1 0 35616 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_367
timestamp 1621261055
transform 1 0 36384 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_375
timestamp 1621261055
transform 1 0 37152 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_383
timestamp 1621261055
transform 1 0 37920 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_391
timestamp 1621261055
transform 1 0 38688 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_958
timestamp 1621261055
transform 1 0 40800 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_399
timestamp 1621261055
transform 1 0 39456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_407
timestamp 1621261055
transform 1 0 40224 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_411
timestamp 1621261055
transform 1 0 40608 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_414
timestamp 1621261055
transform 1 0 40896 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_422
timestamp 1621261055
transform 1 0 41664 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_430
timestamp 1621261055
transform 1 0 42432 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_438
timestamp 1621261055
transform 1 0 43200 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_446
timestamp 1621261055
transform 1 0 43968 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_454
timestamp 1621261055
transform 1 0 44736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_462
timestamp 1621261055
transform 1 0 45504 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_959
timestamp 1621261055
transform 1 0 46080 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_466
timestamp 1621261055
transform 1 0 45888 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_469
timestamp 1621261055
transform 1 0 46176 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_477
timestamp 1621261055
transform 1 0 46944 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_485
timestamp 1621261055
transform 1 0 47712 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_493
timestamp 1621261055
transform 1 0 48480 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_960
timestamp 1621261055
transform 1 0 51360 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_501
timestamp 1621261055
transform 1 0 49248 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_509
timestamp 1621261055
transform 1 0 50016 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_517
timestamp 1621261055
transform 1 0 50784 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_521
timestamp 1621261055
transform 1 0 51168 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_524
timestamp 1621261055
transform 1 0 51456 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_532
timestamp 1621261055
transform 1 0 52224 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_540
timestamp 1621261055
transform 1 0 52992 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_548
timestamp 1621261055
transform 1 0 53760 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_556
timestamp 1621261055
transform 1 0 54528 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_961
timestamp 1621261055
transform 1 0 56640 0 -1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_74_564
timestamp 1621261055
transform 1 0 55296 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_74_572
timestamp 1621261055
transform 1 0 56064 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_576
timestamp 1621261055
transform 1 0 56448 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_74_579
timestamp 1621261055
transform 1 0 56736 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_74_587
timestamp 1621261055
transform 1 0 57504 0 -1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_149
timestamp 1621261055
transform -1 0 58848 0 -1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_74_595
timestamp 1621261055
transform 1 0 58272 0 -1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_150
timestamp 1621261055
transform 1 0 1152 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_75_4
timestamp 1621261055
transform 1 0 1536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_12
timestamp 1621261055
transform 1 0 2304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_20
timestamp 1621261055
transform 1 0 3072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_28
timestamp 1621261055
transform 1 0 3840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_962
timestamp 1621261055
transform 1 0 6432 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_36
timestamp 1621261055
transform 1 0 4608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_44
timestamp 1621261055
transform 1 0 5376 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_52
timestamp 1621261055
transform 1 0 6144 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_54
timestamp 1621261055
transform 1 0 6336 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_56
timestamp 1621261055
transform 1 0 6528 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_64
timestamp 1621261055
transform 1 0 7296 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_72
timestamp 1621261055
transform 1 0 8064 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_80
timestamp 1621261055
transform 1 0 8832 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_88
timestamp 1621261055
transform 1 0 9600 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_96
timestamp 1621261055
transform 1 0 10368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _186_
timestamp 1621261055
transform -1 0 12864 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_963
timestamp 1621261055
transform 1 0 11712 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_254
timestamp 1621261055
transform -1 0 12576 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_75_104
timestamp 1621261055
transform 1 0 11136 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_108
timestamp 1621261055
transform 1 0 11520 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_75_111
timestamp 1621261055
transform 1 0 11808 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_115
timestamp 1621261055
transform 1 0 12192 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_122
timestamp 1621261055
transform 1 0 12864 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_130
timestamp 1621261055
transform 1 0 13632 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_964
timestamp 1621261055
transform 1 0 16992 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_138
timestamp 1621261055
transform 1 0 14400 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_146
timestamp 1621261055
transform 1 0 15168 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_154
timestamp 1621261055
transform 1 0 15936 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_162
timestamp 1621261055
transform 1 0 16704 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_164
timestamp 1621261055
transform 1 0 16896 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_166
timestamp 1621261055
transform 1 0 17088 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_174
timestamp 1621261055
transform 1 0 17856 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_182
timestamp 1621261055
transform 1 0 18624 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_190
timestamp 1621261055
transform 1 0 19392 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_198
timestamp 1621261055
transform 1 0 20160 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_965
timestamp 1621261055
transform 1 0 22272 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_246
timestamp 1621261055
transform -1 0 23520 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_206
timestamp 1621261055
transform 1 0 20928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_214
timestamp 1621261055
transform 1 0 21696 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_218
timestamp 1621261055
transform 1 0 22080 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_221
timestamp 1621261055
transform 1 0 22368 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_229
timestamp 1621261055
transform 1 0 23136 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _206_
timestamp 1621261055
transform -1 0 23808 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_75_236
timestamp 1621261055
transform 1 0 23808 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_244
timestamp 1621261055
transform 1 0 24576 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_252
timestamp 1621261055
transform 1 0 25344 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_260
timestamp 1621261055
transform 1 0 26112 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_966
timestamp 1621261055
transform 1 0 27552 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_75_268
timestamp 1621261055
transform 1 0 26880 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_272
timestamp 1621261055
transform 1 0 27264 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_75_274
timestamp 1621261055
transform 1 0 27456 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_276
timestamp 1621261055
transform 1 0 27648 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_284
timestamp 1621261055
transform 1 0 28416 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_292
timestamp 1621261055
transform 1 0 29184 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_967
timestamp 1621261055
transform 1 0 32832 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_300
timestamp 1621261055
transform 1 0 29952 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_308
timestamp 1621261055
transform 1 0 30720 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_316
timestamp 1621261055
transform 1 0 31488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_324
timestamp 1621261055
transform 1 0 32256 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_328
timestamp 1621261055
transform 1 0 32640 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_331
timestamp 1621261055
transform 1 0 32928 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_339
timestamp 1621261055
transform 1 0 33696 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_347
timestamp 1621261055
transform 1 0 34464 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_355
timestamp 1621261055
transform 1 0 35232 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_363
timestamp 1621261055
transform 1 0 36000 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_968
timestamp 1621261055
transform 1 0 38112 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_371
timestamp 1621261055
transform 1 0 36768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_379
timestamp 1621261055
transform 1 0 37536 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_383
timestamp 1621261055
transform 1 0 37920 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_386
timestamp 1621261055
transform 1 0 38208 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_394
timestamp 1621261055
transform 1 0 38976 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _085_
timestamp 1621261055
transform -1 0 40992 0 1 52614
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_159
timestamp 1621261055
transform -1 0 40704 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_402
timestamp 1621261055
transform 1 0 39744 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_415
timestamp 1621261055
transform 1 0 40992 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_423
timestamp 1621261055
transform 1 0 41760 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_969
timestamp 1621261055
transform 1 0 43392 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_431
timestamp 1621261055
transform 1 0 42528 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_75_439
timestamp 1621261055
transform 1 0 43296 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_441
timestamp 1621261055
transform 1 0 43488 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_449
timestamp 1621261055
transform 1 0 44256 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_457
timestamp 1621261055
transform 1 0 45024 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_970
timestamp 1621261055
transform 1 0 48672 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_465
timestamp 1621261055
transform 1 0 45792 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_473
timestamp 1621261055
transform 1 0 46560 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_481
timestamp 1621261055
transform 1 0 47328 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_489
timestamp 1621261055
transform 1 0 48096 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_493
timestamp 1621261055
transform 1 0 48480 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_496
timestamp 1621261055
transform 1 0 48768 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_504
timestamp 1621261055
transform 1 0 49536 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_512
timestamp 1621261055
transform 1 0 50304 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_520
timestamp 1621261055
transform 1 0 51072 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_528
timestamp 1621261055
transform 1 0 51840 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_971
timestamp 1621261055
transform 1 0 53952 0 1 52614
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_75_536
timestamp 1621261055
transform 1 0 52608 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_544
timestamp 1621261055
transform 1 0 53376 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_548
timestamp 1621261055
transform 1 0 53760 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_75_551
timestamp 1621261055
transform 1 0 54048 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_559
timestamp 1621261055
transform 1 0 54816 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_567
timestamp 1621261055
transform 1 0 55584 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_575
timestamp 1621261055
transform 1 0 56352 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_75_583
timestamp 1621261055
transform 1 0 57120 0 1 52614
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_75_591
timestamp 1621261055
transform 1 0 57888 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_151
timestamp 1621261055
transform -1 0 58848 0 1 52614
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_75_595
timestamp 1621261055
transform 1 0 58272 0 1 52614
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  PHY_152
timestamp 1621261055
transform 1 0 1152 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_972
timestamp 1621261055
transform 1 0 3840 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_4
timestamp 1621261055
transform 1 0 1536 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_12
timestamp 1621261055
transform 1 0 2304 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_20
timestamp 1621261055
transform 1 0 3072 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_29
timestamp 1621261055
transform 1 0 3936 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _174_
timestamp 1621261055
transform 1 0 5280 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__diode_2  ANTENNA_132
timestamp 1621261055
transform 1 0 5088 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_76_37
timestamp 1621261055
transform 1 0 4704 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_76_46
timestamp 1621261055
transform 1 0 5568 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_54
timestamp 1621261055
transform 1 0 6336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_62
timestamp 1621261055
transform 1 0 7104 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_66
timestamp 1621261055
transform 1 0 7488 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _087_
timestamp 1621261055
transform 1 0 7968 0 -1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_973
timestamp 1621261055
transform 1 0 9120 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_163
timestamp 1621261055
transform 1 0 7776 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_76_68
timestamp 1621261055
transform 1 0 7680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_74
timestamp 1621261055
transform 1 0 8256 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_76_82
timestamp 1621261055
transform 1 0 9024 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_84
timestamp 1621261055
transform 1 0 9216 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_92
timestamp 1621261055
transform 1 0 9984 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_100
timestamp 1621261055
transform 1 0 10752 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_108
timestamp 1621261055
transform 1 0 11520 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_116
timestamp 1621261055
transform 1 0 12288 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_124
timestamp 1621261055
transform 1 0 13056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_132
timestamp 1621261055
transform 1 0 13824 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_974
timestamp 1621261055
transform 1 0 14400 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_136
timestamp 1621261055
transform 1 0 14208 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_139
timestamp 1621261055
transform 1 0 14496 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_147
timestamp 1621261055
transform 1 0 15264 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_155
timestamp 1621261055
transform 1 0 16032 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_163
timestamp 1621261055
transform 1 0 16800 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_975
timestamp 1621261055
transform 1 0 19680 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_171
timestamp 1621261055
transform 1 0 17568 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_179
timestamp 1621261055
transform 1 0 18336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_187
timestamp 1621261055
transform 1 0 19104 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_191
timestamp 1621261055
transform 1 0 19488 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_194
timestamp 1621261055
transform 1 0 19776 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_202
timestamp 1621261055
transform 1 0 20544 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_210
timestamp 1621261055
transform 1 0 21312 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_218
timestamp 1621261055
transform 1 0 22080 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_226
timestamp 1621261055
transform 1 0 22848 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_976
timestamp 1621261055
transform 1 0 24960 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_234
timestamp 1621261055
transform 1 0 23616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_242
timestamp 1621261055
transform 1 0 24384 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_246
timestamp 1621261055
transform 1 0 24768 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_249
timestamp 1621261055
transform 1 0 25056 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_257
timestamp 1621261055
transform 1 0 25824 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_265
timestamp 1621261055
transform 1 0 26592 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_273
timestamp 1621261055
transform 1 0 27360 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_281
timestamp 1621261055
transform 1 0 28128 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_289
timestamp 1621261055
transform 1 0 28896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_297
timestamp 1621261055
transform 1 0 29664 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_977
timestamp 1621261055
transform 1 0 30240 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_301
timestamp 1621261055
transform 1 0 30048 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_304
timestamp 1621261055
transform 1 0 30336 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_312
timestamp 1621261055
transform 1 0 31104 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_320
timestamp 1621261055
transform 1 0 31872 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_328
timestamp 1621261055
transform 1 0 32640 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_978
timestamp 1621261055
transform 1 0 35520 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_336
timestamp 1621261055
transform 1 0 33408 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_344
timestamp 1621261055
transform 1 0 34176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_352
timestamp 1621261055
transform 1 0 34944 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_356
timestamp 1621261055
transform 1 0 35328 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_359
timestamp 1621261055
transform 1 0 35616 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_367
timestamp 1621261055
transform 1 0 36384 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_375
timestamp 1621261055
transform 1 0 37152 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_383
timestamp 1621261055
transform 1 0 37920 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_391
timestamp 1621261055
transform 1 0 38688 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_979
timestamp 1621261055
transform 1 0 40800 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_399
timestamp 1621261055
transform 1 0 39456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_407
timestamp 1621261055
transform 1 0 40224 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_411
timestamp 1621261055
transform 1 0 40608 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_414
timestamp 1621261055
transform 1 0 40896 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_422
timestamp 1621261055
transform 1 0 41664 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_430
timestamp 1621261055
transform 1 0 42432 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_438
timestamp 1621261055
transform 1 0 43200 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_446
timestamp 1621261055
transform 1 0 43968 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_454
timestamp 1621261055
transform 1 0 44736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_462
timestamp 1621261055
transform 1 0 45504 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_980
timestamp 1621261055
transform 1 0 46080 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_466
timestamp 1621261055
transform 1 0 45888 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_469
timestamp 1621261055
transform 1 0 46176 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_477
timestamp 1621261055
transform 1 0 46944 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_485
timestamp 1621261055
transform 1 0 47712 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_493
timestamp 1621261055
transform 1 0 48480 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_981
timestamp 1621261055
transform 1 0 51360 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_76_501
timestamp 1621261055
transform 1 0 49248 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_509
timestamp 1621261055
transform 1 0 50016 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_517
timestamp 1621261055
transform 1 0 50784 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_521
timestamp 1621261055
transform 1 0 51168 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_524
timestamp 1621261055
transform 1 0 51456 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_532
timestamp 1621261055
transform 1 0 52224 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_540
timestamp 1621261055
transform 1 0 52992 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_548
timestamp 1621261055
transform 1 0 53760 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_76_556
timestamp 1621261055
transform 1 0 54528 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_982
timestamp 1621261055
transform 1 0 56640 0 -1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output436
timestamp 1621261055
transform -1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_86
timestamp 1621261055
transform -1 0 57696 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_564
timestamp 1621261055
transform 1 0 55296 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_572
timestamp 1621261055
transform 1 0 56064 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_76_576
timestamp 1621261055
transform 1 0 56448 0 -1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_76_579
timestamp 1621261055
transform 1 0 56736 0 -1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_76_593
timestamp 1621261055
transform 1 0 58080 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_153
timestamp 1621261055
transform -1 0 58848 0 -1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_4
timestamp 1621261055
transform 1 0 1536 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_4
timestamp 1621261055
transform 1 0 1536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_156
timestamp 1621261055
transform 1 0 1152 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_154
timestamp 1621261055
transform 1 0 1152 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_12
timestamp 1621261055
transform 1 0 2304 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_16
timestamp 1621261055
transform 1 0 2688 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_12
timestamp 1621261055
transform 1 0 2304 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _005_
timestamp 1621261055
transform 1 0 2400 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_20
timestamp 1621261055
transform 1 0 3072 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_24
timestamp 1621261055
transform 1 0 3456 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_29
timestamp 1621261055
transform 1 0 3936 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_32
timestamp 1621261055
transform 1 0 4224 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_993
timestamp 1621261055
transform 1 0 3840 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_37
timestamp 1621261055
transform 1 0 4704 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_40
timestamp 1621261055
transform 1 0 4992 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_45
timestamp 1621261055
transform 1 0 5472 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_48
timestamp 1621261055
transform 1 0 5760 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_53
timestamp 1621261055
transform 1 0 6240 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_56
timestamp 1621261055
transform 1 0 6528 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_54
timestamp 1621261055
transform 1 0 6336 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_52
timestamp 1621261055
transform 1 0 6144 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_983
timestamp 1621261055
transform 1 0 6432 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_61
timestamp 1621261055
transform 1 0 7008 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_64
timestamp 1621261055
transform 1 0 7296 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_69
timestamp 1621261055
transform 1 0 7776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_72
timestamp 1621261055
transform 1 0 8064 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_81
timestamp 1621261055
transform 1 0 8928 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_77
timestamp 1621261055
transform 1 0 8544 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_80
timestamp 1621261055
transform 1 0 8832 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_994
timestamp 1621261055
transform 1 0 9120 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_92
timestamp 1621261055
transform 1 0 9984 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_84
timestamp 1621261055
transform 1 0 9216 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_88
timestamp 1621261055
transform 1 0 9600 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_96
timestamp 1621261055
transform 1 0 10368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_100
timestamp 1621261055
transform 1 0 10752 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_104
timestamp 1621261055
transform 1 0 11136 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_116
timestamp 1621261055
transform 1 0 12288 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_108
timestamp 1621261055
transform 1 0 11520 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_111
timestamp 1621261055
transform 1 0 11808 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_108
timestamp 1621261055
transform 1 0 11520 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_984
timestamp 1621261055
transform 1 0 11712 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_124
timestamp 1621261055
transform 1 0 13056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_119
timestamp 1621261055
transform 1 0 12576 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_132
timestamp 1621261055
transform 1 0 13824 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_127
timestamp 1621261055
transform 1 0 13344 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_139
timestamp 1621261055
transform 1 0 14496 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_136
timestamp 1621261055
transform 1 0 14208 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_135
timestamp 1621261055
transform 1 0 14112 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_995
timestamp 1621261055
transform 1 0 14400 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_147
timestamp 1621261055
transform 1 0 15264 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_143
timestamp 1621261055
transform 1 0 14880 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_155
timestamp 1621261055
transform 1 0 16032 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_151
timestamp 1621261055
transform 1 0 15648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_163
timestamp 1621261055
transform 1 0 16800 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_163
timestamp 1621261055
transform 1 0 16800 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_159
timestamp 1621261055
transform 1 0 16416 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_985
timestamp 1621261055
transform 1 0 16992 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_171
timestamp 1621261055
transform 1 0 17568 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_166
timestamp 1621261055
transform 1 0 17088 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_179
timestamp 1621261055
transform 1 0 18336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_182
timestamp 1621261055
transform 1 0 18624 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_174
timestamp 1621261055
transform 1 0 17856 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_191
timestamp 1621261055
transform 1 0 19488 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_187
timestamp 1621261055
transform 1 0 19104 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_190
timestamp 1621261055
transform 1 0 19392 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_194
timestamp 1621261055
transform 1 0 19776 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_198
timestamp 1621261055
transform 1 0 20160 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_996
timestamp 1621261055
transform 1 0 19680 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_202
timestamp 1621261055
transform 1 0 20544 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_206
timestamp 1621261055
transform 1 0 20928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_214
timestamp 1621261055
transform 1 0 21696 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_210
timestamp 1621261055
transform 1 0 21312 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_77_214
timestamp 1621261055
transform 1 0 21696 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_219
timestamp 1621261055
transform 1 0 22176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_221
timestamp 1621261055
transform 1 0 22368 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_218
timestamp 1621261055
transform 1 0 22080 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_986
timestamp 1621261055
transform 1 0 22272 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _051_
timestamp 1621261055
transform 1 0 21888 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_227
timestamp 1621261055
transform 1 0 22944 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_229
timestamp 1621261055
transform 1 0 23136 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_235
timestamp 1621261055
transform 1 0 23712 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_237
timestamp 1621261055
transform 1 0 23904 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_247
timestamp 1621261055
transform 1 0 24864 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_243
timestamp 1621261055
transform 1 0 24480 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_245
timestamp 1621261055
transform 1 0 24672 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_997
timestamp 1621261055
transform 1 0 24960 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_257
timestamp 1621261055
transform 1 0 25824 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_249
timestamp 1621261055
transform 1 0 25056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_253
timestamp 1621261055
transform 1 0 25440 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_261
timestamp 1621261055
transform 1 0 26208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_269
timestamp 1621261055
transform 1 0 26976 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_265
timestamp 1621261055
transform 1 0 26592 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_77_269
timestamp 1621261055
transform 1 0 26976 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__conb_1  _022_
timestamp 1621261055
transform 1 0 26688 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_277
timestamp 1621261055
transform 1 0 27744 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_276
timestamp 1621261055
transform 1 0 27648 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_273
timestamp 1621261055
transform 1 0 27360 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_987
timestamp 1621261055
transform 1 0 27552 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_285
timestamp 1621261055
transform 1 0 28512 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_284
timestamp 1621261055
transform 1 0 28416 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_293
timestamp 1621261055
transform 1 0 29280 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_292
timestamp 1621261055
transform 1 0 29184 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_304
timestamp 1621261055
transform 1 0 30336 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_301
timestamp 1621261055
transform 1 0 30048 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_300
timestamp 1621261055
transform 1 0 29952 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_998
timestamp 1621261055
transform 1 0 30240 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_312
timestamp 1621261055
transform 1 0 31104 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_313
timestamp 1621261055
transform 1 0 31200 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_183
timestamp 1621261055
transform 1 0 30720 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _107_
timestamp 1621261055
transform 1 0 30912 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_320
timestamp 1621261055
transform 1 0 31872 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_321
timestamp 1621261055
transform 1 0 31968 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_328
timestamp 1621261055
transform 1 0 32640 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_329
timestamp 1621261055
transform 1 0 32736 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_988
timestamp 1621261055
transform 1 0 32832 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_336
timestamp 1621261055
transform 1 0 33408 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_331
timestamp 1621261055
transform 1 0 32928 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_344
timestamp 1621261055
transform 1 0 34176 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_347
timestamp 1621261055
transform 1 0 34464 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_339
timestamp 1621261055
transform 1 0 33696 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_356
timestamp 1621261055
transform 1 0 35328 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_352
timestamp 1621261055
transform 1 0 34944 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_355
timestamp 1621261055
transform 1 0 35232 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_359
timestamp 1621261055
transform 1 0 35616 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_363
timestamp 1621261055
transform 1 0 36000 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_999
timestamp 1621261055
transform 1 0 35520 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_367
timestamp 1621261055
transform 1 0 36384 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_371
timestamp 1621261055
transform 1 0 36768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_130
timestamp 1621261055
transform -1 0 36768 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _067_
timestamp 1621261055
transform -1 0 37056 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_374
timestamp 1621261055
transform 1 0 37056 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_379
timestamp 1621261055
transform 1 0 37536 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_78_382
timestamp 1621261055
transform 1 0 37824 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_386
timestamp 1621261055
transform 1 0 38208 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_383
timestamp 1621261055
transform 1 0 37920 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_989
timestamp 1621261055
transform 1 0 38112 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_390
timestamp 1621261055
transform 1 0 38592 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_394
timestamp 1621261055
transform 1 0 38976 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_398
timestamp 1621261055
transform 1 0 39360 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_402
timestamp 1621261055
transform 1 0 39744 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_412
timestamp 1621261055
transform 1 0 40704 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_410
timestamp 1621261055
transform 1 0 40512 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_406
timestamp 1621261055
transform 1 0 40128 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_410
timestamp 1621261055
transform 1 0 40512 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1000
timestamp 1621261055
transform 1 0 40800 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_422
timestamp 1621261055
transform 1 0 41664 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_414
timestamp 1621261055
transform 1 0 40896 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_418
timestamp 1621261055
transform 1 0 41280 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_426
timestamp 1621261055
transform 1 0 42048 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_227
timestamp 1621261055
transform -1 0 42336 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _182_
timestamp 1621261055
transform -1 0 42624 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_430
timestamp 1621261055
transform 1 0 42432 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_432
timestamp 1621261055
transform 1 0 42624 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_446
timestamp 1621261055
transform 1 0 43968 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_438
timestamp 1621261055
transform 1 0 43200 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_441
timestamp 1621261055
transform 1 0 43488 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_990
timestamp 1621261055
transform 1 0 43392 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_454
timestamp 1621261055
transform 1 0 44736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_453
timestamp 1621261055
transform 1 0 44640 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_77_449
timestamp 1621261055
transform 1 0 44256 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_109
timestamp 1621261055
transform 1 0 44832 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_462
timestamp 1621261055
transform 1 0 45504 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_460
timestamp 1621261055
transform 1 0 45312 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _159_
timestamp 1621261055
transform 1 0 45024 0 1 53946
box -38 -49 326 715
use sky130_fd_sc_ls__decap_4  FILLER_78_469
timestamp 1621261055
transform 1 0 46176 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_466
timestamp 1621261055
transform 1 0 45888 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_77_468
timestamp 1621261055
transform 1 0 46080 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1001
timestamp 1621261055
transform 1 0 46080 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_478
timestamp 1621261055
transform 1 0 47040 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_476
timestamp 1621261055
transform 1 0 46848 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_233
timestamp 1621261055
transform -1 0 46752 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _198_
timestamp 1621261055
transform -1 0 47040 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_486
timestamp 1621261055
transform 1 0 47808 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_484
timestamp 1621261055
transform 1 0 47616 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_494
timestamp 1621261055
transform 1 0 48576 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_77_494
timestamp 1621261055
transform 1 0 48576 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_492
timestamp 1621261055
transform 1 0 48384 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_991
timestamp 1621261055
transform 1 0 48672 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_502
timestamp 1621261055
transform 1 0 49344 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_496
timestamp 1621261055
transform 1 0 48768 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_510
timestamp 1621261055
transform 1 0 50112 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_512
timestamp 1621261055
transform 1 0 50304 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_504
timestamp 1621261055
transform 1 0 49536 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_78_518
timestamp 1621261055
transform 1 0 50880 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_520
timestamp 1621261055
transform 1 0 51072 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_524
timestamp 1621261055
transform 1 0 51456 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_78_522
timestamp 1621261055
transform 1 0 51264 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_77_528
timestamp 1621261055
transform 1 0 51840 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1002
timestamp 1621261055
transform 1 0 51360 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_78_532
timestamp 1621261055
transform 1 0 52224 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_536
timestamp 1621261055
transform 1 0 52608 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_540
timestamp 1621261055
transform 1 0 52992 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_544
timestamp 1621261055
transform 1 0 53376 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_78_552
timestamp 1621261055
transform 1 0 54144 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_78_548
timestamp 1621261055
transform 1 0 53760 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_551
timestamp 1621261055
transform 1 0 54048 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_77_548
timestamp 1621261055
transform 1 0 53760 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_992
timestamp 1621261055
transform 1 0 53952 0 1 53946
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _031_
timestamp 1621261055
transform 1 0 54240 0 -1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__decap_8  FILLER_78_556
timestamp 1621261055
transform 1 0 54528 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_559
timestamp 1621261055
transform 1 0 54816 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_78_564
timestamp 1621261055
transform 1 0 55296 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_77_567
timestamp 1621261055
transform 1 0 55584 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_576
timestamp 1621261055
transform 1 0 56448 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_572
timestamp 1621261055
transform 1 0 56064 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_77_575
timestamp 1621261055
transform 1 0 56352 0 1 53946
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1003
timestamp 1621261055
transform 1 0 56640 0 -1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_78_587
timestamp 1621261055
transform 1 0 57504 0 -1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_78_579
timestamp 1621261055
transform 1 0 56736 0 -1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_77_583
timestamp 1621261055
transform 1 0 57120 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_84
timestamp 1621261055
transform -1 0 57696 0 1 53946
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_78_593
timestamp 1621261055
transform 1 0 58080 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_77_593
timestamp 1621261055
transform 1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output435
timestamp 1621261055
transform -1 0 58080 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output398
timestamp 1621261055
transform 1 0 57696 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_155
timestamp 1621261055
transform -1 0 58848 0 1 53946
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_157
timestamp 1621261055
transform -1 0 58848 0 -1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_158
timestamp 1621261055
transform 1 0 1152 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output406
timestamp 1621261055
transform 1 0 1536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output428
timestamp 1621261055
transform 1 0 4320 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_36
timestamp 1621261055
transform 1 0 1920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_72
timestamp 1621261055
transform 1 0 4128 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_10
timestamp 1621261055
transform 1 0 2112 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_18
timestamp 1621261055
transform 1 0 2880 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_26
timestamp 1621261055
transform 1 0 3648 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_30
timestamp 1621261055
transform 1 0 4032 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1004
timestamp 1621261055
transform 1 0 6432 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output438
timestamp 1621261055
transform 1 0 7488 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_37
timestamp 1621261055
transform 1 0 4704 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_45
timestamp 1621261055
transform 1 0 5472 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_53
timestamp 1621261055
transform 1 0 6240 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_56
timestamp 1621261055
transform 1 0 6528 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_64
timestamp 1621261055
transform 1 0 7296 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _156_
timestamp 1621261055
transform 1 0 8256 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output439
timestamp 1621261055
transform -1 0 9504 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_88
timestamp 1621261055
transform -1 0 9120 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_106
timestamp 1621261055
transform 1 0 8064 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_70
timestamp 1621261055
transform 1 0 7872 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_77
timestamp 1621261055
transform 1 0 8544 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_87
timestamp 1621261055
transform 1 0 9504 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_95
timestamp 1621261055
transform 1 0 10272 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_107
timestamp 1621261055
transform 1 0 11424 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_103
timestamp 1621261055
transform 1 0 11040 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_111
timestamp 1621261055
transform 1 0 11808 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_79_109
timestamp 1621261055
transform 1 0 11616 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1005
timestamp 1621261055
transform 1 0 11712 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_119
timestamp 1621261055
transform 1 0 12576 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_79_129
timestamp 1621261055
transform 1 0 13536 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_127
timestamp 1621261055
transform 1 0 13344 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_94
timestamp 1621261055
transform 1 0 13632 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output442
timestamp 1621261055
transform 1 0 13824 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1006
timestamp 1621261055
transform 1 0 16992 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_136
timestamp 1621261055
transform 1 0 14208 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_144
timestamp 1621261055
transform 1 0 14976 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_152
timestamp 1621261055
transform 1 0 15744 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_160
timestamp 1621261055
transform 1 0 16512 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_164
timestamp 1621261055
transform 1 0 16896 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _086_
timestamp 1621261055
transform 1 0 18048 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output409
timestamp 1621261055
transform 1 0 20160 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_161
timestamp 1621261055
transform 1 0 17856 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_166
timestamp 1621261055
transform 1 0 17088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_179
timestamp 1621261055
transform 1 0 18336 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_187
timestamp 1621261055
transform 1 0 19104 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_195
timestamp 1621261055
transform 1 0 19872 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_197
timestamp 1621261055
transform 1 0 20064 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__conb_1  _029_
timestamp 1621261055
transform 1 0 21216 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1007
timestamp 1621261055
transform 1 0 22272 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output411
timestamp 1621261055
transform -1 0 23712 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_44
timestamp 1621261055
transform -1 0 23328 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_202
timestamp 1621261055
transform 1 0 20544 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_206
timestamp 1621261055
transform 1 0 20928 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_208
timestamp 1621261055
transform 1 0 21120 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_212
timestamp 1621261055
transform 1 0 21504 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_221
timestamp 1621261055
transform 1 0 22368 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output412
timestamp 1621261055
transform -1 0 25248 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_46
timestamp 1621261055
transform -1 0 24864 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_235
timestamp 1621261055
transform 1 0 23712 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_243
timestamp 1621261055
transform 1 0 24480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_251
timestamp 1621261055
transform 1 0 25248 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_259
timestamp 1621261055
transform 1 0 26016 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _193_
timestamp 1621261055
transform -1 0 29184 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1008
timestamp 1621261055
transform 1 0 27552 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_229
timestamp 1621261055
transform -1 0 28896 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_267
timestamp 1621261055
transform 1 0 26784 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_276
timestamp 1621261055
transform 1 0 27648 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_284
timestamp 1621261055
transform 1 0 28416 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_286
timestamp 1621261055
transform 1 0 28608 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_79_292
timestamp 1621261055
transform 1 0 29184 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_296
timestamp 1621261055
transform 1 0 29568 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _177_
timestamp 1621261055
transform 1 0 29952 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1009
timestamp 1621261055
transform 1 0 32832 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_135
timestamp 1621261055
transform 1 0 29760 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_303
timestamp 1621261055
transform 1 0 30240 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_311
timestamp 1621261055
transform 1 0 31008 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_319
timestamp 1621261055
transform 1 0 31776 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_327
timestamp 1621261055
transform 1 0 32544 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_329
timestamp 1621261055
transform 1 0 32736 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_331
timestamp 1621261055
transform 1 0 32928 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_339
timestamp 1621261055
transform 1 0 33696 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_347
timestamp 1621261055
transform 1 0 34464 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_355
timestamp 1621261055
transform 1 0 35232 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_363
timestamp 1621261055
transform 1 0 36000 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1010
timestamp 1621261055
transform 1 0 38112 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output422
timestamp 1621261055
transform -1 0 39456 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_64
timestamp 1621261055
transform -1 0 39072 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_371
timestamp 1621261055
transform 1 0 36768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_379
timestamp 1621261055
transform 1 0 37536 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_383
timestamp 1621261055
transform 1 0 37920 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_386
timestamp 1621261055
transform 1 0 38208 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_390
timestamp 1621261055
transform 1 0 38592 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_392
timestamp 1621261055
transform 1 0 38784 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output423
timestamp 1621261055
transform 1 0 40704 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_79_399
timestamp 1621261055
transform 1 0 39456 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_407
timestamp 1621261055
transform 1 0 40224 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_411
timestamp 1621261055
transform 1 0 40608 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_79_416
timestamp 1621261055
transform 1 0 41088 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_424
timestamp 1621261055
transform 1 0 41856 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1011
timestamp 1621261055
transform 1 0 43392 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output426
timestamp 1621261055
transform -1 0 45792 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_68
timestamp 1621261055
transform -1 0 45408 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_432
timestamp 1621261055
transform 1 0 42624 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_441
timestamp 1621261055
transform 1 0 43488 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_449
timestamp 1621261055
transform 1 0 44256 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_457
timestamp 1621261055
transform 1 0 45024 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1012
timestamp 1621261055
transform 1 0 48672 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output427
timestamp 1621261055
transform -1 0 47328 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_70
timestamp 1621261055
transform -1 0 46944 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_465
timestamp 1621261055
transform 1 0 45792 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_473
timestamp 1621261055
transform 1 0 46560 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_481
timestamp 1621261055
transform 1 0 47328 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_79_489
timestamp 1621261055
transform 1 0 48096 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_493
timestamp 1621261055
transform 1 0 48480 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _081_
timestamp 1621261055
transform -1 0 50784 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__clkbuf_2  output431
timestamp 1621261055
transform -1 0 52128 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_75
timestamp 1621261055
transform -1 0 51744 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_155
timestamp 1621261055
transform -1 0 50496 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_496
timestamp 1621261055
transform 1 0 48768 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_504
timestamp 1621261055
transform 1 0 49536 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_517
timestamp 1621261055
transform 1 0 50784 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__conb_1  _072_
timestamp 1621261055
transform -1 0 54720 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1013
timestamp 1621261055
transform 1 0 53952 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_145
timestamp 1621261055
transform -1 0 54432 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_531
timestamp 1621261055
transform 1 0 52128 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__decap_8  FILLER_79_539
timestamp 1621261055
transform 1 0 52896 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_547
timestamp 1621261055
transform 1 0 53664 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_79_549
timestamp 1621261055
transform 1 0 53856 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_551
timestamp 1621261055
transform 1 0 54048 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_79_558
timestamp 1621261055
transform 1 0 54720 0 1 55278
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_79_566
timestamp 1621261055
transform 1 0 55488 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_177
timestamp 1621261055
transform -1 0 55776 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__conb_1  _098_
timestamp 1621261055
transform -1 0 56064 0 1 55278
box -38 -49 326 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_572
timestamp 1621261055
transform 1 0 56064 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_82
timestamp 1621261055
transform 1 0 56256 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_79_580
timestamp 1621261055
transform 1 0 56832 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output434
timestamp 1621261055
transform 1 0 56448 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_79_584
timestamp 1621261055
transform 1 0 57216 0 1 55278
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_30
timestamp 1621261055
transform -1 0 57504 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output397
timestamp 1621261055
transform -1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_79_591
timestamp 1621261055
transform 1 0 57888 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_159
timestamp 1621261055
transform -1 0 58848 0 1 55278
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_79_595
timestamp 1621261055
transform 1 0 58272 0 1 55278
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output368
timestamp 1621261055
transform 1 0 1536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_160
timestamp 1621261055
transform 1 0 1152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_8
timestamp 1621261055
transform 1 0 1920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output379
timestamp 1621261055
transform 1 0 2304 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_16
timestamp 1621261055
transform 1 0 2688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_56
timestamp 1621261055
transform 1 0 2880 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_24
timestamp 1621261055
transform 1 0 3456 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output417
timestamp 1621261055
transform 1 0 3072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1014
timestamp 1621261055
transform 1 0 3840 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_29
timestamp 1621261055
transform 1 0 3936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_26
timestamp 1621261055
transform 1 0 4128 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output390
timestamp 1621261055
transform 1 0 4320 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_41
timestamp 1621261055
transform 1 0 5088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_37
timestamp 1621261055
transform 1 0 4704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_48
timestamp 1621261055
transform 1 0 5760 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_43
timestamp 1621261055
transform 1 0 5280 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output399
timestamp 1621261055
transform 1 0 5376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_58
timestamp 1621261055
transform 1 0 6720 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_56
timestamp 1621261055
transform 1 0 6528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_32
timestamp 1621261055
transform 1 0 6816 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output437
timestamp 1621261055
transform 1 0 6144 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_65
timestamp 1621261055
transform 1 0 7392 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output400
timestamp 1621261055
transform 1 0 7008 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1015
timestamp 1621261055
transform 1 0 9120 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output401
timestamp 1621261055
transform 1 0 8352 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output402
timestamp 1621261055
transform -1 0 10560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_34
timestamp 1621261055
transform -1 0 10176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_73
timestamp 1621261055
transform 1 0 8160 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_79
timestamp 1621261055
transform 1 0 8736 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_84
timestamp 1621261055
transform 1 0 9216 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_98
timestamp 1621261055
transform 1 0 10560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_90
timestamp 1621261055
transform 1 0 10752 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output440
timestamp 1621261055
transform 1 0 10944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_106
timestamp 1621261055
transform 1 0 11328 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output403
timestamp 1621261055
transform 1 0 11712 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_114
timestamp 1621261055
transform 1 0 12096 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_92
timestamp 1621261055
transform 1 0 12288 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output441
timestamp 1621261055
transform 1 0 12480 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_122
timestamp 1621261055
transform 1 0 12864 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_126
timestamp 1621261055
transform 1 0 13248 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output404
timestamp 1621261055
transform 1 0 13344 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_131
timestamp 1621261055
transform 1 0 13728 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_139
timestamp 1621261055
transform 1 0 14496 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_137
timestamp 1621261055
transform 1 0 14304 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_135
timestamp 1621261055
transform 1 0 14112 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1016
timestamp 1621261055
transform 1 0 14400 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_147
timestamp 1621261055
transform 1 0 15264 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_96
timestamp 1621261055
transform -1 0 15648 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output405
timestamp 1621261055
transform 1 0 14880 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_155
timestamp 1621261055
transform 1 0 16032 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output443
timestamp 1621261055
transform -1 0 16032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_38
timestamp 1621261055
transform -1 0 16992 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output407
timestamp 1621261055
transform -1 0 17376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_169
timestamp 1621261055
transform 1 0 17376 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_173
timestamp 1621261055
transform 1 0 17760 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_1
timestamp 1621261055
transform 1 0 17856 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output370
timestamp 1621261055
transform 1 0 18048 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_180
timestamp 1621261055
transform 1 0 18432 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_40
timestamp 1621261055
transform -1 0 18816 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output408
timestamp 1621261055
transform -1 0 19200 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_188
timestamp 1621261055
transform 1 0 19200 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_192
timestamp 1621261055
transform 1 0 19584 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1017
timestamp 1621261055
transform 1 0 19680 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_194
timestamp 1621261055
transform 1 0 19776 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_3
timestamp 1621261055
transform -1 0 20160 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output371
timestamp 1621261055
transform -1 0 20544 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_206
timestamp 1621261055
transform 1 0 20928 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_202
timestamp 1621261055
transform 1 0 20544 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_213
timestamp 1621261055
transform 1 0 21600 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_42
timestamp 1621261055
transform 1 0 21792 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_5
timestamp 1621261055
transform 1 0 21024 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output372
timestamp 1621261055
transform 1 0 21216 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_221
timestamp 1621261055
transform 1 0 22368 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output410
timestamp 1621261055
transform 1 0 21984 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_229
timestamp 1621261055
transform 1 0 23136 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output373
timestamp 1621261055
transform 1 0 22752 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_237
timestamp 1621261055
transform 1 0 23904 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__diode_2  ANTENNA_7
timestamp 1621261055
transform -1 0 24192 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output374
timestamp 1621261055
transform -1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_244
timestamp 1621261055
transform 1 0 24576 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_249
timestamp 1621261055
transform 1 0 25056 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1018
timestamp 1621261055
transform 1 0 24960 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_80_255
timestamp 1621261055
transform 1 0 25632 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_253
timestamp 1621261055
transform 1 0 25440 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_9
timestamp 1621261055
transform 1 0 25728 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output375
timestamp 1621261055
transform 1 0 25920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_262
timestamp 1621261055
transform 1 0 26304 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_48
timestamp 1621261055
transform -1 0 26688 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output413
timestamp 1621261055
transform -1 0 27072 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_272
timestamp 1621261055
transform 1 0 27264 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_270
timestamp 1621261055
transform 1 0 27072 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_11
timestamp 1621261055
transform -1 0 27552 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output376
timestamp 1621261055
transform -1 0 27936 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_279
timestamp 1621261055
transform 1 0 27936 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_50
timestamp 1621261055
transform -1 0 28320 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output414
timestamp 1621261055
transform -1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_287
timestamp 1621261055
transform 1 0 28704 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_291
timestamp 1621261055
transform 1 0 29088 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_52
timestamp 1621261055
transform -1 0 29472 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output415
timestamp 1621261055
transform -1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_299
timestamp 1621261055
transform 1 0 29856 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_304
timestamp 1621261055
transform 1 0 30336 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1019
timestamp 1621261055
transform 1 0 30240 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output378
timestamp 1621261055
transform 1 0 30720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_312
timestamp 1621261055
transform 1 0 31104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_54
timestamp 1621261055
transform -1 0 31488 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output416
timestamp 1621261055
transform -1 0 31872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_320
timestamp 1621261055
transform 1 0 31872 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_15
timestamp 1621261055
transform 1 0 32064 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output380
timestamp 1621261055
transform 1 0 32256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_328
timestamp 1621261055
transform 1 0 32640 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_58
timestamp 1621261055
transform -1 0 33024 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output418
timestamp 1621261055
transform -1 0 33408 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_336
timestamp 1621261055
transform 1 0 33408 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_344
timestamp 1621261055
transform 1 0 34176 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output381
timestamp 1621261055
transform 1 0 33792 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output419
timestamp 1621261055
transform 1 0 34560 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_352
timestamp 1621261055
transform 1 0 34944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_356
timestamp 1621261055
transform 1 0 35328 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1020
timestamp 1621261055
transform 1 0 35520 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_359
timestamp 1621261055
transform 1 0 35616 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_17
timestamp 1621261055
transform -1 0 36000 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output382
timestamp 1621261055
transform -1 0 36384 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_367
timestamp 1621261055
transform 1 0 36384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_60
timestamp 1621261055
transform -1 0 36768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output420
timestamp 1621261055
transform -1 0 37152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_375
timestamp 1621261055
transform 1 0 37152 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_62
timestamp 1621261055
transform 1 0 37344 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output421
timestamp 1621261055
transform 1 0 37536 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_389
timestamp 1621261055
transform 1 0 38496 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_387
timestamp 1621261055
transform 1 0 38304 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_383
timestamp 1621261055
transform 1 0 37920 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_394
timestamp 1621261055
transform 1 0 38976 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output384
timestamp 1621261055
transform 1 0 38592 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_404
timestamp 1621261055
transform 1 0 39936 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_402
timestamp 1621261055
transform 1 0 39744 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_80_409
timestamp 1621261055
transform 1 0 40416 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output385
timestamp 1621261055
transform 1 0 40032 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1021
timestamp 1621261055
transform 1 0 40800 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_1  FILLER_80_422
timestamp 1621261055
transform 1 0 41664 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_414
timestamp 1621261055
transform 1 0 40896 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_427
timestamp 1621261055
transform 1 0 42144 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_66
timestamp 1621261055
transform -1 0 42528 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output386
timestamp 1621261055
transform 1 0 41760 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_435
timestamp 1621261055
transform 1 0 42912 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_21
timestamp 1621261055
transform -1 0 43296 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output424
timestamp 1621261055
transform -1 0 42912 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_443
timestamp 1621261055
transform 1 0 43680 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output387
timestamp 1621261055
transform -1 0 43680 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_455
timestamp 1621261055
transform 1 0 44832 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_451
timestamp 1621261055
transform 1 0 44448 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output425
timestamp 1621261055
transform 1 0 44064 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_80_460
timestamp 1621261055
transform 1 0 45312 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_2  output388
timestamp 1621261055
transform 1 0 44928 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_469
timestamp 1621261055
transform 1 0 46176 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1022
timestamp 1621261055
transform 1 0 46080 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_80_479
timestamp 1621261055
transform 1 0 47136 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__diode_2  ANTENNA_24
timestamp 1621261055
transform -1 0 47136 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_23
timestamp 1621261055
transform -1 0 46560 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output389
timestamp 1621261055
transform -1 0 46944 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_487
timestamp 1621261055
transform 1 0 47904 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_2  output391
timestamp 1621261055
transform 1 0 48000 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_492
timestamp 1621261055
transform 1 0 48384 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_74
timestamp 1621261055
transform -1 0 48768 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output429
timestamp 1621261055
transform -1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_80_504
timestamp 1621261055
transform 1 0 49536 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_500
timestamp 1621261055
transform 1 0 49152 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_509
timestamp 1621261055
transform 1 0 50016 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output392
timestamp 1621261055
transform 1 0 49632 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output430
timestamp 1621261055
transform 1 0 50400 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_517
timestamp 1621261055
transform 1 0 50784 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_521
timestamp 1621261055
transform 1 0 51168 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1023
timestamp 1621261055
transform 1 0 51360 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_80_524
timestamp 1621261055
transform 1 0 51456 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output393
timestamp 1621261055
transform 1 0 51840 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_532
timestamp 1621261055
transform 1 0 52224 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_536
timestamp 1621261055
transform 1 0 52608 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_542
timestamp 1621261055
transform 1 0 53184 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output394
timestamp 1621261055
transform 1 0 52800 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_77
timestamp 1621261055
transform -1 0 53568 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output432
timestamp 1621261055
transform -1 0 53952 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_550
timestamp 1621261055
transform 1 0 53952 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_28
timestamp 1621261055
transform -1 0 54336 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output395
timestamp 1621261055
transform -1 0 54720 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_558
timestamp 1621261055
transform 1 0 54720 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_79
timestamp 1621261055
transform -1 0 55104 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_568
timestamp 1621261055
transform 1 0 55680 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_80
timestamp 1621261055
transform -1 0 55680 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output433
timestamp 1621261055
transform -1 0 55488 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_80_574
timestamp 1621261055
transform 1 0 56256 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output396
timestamp 1621261055
transform 1 0 55872 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1024
timestamp 1621261055
transform 1 0 56640 0 -1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_80_587
timestamp 1621261055
transform 1 0 57504 0 -1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_80_579
timestamp 1621261055
transform 1 0 56736 0 -1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_80_593
timestamp 1621261055
transform 1 0 58080 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input31
timestamp 1621261055
transform 1 0 57696 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_161
timestamp 1621261055
transform -1 0 58848 0 -1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  PHY_162
timestamp 1621261055
transform 1 0 1152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1025
timestamp 1621261055
transform 1 0 3840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 1536 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input12
timestamp 1621261055
transform 1 0 2400 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_9
timestamp 1621261055
transform 1 0 2016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_18
timestamp 1621261055
transform 1 0 2880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_26
timestamp 1621261055
transform 1 0 3648 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_29
timestamp 1621261055
transform 1 0 3936 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1026
timestamp 1621261055
transform 1 0 6528 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input23
timestamp 1621261055
transform 1 0 5760 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__buf_2  input32
timestamp 1621261055
transform 1 0 4896 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input33
timestamp 1621261055
transform 1 0 7008 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_37
timestamp 1621261055
transform 1 0 4704 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_44
timestamp 1621261055
transform 1 0 5376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_52
timestamp 1621261055
transform 1 0 6144 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_57
timestamp 1621261055
transform 1 0 6624 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_66
timestamp 1621261055
transform 1 0 7488 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1027
timestamp 1621261055
transform 1 0 9216 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input34
timestamp 1621261055
transform 1 0 8064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  input35
timestamp 1621261055
transform 1 0 9696 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_70
timestamp 1621261055
transform 1 0 7872 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_76
timestamp 1621261055
transform 1 0 8448 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_85
timestamp 1621261055
transform 1 0 9312 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_93
timestamp 1621261055
transform 1 0 10080 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1028
timestamp 1621261055
transform 1 0 11904 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input36
timestamp 1621261055
transform 1 0 11040 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input37
timestamp 1621261055
transform 1 0 12768 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_2  output369
timestamp 1621261055
transform 1 0 13824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_101
timestamp 1621261055
transform 1 0 10848 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_108
timestamp 1621261055
transform 1 0 11520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_113
timestamp 1621261055
transform 1 0 12000 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_126
timestamp 1621261055
transform 1 0 13248 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_130
timestamp 1621261055
transform 1 0 13632 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1029
timestamp 1621261055
transform 1 0 14592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input2
timestamp 1621261055
transform 1 0 15936 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input38
timestamp 1621261055
transform 1 0 15072 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_136
timestamp 1621261055
transform 1 0 14208 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_141
timestamp 1621261055
transform 1 0 14688 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_149
timestamp 1621261055
transform 1 0 15456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_153
timestamp 1621261055
transform 1 0 15840 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_159
timestamp 1621261055
transform 1 0 16416 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_169
timestamp 1621261055
transform 1 0 17376 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_167
timestamp 1621261055
transform 1 0 17184 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input3
timestamp 1621261055
transform 1 0 17760 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1030
timestamp 1621261055
transform 1 0 17280 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_178
timestamp 1621261055
transform 1 0 18240 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_186
timestamp 1621261055
transform 1 0 19008 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input4
timestamp 1621261055
transform 1 0 19104 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_197
timestamp 1621261055
transform 1 0 20064 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_192
timestamp 1621261055
transform 1 0 19584 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1031
timestamp 1621261055
transform 1 0 19968 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1032
timestamp 1621261055
transform 1 0 22656 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input5
timestamp 1621261055
transform 1 0 20640 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input6
timestamp 1621261055
transform 1 0 21888 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_201
timestamp 1621261055
transform 1 0 20448 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_8  FILLER_81_208
timestamp 1621261055
transform 1 0 21120 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_220
timestamp 1621261055
transform 1 0 22272 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_225
timestamp 1621261055
transform 1 0 22752 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_235
timestamp 1621261055
transform 1 0 23712 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_233
timestamp 1621261055
transform 1 0 23520 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__buf_2  input7
timestamp 1621261055
transform 1 0 23808 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_8  FILLER_81_241
timestamp 1621261055
transform 1 0 24288 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_253
timestamp 1621261055
transform 1 0 25440 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_251
timestamp 1621261055
transform 1 0 25248 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_249
timestamp 1621261055
transform 1 0 25056 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_1  input8
timestamp 1621261055
transform 1 0 25824 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1033
timestamp 1621261055
transform 1 0 25344 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_261
timestamp 1621261055
transform 1 0 26208 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1034
timestamp 1621261055
transform 1 0 28032 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input9
timestamp 1621261055
transform 1 0 26976 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__buf_2  input10
timestamp 1621261055
transform 1 0 28608 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__decap_4  FILLER_81_274
timestamp 1621261055
transform 1 0 27456 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_278
timestamp 1621261055
transform 1 0 27840 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_281
timestamp 1621261055
transform 1 0 28128 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_285
timestamp 1621261055
transform 1 0 28512 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_291
timestamp 1621261055
transform 1 0 29088 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_304
timestamp 1621261055
transform 1 0 30336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_299
timestamp 1621261055
transform 1 0 29856 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input11
timestamp 1621261055
transform 1 0 29952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_309
timestamp 1621261055
transform 1 0 30816 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1035
timestamp 1621261055
transform 1 0 30720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_322
timestamp 1621261055
transform 1 0 32064 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_317
timestamp 1621261055
transform 1 0 31584 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_1  input13
timestamp 1621261055
transform 1 0 31680 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_330
timestamp 1621261055
transform 1 0 32832 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__diode_2  ANTENNA_13
timestamp 1621261055
transform -1 0 32448 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_2  output377
timestamp 1621261055
transform -1 0 32832 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1036
timestamp 1621261055
transform 1 0 33408 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__buf_2  input14
timestamp 1621261055
transform 1 0 33888 0 1 56610
box -38 -49 518 715
use sky130_fd_sc_ls__clkbuf_1  input15
timestamp 1621261055
transform 1 0 34848 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_334
timestamp 1621261055
transform 1 0 33216 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_337
timestamp 1621261055
transform 1 0 33504 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_346
timestamp 1621261055
transform 1 0 34368 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_350
timestamp 1621261055
transform 1 0 34752 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_355
timestamp 1621261055
transform 1 0 35232 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_363
timestamp 1621261055
transform 1 0 36000 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1037
timestamp 1621261055
transform 1 0 36096 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1038
timestamp 1621261055
transform 1 0 38784 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input16 $PDKPATH/libs.ref/sky130_fd_sc_ls/mag
timestamp 1621261055
transform 1 0 36576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input17
timestamp 1621261055
transform 1 0 38016 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_365
timestamp 1621261055
transform 1 0 36192 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_375
timestamp 1621261055
transform 1 0 37152 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_383
timestamp 1621261055
transform 1 0 37920 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_388
timestamp 1621261055
transform 1 0 38400 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_393
timestamp 1621261055
transform 1 0 38880 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__clkbuf_4  input18
timestamp 1621261055
transform 1 0 39648 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_407
timestamp 1621261055
transform 1 0 40224 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__diode_2  ANTENNA_19
timestamp 1621261055
transform -1 0 40608 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_415
timestamp 1621261055
transform 1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_2  output383
timestamp 1621261055
transform -1 0 40992 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_421
timestamp 1621261055
transform 1 0 41568 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_419
timestamp 1621261055
transform 1 0 41376 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1039
timestamp 1621261055
transform 1 0 41472 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_429
timestamp 1621261055
transform 1 0 42336 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input19
timestamp 1621261055
transform 1 0 41952 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1040
timestamp 1621261055
transform 1 0 44160 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input20
timestamp 1621261055
transform 1 0 42816 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_1  input21
timestamp 1621261055
transform 1 0 44640 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_433
timestamp 1621261055
transform 1 0 42720 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_440
timestamp 1621261055
transform 1 0 43392 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_449
timestamp 1621261055
transform 1 0 44256 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_457
timestamp 1621261055
transform 1 0 45024 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_1  FILLER_81_465
timestamp 1621261055
transform 1 0 45792 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input22
timestamp 1621261055
transform 1 0 45888 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_472
timestamp 1621261055
transform 1 0 46464 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_481
timestamp 1621261055
transform 1 0 47328 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_477
timestamp 1621261055
transform 1 0 46944 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1041
timestamp 1621261055
transform 1 0 46848 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_487
timestamp 1621261055
transform 1 0 47904 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input24
timestamp 1621261055
transform 1 0 47520 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_493
timestamp 1621261055
transform 1 0 48480 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_491
timestamp 1621261055
transform 1 0 48288 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__clkbuf_4  input25
timestamp 1621261055
transform 1 0 48576 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1042
timestamp 1621261055
transform 1 0 49536 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input26
timestamp 1621261055
transform 1 0 50688 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_500
timestamp 1621261055
transform 1 0 49152 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_505
timestamp 1621261055
transform 1 0 49632 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_513
timestamp 1621261055
transform 1 0 50400 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_515
timestamp 1621261055
transform 1 0 50592 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_8  FILLER_81_522
timestamp 1621261055
transform 1 0 51264 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  FILLER_81_533
timestamp 1621261055
transform 1 0 52320 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_530
timestamp 1621261055
transform 1 0 52032 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1043
timestamp 1621261055
transform 1 0 52224 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input27
timestamp 1621261055
transform 1 0 52704 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_547
timestamp 1621261055
transform 1 0 53664 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__decap_4  FILLER_81_543
timestamp 1621261055
transform 1 0 53280 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_553
timestamp 1621261055
transform 1 0 54240 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__clkbuf_1  input28
timestamp 1621261055
transform 1 0 53856 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_4  FILLER_81_561
timestamp 1621261055
transform 1 0 55008 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_1  FILLER_81_559
timestamp 1621261055
transform 1 0 54816 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_557
timestamp 1621261055
transform 1 0 54624 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1044
timestamp 1621261055
transform 1 0 54912 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__tapvpwrvgnd_1  PHY_1045
timestamp 1621261055
transform 1 0 57600 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__clkbuf_4  input29
timestamp 1621261055
transform 1 0 55392 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__clkbuf_4  input30
timestamp 1621261055
transform 1 0 56640 0 1 56610
box -38 -49 614 715
use sky130_fd_sc_ls__decap_4  FILLER_81_571
timestamp 1621261055
transform 1 0 55968 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__fill_diode_2  FILLER_81_575
timestamp 1621261055
transform 1 0 56352 0 1 56610
box -38 -49 230 715
use sky130_fd_sc_ls__fill_1  FILLER_81_577
timestamp 1621261055
transform 1 0 56544 0 1 56610
box -38 -49 134 715
use sky130_fd_sc_ls__decap_4  FILLER_81_584
timestamp 1621261055
transform 1 0 57216 0 1 56610
box -38 -49 422 715
use sky130_fd_sc_ls__decap_8  FILLER_81_589
timestamp 1621261055
transform 1 0 57696 0 1 56610
box -38 -49 806 715
use sky130_fd_sc_ls__decap_4  PHY_163
timestamp 1621261055
transform -1 0 58848 0 1 56610
box -38 -49 422 715
<< labels >>
rlabel metal2 s 212 59200 268 60000 6 io_in[0]
port 0 nsew signal input
rlabel metal2 s 15956 59200 16012 60000 6 io_in[10]
port 1 nsew signal input
rlabel metal2 s 17492 59200 17548 60000 6 io_in[11]
port 2 nsew signal input
rlabel metal2 s 19124 59200 19180 60000 6 io_in[12]
port 3 nsew signal input
rlabel metal2 s 20660 59200 20716 60000 6 io_in[13]
port 4 nsew signal input
rlabel metal2 s 22292 59200 22348 60000 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew signal input
rlabel metal2 s 25460 59200 25516 60000 6 io_in[16]
port 7 nsew signal input
rlabel metal2 s 26996 59200 27052 60000 6 io_in[17]
port 8 nsew signal input
rlabel metal2 s 28628 59200 28684 60000 6 io_in[18]
port 9 nsew signal input
rlabel metal2 s 30164 59200 30220 60000 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew signal input
rlabel metal2 s 31700 59200 31756 60000 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 33332 59200 33388 60000 6 io_in[21]
port 13 nsew signal input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew signal input
rlabel metal2 s 36500 59200 36556 60000 6 io_in[23]
port 15 nsew signal input
rlabel metal2 s 38036 59200 38092 60000 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 39668 59200 39724 60000 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 41204 59200 41260 60000 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 42836 59200 42892 60000 6 io_in[27]
port 19 nsew signal input
rlabel metal2 s 44372 59200 44428 60000 6 io_in[28]
port 20 nsew signal input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew signal input
rlabel metal2 s 3284 59200 3340 60000 6 io_in[2]
port 22 nsew signal input
rlabel metal2 s 47540 59200 47596 60000 6 io_in[30]
port 23 nsew signal input
rlabel metal2 s 49076 59200 49132 60000 6 io_in[31]
port 24 nsew signal input
rlabel metal2 s 50708 59200 50764 60000 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 52244 59200 52300 60000 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 53876 59200 53932 60000 6 io_in[34]
port 27 nsew signal input
rlabel metal2 s 55412 59200 55468 60000 6 io_in[35]
port 28 nsew signal input
rlabel metal2 s 57044 59200 57100 60000 6 io_in[36]
port 29 nsew signal input
rlabel metal2 s 58580 59200 58636 60000 6 io_in[37]
port 30 nsew signal input
rlabel metal2 s 4916 59200 4972 60000 6 io_in[3]
port 31 nsew signal input
rlabel metal2 s 6452 59200 6508 60000 6 io_in[4]
port 32 nsew signal input
rlabel metal2 s 8084 59200 8140 60000 6 io_in[5]
port 33 nsew signal input
rlabel metal2 s 9620 59200 9676 60000 6 io_in[6]
port 34 nsew signal input
rlabel metal2 s 11252 59200 11308 60000 6 io_in[7]
port 35 nsew signal input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew signal input
rlabel metal2 s 14420 59200 14476 60000 6 io_in[9]
port 37 nsew signal input
rlabel metal2 s 692 59200 748 60000 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal2 s 16436 59200 16492 60000 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 18068 59200 18124 60000 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 19604 59200 19660 60000 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 21236 59200 21292 60000 6 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 22772 59200 22828 60000 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal2 s 24404 59200 24460 60000 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 25940 59200 25996 60000 6 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 27572 59200 27628 60000 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 29108 59200 29164 60000 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal2 s 30644 59200 30700 60000 6 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 2228 59200 2284 60000 6 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 32276 59200 32332 60000 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 33812 59200 33868 60000 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal2 s 35444 59200 35500 60000 6 io_oeb[22]
port 52 nsew signal tristate
rlabel metal2 s 36980 59200 37036 60000 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal2 s 38612 59200 38668 60000 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal2 s 40148 59200 40204 60000 6 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 41780 59200 41836 60000 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal2 s 43316 59200 43372 60000 6 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 44948 59200 45004 60000 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal2 s 46484 59200 46540 60000 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal2 s 3860 59200 3916 60000 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 48020 59200 48076 60000 6 io_oeb[30]
port 61 nsew signal tristate
rlabel metal2 s 49652 59200 49708 60000 6 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 51188 59200 51244 60000 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 52820 59200 52876 60000 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 54356 59200 54412 60000 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal2 s 55988 59200 56044 60000 6 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 57524 59200 57580 60000 6 io_oeb[36]
port 67 nsew signal tristate
rlabel metal2 s 59156 59200 59212 60000 6 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 5396 59200 5452 60000 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 7028 59200 7084 60000 6 io_oeb[4]
port 70 nsew signal tristate
rlabel metal2 s 8564 59200 8620 60000 6 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 10196 59200 10252 60000 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 11732 59200 11788 60000 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal2 s 13364 59200 13420 60000 6 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 14900 59200 14956 60000 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 1172 59200 1228 60000 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 17012 59200 17068 60000 6 io_out[10]
port 77 nsew signal tristate
rlabel metal2 s 18548 59200 18604 60000 6 io_out[11]
port 78 nsew signal tristate
rlabel metal2 s 20180 59200 20236 60000 6 io_out[12]
port 79 nsew signal tristate
rlabel metal2 s 21716 59200 21772 60000 6 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 23348 59200 23404 60000 6 io_out[14]
port 81 nsew signal tristate
rlabel metal2 s 24884 59200 24940 60000 6 io_out[15]
port 82 nsew signal tristate
rlabel metal2 s 26516 59200 26572 60000 6 io_out[16]
port 83 nsew signal tristate
rlabel metal2 s 28052 59200 28108 60000 6 io_out[17]
port 84 nsew signal tristate
rlabel metal2 s 29684 59200 29740 60000 6 io_out[18]
port 85 nsew signal tristate
rlabel metal2 s 31220 59200 31276 60000 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 2804 59200 2860 60000 6 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 32756 59200 32812 60000 6 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 34388 59200 34444 60000 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 35924 59200 35980 60000 6 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 37556 59200 37612 60000 6 io_out[23]
port 91 nsew signal tristate
rlabel metal2 s 39092 59200 39148 60000 6 io_out[24]
port 92 nsew signal tristate
rlabel metal2 s 40724 59200 40780 60000 6 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 42260 59200 42316 60000 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 43892 59200 43948 60000 6 io_out[27]
port 95 nsew signal tristate
rlabel metal2 s 45428 59200 45484 60000 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 46964 59200 47020 60000 6 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 4340 59200 4396 60000 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 48596 59200 48652 60000 6 io_out[30]
port 99 nsew signal tristate
rlabel metal2 s 50132 59200 50188 60000 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 51764 59200 51820 60000 6 io_out[32]
port 101 nsew signal tristate
rlabel metal2 s 53300 59200 53356 60000 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 54932 59200 54988 60000 6 io_out[34]
port 103 nsew signal tristate
rlabel metal2 s 56468 59200 56524 60000 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 58100 59200 58156 60000 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 59636 59200 59692 60000 6 io_out[37]
port 106 nsew signal tristate
rlabel metal2 s 5972 59200 6028 60000 6 io_out[3]
port 107 nsew signal tristate
rlabel metal2 s 7508 59200 7564 60000 6 io_out[4]
port 108 nsew signal tristate
rlabel metal2 s 9140 59200 9196 60000 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 10676 59200 10732 60000 6 io_out[6]
port 110 nsew signal tristate
rlabel metal2 s 12308 59200 12364 60000 6 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 13844 59200 13900 60000 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 15380 59200 15436 60000 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 12980 0 13036 800 6 la_data_in[0]
port 114 nsew signal input
rlabel metal2 s 49652 0 49708 800 6 la_data_in[100]
port 115 nsew signal input
rlabel metal2 s 50036 0 50092 800 6 la_data_in[101]
port 116 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[102]
port 117 nsew signal input
rlabel metal2 s 50804 0 50860 800 6 la_data_in[103]
port 118 nsew signal input
rlabel metal2 s 51188 0 51244 800 6 la_data_in[104]
port 119 nsew signal input
rlabel metal2 s 51476 0 51532 800 6 la_data_in[105]
port 120 nsew signal input
rlabel metal2 s 51860 0 51916 800 6 la_data_in[106]
port 121 nsew signal input
rlabel metal2 s 52244 0 52300 800 6 la_data_in[107]
port 122 nsew signal input
rlabel metal2 s 52628 0 52684 800 6 la_data_in[108]
port 123 nsew signal input
rlabel metal2 s 53012 0 53068 800 6 la_data_in[109]
port 124 nsew signal input
rlabel metal2 s 16628 0 16684 800 6 la_data_in[10]
port 125 nsew signal input
rlabel metal2 s 53396 0 53452 800 6 la_data_in[110]
port 126 nsew signal input
rlabel metal2 s 53684 0 53740 800 6 la_data_in[111]
port 127 nsew signal input
rlabel metal2 s 54068 0 54124 800 6 la_data_in[112]
port 128 nsew signal input
rlabel metal2 s 54452 0 54508 800 6 la_data_in[113]
port 129 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[114]
port 130 nsew signal input
rlabel metal2 s 55220 0 55276 800 6 la_data_in[115]
port 131 nsew signal input
rlabel metal2 s 55604 0 55660 800 6 la_data_in[116]
port 132 nsew signal input
rlabel metal2 s 55892 0 55948 800 6 la_data_in[117]
port 133 nsew signal input
rlabel metal2 s 56276 0 56332 800 6 la_data_in[118]
port 134 nsew signal input
rlabel metal2 s 56660 0 56716 800 6 la_data_in[119]
port 135 nsew signal input
rlabel metal2 s 17012 0 17068 800 6 la_data_in[11]
port 136 nsew signal input
rlabel metal2 s 57044 0 57100 800 6 la_data_in[120]
port 137 nsew signal input
rlabel metal2 s 57428 0 57484 800 6 la_data_in[121]
port 138 nsew signal input
rlabel metal2 s 57812 0 57868 800 6 la_data_in[122]
port 139 nsew signal input
rlabel metal2 s 58100 0 58156 800 6 la_data_in[123]
port 140 nsew signal input
rlabel metal2 s 58484 0 58540 800 6 la_data_in[124]
port 141 nsew signal input
rlabel metal2 s 58868 0 58924 800 6 la_data_in[125]
port 142 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[126]
port 143 nsew signal input
rlabel metal2 s 59636 0 59692 800 6 la_data_in[127]
port 144 nsew signal input
rlabel metal2 s 17396 0 17452 800 6 la_data_in[12]
port 145 nsew signal input
rlabel metal2 s 17684 0 17740 800 6 la_data_in[13]
port 146 nsew signal input
rlabel metal2 s 18068 0 18124 800 6 la_data_in[14]
port 147 nsew signal input
rlabel metal2 s 18452 0 18508 800 6 la_data_in[15]
port 148 nsew signal input
rlabel metal2 s 18836 0 18892 800 6 la_data_in[16]
port 149 nsew signal input
rlabel metal2 s 19220 0 19276 800 6 la_data_in[17]
port 150 nsew signal input
rlabel metal2 s 19604 0 19660 800 6 la_data_in[18]
port 151 nsew signal input
rlabel metal2 s 19892 0 19948 800 6 la_data_in[19]
port 152 nsew signal input
rlabel metal2 s 13364 0 13420 800 6 la_data_in[1]
port 153 nsew signal input
rlabel metal2 s 20276 0 20332 800 6 la_data_in[20]
port 154 nsew signal input
rlabel metal2 s 20660 0 20716 800 6 la_data_in[21]
port 155 nsew signal input
rlabel metal2 s 21044 0 21100 800 6 la_data_in[22]
port 156 nsew signal input
rlabel metal2 s 21428 0 21484 800 6 la_data_in[23]
port 157 nsew signal input
rlabel metal2 s 21812 0 21868 800 6 la_data_in[24]
port 158 nsew signal input
rlabel metal2 s 22100 0 22156 800 6 la_data_in[25]
port 159 nsew signal input
rlabel metal2 s 22484 0 22540 800 6 la_data_in[26]
port 160 nsew signal input
rlabel metal2 s 22868 0 22924 800 6 la_data_in[27]
port 161 nsew signal input
rlabel metal2 s 23252 0 23308 800 6 la_data_in[28]
port 162 nsew signal input
rlabel metal2 s 23636 0 23692 800 6 la_data_in[29]
port 163 nsew signal input
rlabel metal2 s 13652 0 13708 800 6 la_data_in[2]
port 164 nsew signal input
rlabel metal2 s 24020 0 24076 800 6 la_data_in[30]
port 165 nsew signal input
rlabel metal2 s 24308 0 24364 800 6 la_data_in[31]
port 166 nsew signal input
rlabel metal2 s 24692 0 24748 800 6 la_data_in[32]
port 167 nsew signal input
rlabel metal2 s 25076 0 25132 800 6 la_data_in[33]
port 168 nsew signal input
rlabel metal2 s 25460 0 25516 800 6 la_data_in[34]
port 169 nsew signal input
rlabel metal2 s 25844 0 25900 800 6 la_data_in[35]
port 170 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_in[36]
port 171 nsew signal input
rlabel metal2 s 26516 0 26572 800 6 la_data_in[37]
port 172 nsew signal input
rlabel metal2 s 26900 0 26956 800 6 la_data_in[38]
port 173 nsew signal input
rlabel metal2 s 27284 0 27340 800 6 la_data_in[39]
port 174 nsew signal input
rlabel metal2 s 14036 0 14092 800 6 la_data_in[3]
port 175 nsew signal input
rlabel metal2 s 27668 0 27724 800 6 la_data_in[40]
port 176 nsew signal input
rlabel metal2 s 28052 0 28108 800 6 la_data_in[41]
port 177 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 la_data_in[42]
port 178 nsew signal input
rlabel metal2 s 28724 0 28780 800 6 la_data_in[43]
port 179 nsew signal input
rlabel metal2 s 29108 0 29164 800 6 la_data_in[44]
port 180 nsew signal input
rlabel metal2 s 29492 0 29548 800 6 la_data_in[45]
port 181 nsew signal input
rlabel metal2 s 29876 0 29932 800 6 la_data_in[46]
port 182 nsew signal input
rlabel metal2 s 30260 0 30316 800 6 la_data_in[47]
port 183 nsew signal input
rlabel metal2 s 30548 0 30604 800 6 la_data_in[48]
port 184 nsew signal input
rlabel metal2 s 30932 0 30988 800 6 la_data_in[49]
port 185 nsew signal input
rlabel metal2 s 14420 0 14476 800 6 la_data_in[4]
port 186 nsew signal input
rlabel metal2 s 31316 0 31372 800 6 la_data_in[50]
port 187 nsew signal input
rlabel metal2 s 31700 0 31756 800 6 la_data_in[51]
port 188 nsew signal input
rlabel metal2 s 32084 0 32140 800 6 la_data_in[52]
port 189 nsew signal input
rlabel metal2 s 32468 0 32524 800 6 la_data_in[53]
port 190 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 la_data_in[54]
port 191 nsew signal input
rlabel metal2 s 33140 0 33196 800 6 la_data_in[55]
port 192 nsew signal input
rlabel metal2 s 33524 0 33580 800 6 la_data_in[56]
port 193 nsew signal input
rlabel metal2 s 33908 0 33964 800 6 la_data_in[57]
port 194 nsew signal input
rlabel metal2 s 34292 0 34348 800 6 la_data_in[58]
port 195 nsew signal input
rlabel metal2 s 34580 0 34636 800 6 la_data_in[59]
port 196 nsew signal input
rlabel metal2 s 14804 0 14860 800 6 la_data_in[5]
port 197 nsew signal input
rlabel metal2 s 34964 0 35020 800 6 la_data_in[60]
port 198 nsew signal input
rlabel metal2 s 35348 0 35404 800 6 la_data_in[61]
port 199 nsew signal input
rlabel metal2 s 35732 0 35788 800 6 la_data_in[62]
port 200 nsew signal input
rlabel metal2 s 36116 0 36172 800 6 la_data_in[63]
port 201 nsew signal input
rlabel metal2 s 36500 0 36556 800 6 la_data_in[64]
port 202 nsew signal input
rlabel metal2 s 36788 0 36844 800 6 la_data_in[65]
port 203 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 la_data_in[66]
port 204 nsew signal input
rlabel metal2 s 37556 0 37612 800 6 la_data_in[67]
port 205 nsew signal input
rlabel metal2 s 37940 0 37996 800 6 la_data_in[68]
port 206 nsew signal input
rlabel metal2 s 38324 0 38380 800 6 la_data_in[69]
port 207 nsew signal input
rlabel metal2 s 15188 0 15244 800 6 la_data_in[6]
port 208 nsew signal input
rlabel metal2 s 38708 0 38764 800 6 la_data_in[70]
port 209 nsew signal input
rlabel metal2 s 38996 0 39052 800 6 la_data_in[71]
port 210 nsew signal input
rlabel metal2 s 39380 0 39436 800 6 la_data_in[72]
port 211 nsew signal input
rlabel metal2 s 39764 0 39820 800 6 la_data_in[73]
port 212 nsew signal input
rlabel metal2 s 40148 0 40204 800 6 la_data_in[74]
port 213 nsew signal input
rlabel metal2 s 40532 0 40588 800 6 la_data_in[75]
port 214 nsew signal input
rlabel metal2 s 40916 0 40972 800 6 la_data_in[76]
port 215 nsew signal input
rlabel metal2 s 41204 0 41260 800 6 la_data_in[77]
port 216 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 la_data_in[78]
port 217 nsew signal input
rlabel metal2 s 41972 0 42028 800 6 la_data_in[79]
port 218 nsew signal input
rlabel metal2 s 15476 0 15532 800 6 la_data_in[7]
port 219 nsew signal input
rlabel metal2 s 42356 0 42412 800 6 la_data_in[80]
port 220 nsew signal input
rlabel metal2 s 42740 0 42796 800 6 la_data_in[81]
port 221 nsew signal input
rlabel metal2 s 43028 0 43084 800 6 la_data_in[82]
port 222 nsew signal input
rlabel metal2 s 43412 0 43468 800 6 la_data_in[83]
port 223 nsew signal input
rlabel metal2 s 43796 0 43852 800 6 la_data_in[84]
port 224 nsew signal input
rlabel metal2 s 44180 0 44236 800 6 la_data_in[85]
port 225 nsew signal input
rlabel metal2 s 44564 0 44620 800 6 la_data_in[86]
port 226 nsew signal input
rlabel metal2 s 44948 0 45004 800 6 la_data_in[87]
port 227 nsew signal input
rlabel metal2 s 45236 0 45292 800 6 la_data_in[88]
port 228 nsew signal input
rlabel metal2 s 45620 0 45676 800 6 la_data_in[89]
port 229 nsew signal input
rlabel metal2 s 15860 0 15916 800 6 la_data_in[8]
port 230 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 la_data_in[90]
port 231 nsew signal input
rlabel metal2 s 46388 0 46444 800 6 la_data_in[91]
port 232 nsew signal input
rlabel metal2 s 46772 0 46828 800 6 la_data_in[92]
port 233 nsew signal input
rlabel metal2 s 47156 0 47212 800 6 la_data_in[93]
port 234 nsew signal input
rlabel metal2 s 47444 0 47500 800 6 la_data_in[94]
port 235 nsew signal input
rlabel metal2 s 47828 0 47884 800 6 la_data_in[95]
port 236 nsew signal input
rlabel metal2 s 48212 0 48268 800 6 la_data_in[96]
port 237 nsew signal input
rlabel metal2 s 48596 0 48652 800 6 la_data_in[97]
port 238 nsew signal input
rlabel metal2 s 48980 0 49036 800 6 la_data_in[98]
port 239 nsew signal input
rlabel metal2 s 49364 0 49420 800 6 la_data_in[99]
port 240 nsew signal input
rlabel metal2 s 16244 0 16300 800 6 la_data_in[9]
port 241 nsew signal input
rlabel metal2 s 13076 0 13132 800 6 la_data_out[0]
port 242 nsew signal tristate
rlabel metal2 s 49844 0 49900 800 6 la_data_out[100]
port 243 nsew signal tristate
rlabel metal2 s 50132 0 50188 800 6 la_data_out[101]
port 244 nsew signal tristate
rlabel metal2 s 50516 0 50572 800 6 la_data_out[102]
port 245 nsew signal tristate
rlabel metal2 s 50900 0 50956 800 6 la_data_out[103]
port 246 nsew signal tristate
rlabel metal2 s 51284 0 51340 800 6 la_data_out[104]
port 247 nsew signal tristate
rlabel metal2 s 51668 0 51724 800 6 la_data_out[105]
port 248 nsew signal tristate
rlabel metal2 s 52052 0 52108 800 6 la_data_out[106]
port 249 nsew signal tristate
rlabel metal2 s 52340 0 52396 800 6 la_data_out[107]
port 250 nsew signal tristate
rlabel metal2 s 52724 0 52780 800 6 la_data_out[108]
port 251 nsew signal tristate
rlabel metal2 s 53108 0 53164 800 6 la_data_out[109]
port 252 nsew signal tristate
rlabel metal2 s 16724 0 16780 800 6 la_data_out[10]
port 253 nsew signal tristate
rlabel metal2 s 53492 0 53548 800 6 la_data_out[110]
port 254 nsew signal tristate
rlabel metal2 s 53876 0 53932 800 6 la_data_out[111]
port 255 nsew signal tristate
rlabel metal2 s 54260 0 54316 800 6 la_data_out[112]
port 256 nsew signal tristate
rlabel metal2 s 54548 0 54604 800 6 la_data_out[113]
port 257 nsew signal tristate
rlabel metal2 s 54932 0 54988 800 6 la_data_out[114]
port 258 nsew signal tristate
rlabel metal2 s 55316 0 55372 800 6 la_data_out[115]
port 259 nsew signal tristate
rlabel metal2 s 55700 0 55756 800 6 la_data_out[116]
port 260 nsew signal tristate
rlabel metal2 s 56084 0 56140 800 6 la_data_out[117]
port 261 nsew signal tristate
rlabel metal2 s 56468 0 56524 800 6 la_data_out[118]
port 262 nsew signal tristate
rlabel metal2 s 56756 0 56812 800 6 la_data_out[119]
port 263 nsew signal tristate
rlabel metal2 s 17108 0 17164 800 6 la_data_out[11]
port 264 nsew signal tristate
rlabel metal2 s 57140 0 57196 800 6 la_data_out[120]
port 265 nsew signal tristate
rlabel metal2 s 57524 0 57580 800 6 la_data_out[121]
port 266 nsew signal tristate
rlabel metal2 s 57908 0 57964 800 6 la_data_out[122]
port 267 nsew signal tristate
rlabel metal2 s 58292 0 58348 800 6 la_data_out[123]
port 268 nsew signal tristate
rlabel metal2 s 58580 0 58636 800 6 la_data_out[124]
port 269 nsew signal tristate
rlabel metal2 s 58964 0 59020 800 6 la_data_out[125]
port 270 nsew signal tristate
rlabel metal2 s 59348 0 59404 800 6 la_data_out[126]
port 271 nsew signal tristate
rlabel metal2 s 59732 0 59788 800 6 la_data_out[127]
port 272 nsew signal tristate
rlabel metal2 s 17492 0 17548 800 6 la_data_out[12]
port 273 nsew signal tristate
rlabel metal2 s 17876 0 17932 800 6 la_data_out[13]
port 274 nsew signal tristate
rlabel metal2 s 18260 0 18316 800 6 la_data_out[14]
port 275 nsew signal tristate
rlabel metal2 s 18548 0 18604 800 6 la_data_out[15]
port 276 nsew signal tristate
rlabel metal2 s 18932 0 18988 800 6 la_data_out[16]
port 277 nsew signal tristate
rlabel metal2 s 19316 0 19372 800 6 la_data_out[17]
port 278 nsew signal tristate
rlabel metal2 s 19700 0 19756 800 6 la_data_out[18]
port 279 nsew signal tristate
rlabel metal2 s 20084 0 20140 800 6 la_data_out[19]
port 280 nsew signal tristate
rlabel metal2 s 13460 0 13516 800 6 la_data_out[1]
port 281 nsew signal tristate
rlabel metal2 s 20468 0 20524 800 6 la_data_out[20]
port 282 nsew signal tristate
rlabel metal2 s 20756 0 20812 800 6 la_data_out[21]
port 283 nsew signal tristate
rlabel metal2 s 21140 0 21196 800 6 la_data_out[22]
port 284 nsew signal tristate
rlabel metal2 s 21524 0 21580 800 6 la_data_out[23]
port 285 nsew signal tristate
rlabel metal2 s 21908 0 21964 800 6 la_data_out[24]
port 286 nsew signal tristate
rlabel metal2 s 22292 0 22348 800 6 la_data_out[25]
port 287 nsew signal tristate
rlabel metal2 s 22580 0 22636 800 6 la_data_out[26]
port 288 nsew signal tristate
rlabel metal2 s 22964 0 23020 800 6 la_data_out[27]
port 289 nsew signal tristate
rlabel metal2 s 23348 0 23404 800 6 la_data_out[28]
port 290 nsew signal tristate
rlabel metal2 s 23732 0 23788 800 6 la_data_out[29]
port 291 nsew signal tristate
rlabel metal2 s 13844 0 13900 800 6 la_data_out[2]
port 292 nsew signal tristate
rlabel metal2 s 24116 0 24172 800 6 la_data_out[30]
port 293 nsew signal tristate
rlabel metal2 s 24500 0 24556 800 6 la_data_out[31]
port 294 nsew signal tristate
rlabel metal2 s 24788 0 24844 800 6 la_data_out[32]
port 295 nsew signal tristate
rlabel metal2 s 25172 0 25228 800 6 la_data_out[33]
port 296 nsew signal tristate
rlabel metal2 s 25556 0 25612 800 6 la_data_out[34]
port 297 nsew signal tristate
rlabel metal2 s 25940 0 25996 800 6 la_data_out[35]
port 298 nsew signal tristate
rlabel metal2 s 26324 0 26380 800 6 la_data_out[36]
port 299 nsew signal tristate
rlabel metal2 s 26708 0 26764 800 6 la_data_out[37]
port 300 nsew signal tristate
rlabel metal2 s 26996 0 27052 800 6 la_data_out[38]
port 301 nsew signal tristate
rlabel metal2 s 27380 0 27436 800 6 la_data_out[39]
port 302 nsew signal tristate
rlabel metal2 s 14132 0 14188 800 6 la_data_out[3]
port 303 nsew signal tristate
rlabel metal2 s 27764 0 27820 800 6 la_data_out[40]
port 304 nsew signal tristate
rlabel metal2 s 28148 0 28204 800 6 la_data_out[41]
port 305 nsew signal tristate
rlabel metal2 s 28532 0 28588 800 6 la_data_out[42]
port 306 nsew signal tristate
rlabel metal2 s 28916 0 28972 800 6 la_data_out[43]
port 307 nsew signal tristate
rlabel metal2 s 29204 0 29260 800 6 la_data_out[44]
port 308 nsew signal tristate
rlabel metal2 s 29588 0 29644 800 6 la_data_out[45]
port 309 nsew signal tristate
rlabel metal2 s 29972 0 30028 800 6 la_data_out[46]
port 310 nsew signal tristate
rlabel metal2 s 30356 0 30412 800 6 la_data_out[47]
port 311 nsew signal tristate
rlabel metal2 s 30740 0 30796 800 6 la_data_out[48]
port 312 nsew signal tristate
rlabel metal2 s 31028 0 31084 800 6 la_data_out[49]
port 313 nsew signal tristate
rlabel metal2 s 14516 0 14572 800 6 la_data_out[4]
port 314 nsew signal tristate
rlabel metal2 s 31412 0 31468 800 6 la_data_out[50]
port 315 nsew signal tristate
rlabel metal2 s 31796 0 31852 800 6 la_data_out[51]
port 316 nsew signal tristate
rlabel metal2 s 32180 0 32236 800 6 la_data_out[52]
port 317 nsew signal tristate
rlabel metal2 s 32564 0 32620 800 6 la_data_out[53]
port 318 nsew signal tristate
rlabel metal2 s 32948 0 33004 800 6 la_data_out[54]
port 319 nsew signal tristate
rlabel metal2 s 33236 0 33292 800 6 la_data_out[55]
port 320 nsew signal tristate
rlabel metal2 s 33620 0 33676 800 6 la_data_out[56]
port 321 nsew signal tristate
rlabel metal2 s 34004 0 34060 800 6 la_data_out[57]
port 322 nsew signal tristate
rlabel metal2 s 34388 0 34444 800 6 la_data_out[58]
port 323 nsew signal tristate
rlabel metal2 s 34772 0 34828 800 6 la_data_out[59]
port 324 nsew signal tristate
rlabel metal2 s 14900 0 14956 800 6 la_data_out[5]
port 325 nsew signal tristate
rlabel metal2 s 35156 0 35212 800 6 la_data_out[60]
port 326 nsew signal tristate
rlabel metal2 s 35444 0 35500 800 6 la_data_out[61]
port 327 nsew signal tristate
rlabel metal2 s 35828 0 35884 800 6 la_data_out[62]
port 328 nsew signal tristate
rlabel metal2 s 36212 0 36268 800 6 la_data_out[63]
port 329 nsew signal tristate
rlabel metal2 s 36596 0 36652 800 6 la_data_out[64]
port 330 nsew signal tristate
rlabel metal2 s 36980 0 37036 800 6 la_data_out[65]
port 331 nsew signal tristate
rlabel metal2 s 37364 0 37420 800 6 la_data_out[66]
port 332 nsew signal tristate
rlabel metal2 s 37652 0 37708 800 6 la_data_out[67]
port 333 nsew signal tristate
rlabel metal2 s 38036 0 38092 800 6 la_data_out[68]
port 334 nsew signal tristate
rlabel metal2 s 38420 0 38476 800 6 la_data_out[69]
port 335 nsew signal tristate
rlabel metal2 s 15284 0 15340 800 6 la_data_out[6]
port 336 nsew signal tristate
rlabel metal2 s 38804 0 38860 800 6 la_data_out[70]
port 337 nsew signal tristate
rlabel metal2 s 39188 0 39244 800 6 la_data_out[71]
port 338 nsew signal tristate
rlabel metal2 s 39476 0 39532 800 6 la_data_out[72]
port 339 nsew signal tristate
rlabel metal2 s 39860 0 39916 800 6 la_data_out[73]
port 340 nsew signal tristate
rlabel metal2 s 40244 0 40300 800 6 la_data_out[74]
port 341 nsew signal tristate
rlabel metal2 s 40628 0 40684 800 6 la_data_out[75]
port 342 nsew signal tristate
rlabel metal2 s 41012 0 41068 800 6 la_data_out[76]
port 343 nsew signal tristate
rlabel metal2 s 41396 0 41452 800 6 la_data_out[77]
port 344 nsew signal tristate
rlabel metal2 s 41684 0 41740 800 6 la_data_out[78]
port 345 nsew signal tristate
rlabel metal2 s 42068 0 42124 800 6 la_data_out[79]
port 346 nsew signal tristate
rlabel metal2 s 15668 0 15724 800 6 la_data_out[7]
port 347 nsew signal tristate
rlabel metal2 s 42452 0 42508 800 6 la_data_out[80]
port 348 nsew signal tristate
rlabel metal2 s 42836 0 42892 800 6 la_data_out[81]
port 349 nsew signal tristate
rlabel metal2 s 43220 0 43276 800 6 la_data_out[82]
port 350 nsew signal tristate
rlabel metal2 s 43604 0 43660 800 6 la_data_out[83]
port 351 nsew signal tristate
rlabel metal2 s 43892 0 43948 800 6 la_data_out[84]
port 352 nsew signal tristate
rlabel metal2 s 44276 0 44332 800 6 la_data_out[85]
port 353 nsew signal tristate
rlabel metal2 s 44660 0 44716 800 6 la_data_out[86]
port 354 nsew signal tristate
rlabel metal2 s 45044 0 45100 800 6 la_data_out[87]
port 355 nsew signal tristate
rlabel metal2 s 45428 0 45484 800 6 la_data_out[88]
port 356 nsew signal tristate
rlabel metal2 s 45812 0 45868 800 6 la_data_out[89]
port 357 nsew signal tristate
rlabel metal2 s 16052 0 16108 800 6 la_data_out[8]
port 358 nsew signal tristate
rlabel metal2 s 46100 0 46156 800 6 la_data_out[90]
port 359 nsew signal tristate
rlabel metal2 s 46484 0 46540 800 6 la_data_out[91]
port 360 nsew signal tristate
rlabel metal2 s 46868 0 46924 800 6 la_data_out[92]
port 361 nsew signal tristate
rlabel metal2 s 47252 0 47308 800 6 la_data_out[93]
port 362 nsew signal tristate
rlabel metal2 s 47636 0 47692 800 6 la_data_out[94]
port 363 nsew signal tristate
rlabel metal2 s 48020 0 48076 800 6 la_data_out[95]
port 364 nsew signal tristate
rlabel metal2 s 48308 0 48364 800 6 la_data_out[96]
port 365 nsew signal tristate
rlabel metal2 s 48692 0 48748 800 6 la_data_out[97]
port 366 nsew signal tristate
rlabel metal2 s 49076 0 49132 800 6 la_data_out[98]
port 367 nsew signal tristate
rlabel metal2 s 49460 0 49516 800 6 la_data_out[99]
port 368 nsew signal tristate
rlabel metal2 s 16340 0 16396 800 6 la_data_out[9]
port 369 nsew signal tristate
rlabel metal2 s 13172 0 13228 800 6 la_oen[0]
port 370 nsew signal input
rlabel metal2 s 49940 0 49996 800 6 la_oen[100]
port 371 nsew signal input
rlabel metal2 s 50324 0 50380 800 6 la_oen[101]
port 372 nsew signal input
rlabel metal2 s 50708 0 50764 800 6 la_oen[102]
port 373 nsew signal input
rlabel metal2 s 50996 0 51052 800 6 la_oen[103]
port 374 nsew signal input
rlabel metal2 s 51380 0 51436 800 6 la_oen[104]
port 375 nsew signal input
rlabel metal2 s 51764 0 51820 800 6 la_oen[105]
port 376 nsew signal input
rlabel metal2 s 52148 0 52204 800 6 la_oen[106]
port 377 nsew signal input
rlabel metal2 s 52532 0 52588 800 6 la_oen[107]
port 378 nsew signal input
rlabel metal2 s 52916 0 52972 800 6 la_oen[108]
port 379 nsew signal input
rlabel metal2 s 53204 0 53260 800 6 la_oen[109]
port 380 nsew signal input
rlabel metal2 s 16916 0 16972 800 6 la_oen[10]
port 381 nsew signal input
rlabel metal2 s 53588 0 53644 800 6 la_oen[110]
port 382 nsew signal input
rlabel metal2 s 53972 0 54028 800 6 la_oen[111]
port 383 nsew signal input
rlabel metal2 s 54356 0 54412 800 6 la_oen[112]
port 384 nsew signal input
rlabel metal2 s 54740 0 54796 800 6 la_oen[113]
port 385 nsew signal input
rlabel metal2 s 55028 0 55084 800 6 la_oen[114]
port 386 nsew signal input
rlabel metal2 s 55412 0 55468 800 6 la_oen[115]
port 387 nsew signal input
rlabel metal2 s 55796 0 55852 800 6 la_oen[116]
port 388 nsew signal input
rlabel metal2 s 56180 0 56236 800 6 la_oen[117]
port 389 nsew signal input
rlabel metal2 s 56564 0 56620 800 6 la_oen[118]
port 390 nsew signal input
rlabel metal2 s 56948 0 57004 800 6 la_oen[119]
port 391 nsew signal input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew signal input
rlabel metal2 s 57236 0 57292 800 6 la_oen[120]
port 393 nsew signal input
rlabel metal2 s 57620 0 57676 800 6 la_oen[121]
port 394 nsew signal input
rlabel metal2 s 58004 0 58060 800 6 la_oen[122]
port 395 nsew signal input
rlabel metal2 s 58388 0 58444 800 6 la_oen[123]
port 396 nsew signal input
rlabel metal2 s 58772 0 58828 800 6 la_oen[124]
port 397 nsew signal input
rlabel metal2 s 59156 0 59212 800 6 la_oen[125]
port 398 nsew signal input
rlabel metal2 s 59444 0 59500 800 6 la_oen[126]
port 399 nsew signal input
rlabel metal2 s 59828 0 59884 800 6 la_oen[127]
port 400 nsew signal input
rlabel metal2 s 17588 0 17644 800 6 la_oen[12]
port 401 nsew signal input
rlabel metal2 s 17972 0 18028 800 6 la_oen[13]
port 402 nsew signal input
rlabel metal2 s 18356 0 18412 800 6 la_oen[14]
port 403 nsew signal input
rlabel metal2 s 18740 0 18796 800 6 la_oen[15]
port 404 nsew signal input
rlabel metal2 s 19028 0 19084 800 6 la_oen[16]
port 405 nsew signal input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew signal input
rlabel metal2 s 19796 0 19852 800 6 la_oen[18]
port 407 nsew signal input
rlabel metal2 s 20180 0 20236 800 6 la_oen[19]
port 408 nsew signal input
rlabel metal2 s 13556 0 13612 800 6 la_oen[1]
port 409 nsew signal input
rlabel metal2 s 20564 0 20620 800 6 la_oen[20]
port 410 nsew signal input
rlabel metal2 s 20948 0 21004 800 6 la_oen[21]
port 411 nsew signal input
rlabel metal2 s 21236 0 21292 800 6 la_oen[22]
port 412 nsew signal input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew signal input
rlabel metal2 s 22004 0 22060 800 6 la_oen[24]
port 414 nsew signal input
rlabel metal2 s 22388 0 22444 800 6 la_oen[25]
port 415 nsew signal input
rlabel metal2 s 22772 0 22828 800 6 la_oen[26]
port 416 nsew signal input
rlabel metal2 s 23156 0 23212 800 6 la_oen[27]
port 417 nsew signal input
rlabel metal2 s 23444 0 23500 800 6 la_oen[28]
port 418 nsew signal input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew signal input
rlabel metal2 s 13940 0 13996 800 6 la_oen[2]
port 420 nsew signal input
rlabel metal2 s 24212 0 24268 800 6 la_oen[30]
port 421 nsew signal input
rlabel metal2 s 24596 0 24652 800 6 la_oen[31]
port 422 nsew signal input
rlabel metal2 s 24980 0 25036 800 6 la_oen[32]
port 423 nsew signal input
rlabel metal2 s 25364 0 25420 800 6 la_oen[33]
port 424 nsew signal input
rlabel metal2 s 25652 0 25708 800 6 la_oen[34]
port 425 nsew signal input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew signal input
rlabel metal2 s 26420 0 26476 800 6 la_oen[36]
port 427 nsew signal input
rlabel metal2 s 26804 0 26860 800 6 la_oen[37]
port 428 nsew signal input
rlabel metal2 s 27188 0 27244 800 6 la_oen[38]
port 429 nsew signal input
rlabel metal2 s 27476 0 27532 800 6 la_oen[39]
port 430 nsew signal input
rlabel metal2 s 14324 0 14380 800 6 la_oen[3]
port 431 nsew signal input
rlabel metal2 s 27860 0 27916 800 6 la_oen[40]
port 432 nsew signal input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew signal input
rlabel metal2 s 28628 0 28684 800 6 la_oen[42]
port 434 nsew signal input
rlabel metal2 s 29012 0 29068 800 6 la_oen[43]
port 435 nsew signal input
rlabel metal2 s 29396 0 29452 800 6 la_oen[44]
port 436 nsew signal input
rlabel metal2 s 29684 0 29740 800 6 la_oen[45]
port 437 nsew signal input
rlabel metal2 s 30068 0 30124 800 6 la_oen[46]
port 438 nsew signal input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew signal input
rlabel metal2 s 30836 0 30892 800 6 la_oen[48]
port 440 nsew signal input
rlabel metal2 s 31220 0 31276 800 6 la_oen[49]
port 441 nsew signal input
rlabel metal2 s 14708 0 14764 800 6 la_oen[4]
port 442 nsew signal input
rlabel metal2 s 31604 0 31660 800 6 la_oen[50]
port 443 nsew signal input
rlabel metal2 s 31892 0 31948 800 6 la_oen[51]
port 444 nsew signal input
rlabel metal2 s 32276 0 32332 800 6 la_oen[52]
port 445 nsew signal input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew signal input
rlabel metal2 s 33044 0 33100 800 6 la_oen[54]
port 447 nsew signal input
rlabel metal2 s 33428 0 33484 800 6 la_oen[55]
port 448 nsew signal input
rlabel metal2 s 33812 0 33868 800 6 la_oen[56]
port 449 nsew signal input
rlabel metal2 s 34100 0 34156 800 6 la_oen[57]
port 450 nsew signal input
rlabel metal2 s 34484 0 34540 800 6 la_oen[58]
port 451 nsew signal input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew signal input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew signal input
rlabel metal2 s 35252 0 35308 800 6 la_oen[60]
port 454 nsew signal input
rlabel metal2 s 35636 0 35692 800 6 la_oen[61]
port 455 nsew signal input
rlabel metal2 s 36020 0 36076 800 6 la_oen[62]
port 456 nsew signal input
rlabel metal2 s 36308 0 36364 800 6 la_oen[63]
port 457 nsew signal input
rlabel metal2 s 36692 0 36748 800 6 la_oen[64]
port 458 nsew signal input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew signal input
rlabel metal2 s 37460 0 37516 800 6 la_oen[66]
port 460 nsew signal input
rlabel metal2 s 37844 0 37900 800 6 la_oen[67]
port 461 nsew signal input
rlabel metal2 s 38132 0 38188 800 6 la_oen[68]
port 462 nsew signal input
rlabel metal2 s 38516 0 38572 800 6 la_oen[69]
port 463 nsew signal input
rlabel metal2 s 15380 0 15436 800 6 la_oen[6]
port 464 nsew signal input
rlabel metal2 s 38900 0 38956 800 6 la_oen[70]
port 465 nsew signal input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew signal input
rlabel metal2 s 39668 0 39724 800 6 la_oen[72]
port 467 nsew signal input
rlabel metal2 s 40052 0 40108 800 6 la_oen[73]
port 468 nsew signal input
rlabel metal2 s 40340 0 40396 800 6 la_oen[74]
port 469 nsew signal input
rlabel metal2 s 40724 0 40780 800 6 la_oen[75]
port 470 nsew signal input
rlabel metal2 s 41108 0 41164 800 6 la_oen[76]
port 471 nsew signal input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew signal input
rlabel metal2 s 41876 0 41932 800 6 la_oen[78]
port 473 nsew signal input
rlabel metal2 s 42260 0 42316 800 6 la_oen[79]
port 474 nsew signal input
rlabel metal2 s 15764 0 15820 800 6 la_oen[7]
port 475 nsew signal input
rlabel metal2 s 42548 0 42604 800 6 la_oen[80]
port 476 nsew signal input
rlabel metal2 s 42932 0 42988 800 6 la_oen[81]
port 477 nsew signal input
rlabel metal2 s 43316 0 43372 800 6 la_oen[82]
port 478 nsew signal input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew signal input
rlabel metal2 s 44084 0 44140 800 6 la_oen[84]
port 480 nsew signal input
rlabel metal2 s 44468 0 44524 800 6 la_oen[85]
port 481 nsew signal input
rlabel metal2 s 44756 0 44812 800 6 la_oen[86]
port 482 nsew signal input
rlabel metal2 s 45140 0 45196 800 6 la_oen[87]
port 483 nsew signal input
rlabel metal2 s 45524 0 45580 800 6 la_oen[88]
port 484 nsew signal input
rlabel metal2 s 45908 0 45964 800 6 la_oen[89]
port 485 nsew signal input
rlabel metal2 s 16148 0 16204 800 6 la_oen[8]
port 486 nsew signal input
rlabel metal2 s 46292 0 46348 800 6 la_oen[90]
port 487 nsew signal input
rlabel metal2 s 46580 0 46636 800 6 la_oen[91]
port 488 nsew signal input
rlabel metal2 s 46964 0 47020 800 6 la_oen[92]
port 489 nsew signal input
rlabel metal2 s 47348 0 47404 800 6 la_oen[93]
port 490 nsew signal input
rlabel metal2 s 47732 0 47788 800 6 la_oen[94]
port 491 nsew signal input
rlabel metal2 s 48116 0 48172 800 6 la_oen[95]
port 492 nsew signal input
rlabel metal2 s 48500 0 48556 800 6 la_oen[96]
port 493 nsew signal input
rlabel metal2 s 48788 0 48844 800 6 la_oen[97]
port 494 nsew signal input
rlabel metal2 s 49172 0 49228 800 6 la_oen[98]
port 495 nsew signal input
rlabel metal2 s 49556 0 49612 800 6 la_oen[99]
port 496 nsew signal input
rlabel metal2 s 16532 0 16588 800 6 la_oen[9]
port 497 nsew signal input
rlabel metal2 s 20 0 76 800 6 wb_clk_i
port 498 nsew signal input
rlabel metal2 s 116 0 172 800 6 wb_rst_i
port 499 nsew signal input
rlabel metal2 s 212 0 268 800 6 wbs_ack_o
port 500 nsew signal tristate
rlabel metal2 s 692 0 748 800 6 wbs_adr_i[0]
port 501 nsew signal input
rlabel metal2 s 4916 0 4972 800 6 wbs_adr_i[10]
port 502 nsew signal input
rlabel metal2 s 5204 0 5260 800 6 wbs_adr_i[11]
port 503 nsew signal input
rlabel metal2 s 5588 0 5644 800 6 wbs_adr_i[12]
port 504 nsew signal input
rlabel metal2 s 5972 0 6028 800 6 wbs_adr_i[13]
port 505 nsew signal input
rlabel metal2 s 6356 0 6412 800 6 wbs_adr_i[14]
port 506 nsew signal input
rlabel metal2 s 6740 0 6796 800 6 wbs_adr_i[15]
port 507 nsew signal input
rlabel metal2 s 7028 0 7084 800 6 wbs_adr_i[16]
port 508 nsew signal input
rlabel metal2 s 7412 0 7468 800 6 wbs_adr_i[17]
port 509 nsew signal input
rlabel metal2 s 7796 0 7852 800 6 wbs_adr_i[18]
port 510 nsew signal input
rlabel metal2 s 8180 0 8236 800 6 wbs_adr_i[19]
port 511 nsew signal input
rlabel metal2 s 1172 0 1228 800 6 wbs_adr_i[1]
port 512 nsew signal input
rlabel metal2 s 8564 0 8620 800 6 wbs_adr_i[20]
port 513 nsew signal input
rlabel metal2 s 8948 0 9004 800 6 wbs_adr_i[21]
port 514 nsew signal input
rlabel metal2 s 9236 0 9292 800 6 wbs_adr_i[22]
port 515 nsew signal input
rlabel metal2 s 9620 0 9676 800 6 wbs_adr_i[23]
port 516 nsew signal input
rlabel metal2 s 10004 0 10060 800 6 wbs_adr_i[24]
port 517 nsew signal input
rlabel metal2 s 10388 0 10444 800 6 wbs_adr_i[25]
port 518 nsew signal input
rlabel metal2 s 10772 0 10828 800 6 wbs_adr_i[26]
port 519 nsew signal input
rlabel metal2 s 11156 0 11212 800 6 wbs_adr_i[27]
port 520 nsew signal input
rlabel metal2 s 11444 0 11500 800 6 wbs_adr_i[28]
port 521 nsew signal input
rlabel metal2 s 11828 0 11884 800 6 wbs_adr_i[29]
port 522 nsew signal input
rlabel metal2 s 1652 0 1708 800 6 wbs_adr_i[2]
port 523 nsew signal input
rlabel metal2 s 12212 0 12268 800 6 wbs_adr_i[30]
port 524 nsew signal input
rlabel metal2 s 12596 0 12652 800 6 wbs_adr_i[31]
port 525 nsew signal input
rlabel metal2 s 2132 0 2188 800 6 wbs_adr_i[3]
port 526 nsew signal input
rlabel metal2 s 2708 0 2764 800 6 wbs_adr_i[4]
port 527 nsew signal input
rlabel metal2 s 2996 0 3052 800 6 wbs_adr_i[5]
port 528 nsew signal input
rlabel metal2 s 3380 0 3436 800 6 wbs_adr_i[6]
port 529 nsew signal input
rlabel metal2 s 3764 0 3820 800 6 wbs_adr_i[7]
port 530 nsew signal input
rlabel metal2 s 4148 0 4204 800 6 wbs_adr_i[8]
port 531 nsew signal input
rlabel metal2 s 4532 0 4588 800 6 wbs_adr_i[9]
port 532 nsew signal input
rlabel metal2 s 308 0 364 800 6 wbs_cyc_i
port 533 nsew signal input
rlabel metal2 s 788 0 844 800 6 wbs_dat_i[0]
port 534 nsew signal input
rlabel metal2 s 5012 0 5068 800 6 wbs_dat_i[10]
port 535 nsew signal input
rlabel metal2 s 5396 0 5452 800 6 wbs_dat_i[11]
port 536 nsew signal input
rlabel metal2 s 5684 0 5740 800 6 wbs_dat_i[12]
port 537 nsew signal input
rlabel metal2 s 6068 0 6124 800 6 wbs_dat_i[13]
port 538 nsew signal input
rlabel metal2 s 6452 0 6508 800 6 wbs_dat_i[14]
port 539 nsew signal input
rlabel metal2 s 6836 0 6892 800 6 wbs_dat_i[15]
port 540 nsew signal input
rlabel metal2 s 7220 0 7276 800 6 wbs_dat_i[16]
port 541 nsew signal input
rlabel metal2 s 7604 0 7660 800 6 wbs_dat_i[17]
port 542 nsew signal input
rlabel metal2 s 7892 0 7948 800 6 wbs_dat_i[18]
port 543 nsew signal input
rlabel metal2 s 8276 0 8332 800 6 wbs_dat_i[19]
port 544 nsew signal input
rlabel metal2 s 1364 0 1420 800 6 wbs_dat_i[1]
port 545 nsew signal input
rlabel metal2 s 8660 0 8716 800 6 wbs_dat_i[20]
port 546 nsew signal input
rlabel metal2 s 9044 0 9100 800 6 wbs_dat_i[21]
port 547 nsew signal input
rlabel metal2 s 9428 0 9484 800 6 wbs_dat_i[22]
port 548 nsew signal input
rlabel metal2 s 9812 0 9868 800 6 wbs_dat_i[23]
port 549 nsew signal input
rlabel metal2 s 10100 0 10156 800 6 wbs_dat_i[24]
port 550 nsew signal input
rlabel metal2 s 10484 0 10540 800 6 wbs_dat_i[25]
port 551 nsew signal input
rlabel metal2 s 10868 0 10924 800 6 wbs_dat_i[26]
port 552 nsew signal input
rlabel metal2 s 11252 0 11308 800 6 wbs_dat_i[27]
port 553 nsew signal input
rlabel metal2 s 11636 0 11692 800 6 wbs_dat_i[28]
port 554 nsew signal input
rlabel metal2 s 12020 0 12076 800 6 wbs_dat_i[29]
port 555 nsew signal input
rlabel metal2 s 1844 0 1900 800 6 wbs_dat_i[2]
port 556 nsew signal input
rlabel metal2 s 12308 0 12364 800 6 wbs_dat_i[30]
port 557 nsew signal input
rlabel metal2 s 12692 0 12748 800 6 wbs_dat_i[31]
port 558 nsew signal input
rlabel metal2 s 2324 0 2380 800 6 wbs_dat_i[3]
port 559 nsew signal input
rlabel metal2 s 2804 0 2860 800 6 wbs_dat_i[4]
port 560 nsew signal input
rlabel metal2 s 3188 0 3244 800 6 wbs_dat_i[5]
port 561 nsew signal input
rlabel metal2 s 3476 0 3532 800 6 wbs_dat_i[6]
port 562 nsew signal input
rlabel metal2 s 3860 0 3916 800 6 wbs_dat_i[7]
port 563 nsew signal input
rlabel metal2 s 4244 0 4300 800 6 wbs_dat_i[8]
port 564 nsew signal input
rlabel metal2 s 4628 0 4684 800 6 wbs_dat_i[9]
port 565 nsew signal input
rlabel metal2 s 980 0 1036 800 6 wbs_dat_o[0]
port 566 nsew signal tristate
rlabel metal2 s 5108 0 5164 800 6 wbs_dat_o[10]
port 567 nsew signal tristate
rlabel metal2 s 5492 0 5548 800 6 wbs_dat_o[11]
port 568 nsew signal tristate
rlabel metal2 s 5876 0 5932 800 6 wbs_dat_o[12]
port 569 nsew signal tristate
rlabel metal2 s 6260 0 6316 800 6 wbs_dat_o[13]
port 570 nsew signal tristate
rlabel metal2 s 6548 0 6604 800 6 wbs_dat_o[14]
port 571 nsew signal tristate
rlabel metal2 s 6932 0 6988 800 6 wbs_dat_o[15]
port 572 nsew signal tristate
rlabel metal2 s 7316 0 7372 800 6 wbs_dat_o[16]
port 573 nsew signal tristate
rlabel metal2 s 7700 0 7756 800 6 wbs_dat_o[17]
port 574 nsew signal tristate
rlabel metal2 s 8084 0 8140 800 6 wbs_dat_o[18]
port 575 nsew signal tristate
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_o[19]
port 576 nsew signal tristate
rlabel metal2 s 1460 0 1516 800 6 wbs_dat_o[1]
port 577 nsew signal tristate
rlabel metal2 s 8756 0 8812 800 6 wbs_dat_o[20]
port 578 nsew signal tristate
rlabel metal2 s 9140 0 9196 800 6 wbs_dat_o[21]
port 579 nsew signal tristate
rlabel metal2 s 9524 0 9580 800 6 wbs_dat_o[22]
port 580 nsew signal tristate
rlabel metal2 s 9908 0 9964 800 6 wbs_dat_o[23]
port 581 nsew signal tristate
rlabel metal2 s 10292 0 10348 800 6 wbs_dat_o[24]
port 582 nsew signal tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew signal tristate
rlabel metal2 s 10964 0 11020 800 6 wbs_dat_o[26]
port 584 nsew signal tristate
rlabel metal2 s 11348 0 11404 800 6 wbs_dat_o[27]
port 585 nsew signal tristate
rlabel metal2 s 11732 0 11788 800 6 wbs_dat_o[28]
port 586 nsew signal tristate
rlabel metal2 s 12116 0 12172 800 6 wbs_dat_o[29]
port 587 nsew signal tristate
rlabel metal2 s 1940 0 1996 800 6 wbs_dat_o[2]
port 588 nsew signal tristate
rlabel metal2 s 12500 0 12556 800 6 wbs_dat_o[30]
port 589 nsew signal tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew signal tristate
rlabel metal2 s 2420 0 2476 800 6 wbs_dat_o[3]
port 591 nsew signal tristate
rlabel metal2 s 2900 0 2956 800 6 wbs_dat_o[4]
port 592 nsew signal tristate
rlabel metal2 s 3284 0 3340 800 6 wbs_dat_o[5]
port 593 nsew signal tristate
rlabel metal2 s 3668 0 3724 800 6 wbs_dat_o[6]
port 594 nsew signal tristate
rlabel metal2 s 4052 0 4108 800 6 wbs_dat_o[7]
port 595 nsew signal tristate
rlabel metal2 s 4340 0 4396 800 6 wbs_dat_o[8]
port 596 nsew signal tristate
rlabel metal2 s 4724 0 4780 800 6 wbs_dat_o[9]
port 597 nsew signal tristate
rlabel metal2 s 1076 0 1132 800 6 wbs_sel_i[0]
port 598 nsew signal input
rlabel metal2 s 1556 0 1612 800 6 wbs_sel_i[1]
port 599 nsew signal input
rlabel metal2 s 2036 0 2092 800 6 wbs_sel_i[2]
port 600 nsew signal input
rlabel metal2 s 2516 0 2572 800 6 wbs_sel_i[3]
port 601 nsew signal input
rlabel metal2 s 500 0 556 800 6 wbs_stb_i
port 602 nsew signal input
rlabel metal2 s 596 0 652 800 6 wbs_we_i
port 603 nsew signal input
rlabel metal4 s 34976 2616 35296 57324 6 vccd1
port 604 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 57324 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 50336 2616 50656 57324 6 vssd1
port 606 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 57324 6 vssd1
port 607 nsew ground bidirectional
rlabel metal4 s 35636 2664 35956 57276 6 vccd2
port 608 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 57276 6 vccd2
port 609 nsew power bidirectional
rlabel metal4 s 50996 2664 51316 57276 6 vssd2
port 610 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 57276 6 vssd2
port 611 nsew ground bidirectional
rlabel metal4 s 36296 2664 36616 57276 6 vdda1
port 612 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 57276 6 vdda1
port 613 nsew power bidirectional
rlabel metal4 s 51656 2664 51976 57276 6 vssa1
port 614 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 57276 6 vssa1
port 615 nsew ground bidirectional
rlabel metal4 s 36956 2664 37276 57276 6 vdda2
port 616 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 57276 6 vdda2
port 617 nsew power bidirectional
rlabel metal4 s 52316 2664 52636 57276 6 vssa2
port 618 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 57276 6 vssa2
port 619 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
