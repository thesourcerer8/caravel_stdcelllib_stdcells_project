MACRO NOR2X1
 CLASS CORE ;
 FOREIGN NOR2X1 0 0 ;
 SIZE 4.32 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 4.32000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 4.32000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.81500000 0.44000000 1.10500000 0.51500000 ;
        RECT 3.21500000 0.44000000 3.50500000 0.51500000 ;
        RECT 0.81500000 0.51500000 3.50500000 0.65500000 ;
        RECT 0.81500000 0.65500000 1.10500000 0.73000000 ;
        RECT 3.21500000 0.65500000 3.50500000 0.73000000 ;
        RECT 3.29000000 0.73000000 3.43000000 2.19500000 ;
        RECT 3.21500000 2.19500000 3.50500000 2.48500000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
        RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
        RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 3.27500000 2.25500000 3.44500000 2.42500000 ;
     RECT 0.63500000 2.84000000 0.80500000 3.01000000 ;

    LAYER ndiffc ;
     RECT 1.83500000 0.32000000 2.00500000 0.49000000 ;
     RECT 0.87500000 0.50000000 1.04500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;

    LAYER li1 ;
     RECT 1.83500000 0.09500000 2.00500000 0.24000000 ;
     RECT 1.75500000 0.24000000 2.08500000 0.57000000 ;
     RECT 0.79500000 0.42000000 1.12500000 0.75000000 ;
     RECT 3.19500000 0.42000000 3.52500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 3.19500000 2.17500000 3.52500000 2.50500000 ;
     RECT 0.55500000 2.76000000 0.88500000 3.09000000 ;

    LAYER viali ;
     RECT 1.83500000 0.09500000 2.00500000 0.26500000 ;
     RECT 0.87500000 0.50000000 1.04500000 0.67000000 ;
     RECT 3.27500000 0.50000000 3.44500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 3.27500000 2.25500000 3.44500000 2.42500000 ;
     RECT 0.63500000 2.84000000 0.80500000 3.01000000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 4.32000000 0.24000000 ;
     RECT 1.77500000 0.24000000 2.06500000 0.32500000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
     RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
     RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
     RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
     RECT 0.81500000 0.44000000 1.10500000 0.51500000 ;
     RECT 3.21500000 0.44000000 3.50500000 0.51500000 ;
     RECT 0.81500000 0.51500000 3.50500000 0.65500000 ;
     RECT 0.81500000 0.65500000 1.10500000 0.73000000 ;
     RECT 3.21500000 0.65500000 3.50500000 0.73000000 ;
     RECT 3.29000000 0.73000000 3.43000000 2.19500000 ;
     RECT 3.21500000 2.19500000 3.50500000 2.48500000 ;
     RECT 0.57500000 2.78000000 0.86500000 3.09000000 ;
     RECT 0.00000000 3.09000000 4.32000000 3.57000000 ;

 END
END NOR2X1
