VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.310 0.720 0.360 ;
        RECT 0.080 0.290 0.090 0.310 ;
        RECT 0.200 0.290 0.210 0.310 ;
        RECT 0.060 0.280 0.090 0.290 ;
        RECT 0.180 0.280 0.210 0.290 ;
        RECT 0.320 0.290 0.330 0.310 ;
        RECT 0.320 0.280 0.350 0.290 ;
        RECT 0.610 0.280 0.640 0.290 ;
        RECT 0.330 0.260 0.620 0.280 ;
        RECT 0.630 0.260 0.640 0.280 ;
        RECT 0.330 0.240 0.340 0.260 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.660 2.150 4.950 2.440 ;
        RECT 0.820 0.610 1.110 0.690 ;
        RECT 4.730 0.610 4.870 2.150 ;
        RECT 6.100 0.610 6.390 0.690 ;
        RECT 0.820 0.470 6.390 0.610 ;
        RECT 0.820 0.400 1.110 0.470 ;
        RECT 6.100 0.400 6.390 0.470 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END A
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.750 4.470 2.040 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 4.180 0.800 4.470 1.090 ;
    END
  END C
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.750 5.910 2.040 ;
        RECT 5.690 1.090 5.830 1.750 ;
        RECT 5.620 0.800 5.910 1.090 ;
    END
  END D
  OBS
      LAYER li1 ;
        RECT 0.080 0.290 0.090 0.310 ;
        RECT 0.200 0.290 0.210 0.310 ;
        RECT 0.060 0.280 0.090 0.290 ;
        RECT 0.180 0.280 0.210 0.290 ;
        RECT 0.320 0.290 0.330 0.310 ;
        RECT 0.320 0.280 0.350 0.290 ;
        RECT 0.610 0.280 0.640 0.290 ;
        RECT 0.610 0.260 0.620 0.280 ;
        RECT 0.630 0.260 0.640 0.280 ;
        RECT 0.610 0.250 0.640 0.260 ;
        RECT 0.080 0.240 0.110 0.250 ;
        RECT 0.180 0.240 0.210 0.250 ;
        RECT 0.080 0.220 0.090 0.240 ;
        RECT 0.200 0.220 0.210 0.240 ;
        RECT 0.080 0.210 0.110 0.220 ;
        RECT 0.180 0.210 0.210 0.220 ;
        RECT 0.220 0.240 0.260 0.250 ;
        RECT 0.220 0.220 0.230 0.240 ;
        RECT 0.250 0.220 0.260 0.240 ;
        RECT 0.220 0.210 0.260 0.220 ;
        RECT 0.320 0.240 0.350 0.250 ;
        RECT 0.460 0.240 0.500 0.250 ;
        RECT 0.320 0.220 0.330 0.240 ;
        RECT 0.460 0.220 0.470 0.240 ;
        RECT 0.490 0.220 0.500 0.240 ;
        RECT 0.320 0.210 0.350 0.220 ;
        RECT 0.470 0.210 0.500 0.220 ;
        RECT 0.130 0.200 0.160 0.210 ;
        RECT 0.130 0.180 0.140 0.200 ;
        RECT 0.150 0.180 0.160 0.200 ;
        RECT 0.130 0.170 0.160 0.180 ;
        RECT 0.270 0.200 0.310 0.210 ;
        RECT 0.420 0.200 0.450 0.210 ;
        RECT 0.270 0.180 0.280 0.200 ;
        RECT 0.300 0.180 0.310 0.200 ;
        RECT 0.440 0.180 0.450 0.200 ;
        RECT 0.270 0.170 0.310 0.180 ;
        RECT 0.420 0.170 0.450 0.180 ;
        RECT 0.560 0.200 0.590 0.210 ;
        RECT 0.560 0.180 0.570 0.200 ;
        RECT 0.560 0.170 0.590 0.180 ;
        RECT 0.130 0.100 0.160 0.110 ;
        RECT 0.130 0.090 0.140 0.100 ;
        RECT 0.150 0.090 0.160 0.100 ;
        RECT 0.130 0.080 0.160 0.090 ;
        RECT 0.270 0.100 0.310 0.110 ;
        RECT 0.420 0.100 0.450 0.110 ;
        RECT 0.270 0.090 0.280 0.100 ;
        RECT 0.300 0.090 0.310 0.100 ;
        RECT 0.440 0.090 0.450 0.100 ;
        RECT 0.270 0.080 0.310 0.090 ;
        RECT 0.420 0.080 0.450 0.090 ;
        RECT 0.560 0.100 0.590 0.110 ;
        RECT 0.560 0.090 0.570 0.100 ;
        RECT 0.560 0.080 0.590 0.090 ;
        RECT 0.080 0.060 0.110 0.070 ;
        RECT 0.460 0.060 0.500 0.070 ;
        RECT 0.080 0.050 0.090 0.060 ;
        RECT 0.460 0.050 0.470 0.060 ;
        RECT 0.490 0.050 0.500 0.060 ;
        RECT 0.080 0.040 0.110 0.050 ;
        RECT 0.460 0.040 0.500 0.050 ;
        RECT 0.610 0.060 0.640 0.070 ;
        RECT 0.610 0.050 0.620 0.060 ;
        RECT 0.630 0.050 0.640 0.060 ;
        RECT 0.610 0.040 0.640 0.050 ;
        RECT 0.200 0.010 0.210 0.040 ;
        RECT 0.320 0.020 0.330 0.040 ;
        RECT 0.320 0.010 0.350 0.020 ;
  END
END AOI22X1
END LIBRARY

