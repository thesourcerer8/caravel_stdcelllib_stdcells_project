VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MUX2X1
  CLASS CORE ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 8.640 3.570 ;
        RECT 1.780 3.060 2.070 3.090 ;
        RECT 1.780 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.070 3.060 ;
        RECT 1.780 2.830 2.070 2.890 ;
        RECT 7.540 3.060 7.830 3.090 ;
        RECT 7.540 2.890 7.600 3.060 ;
        RECT 7.770 2.890 7.830 3.060 ;
        RECT 7.540 2.830 7.830 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.360 2.070 0.420 ;
        RECT 1.780 0.240 1.840 0.360 ;
        RECT 2.010 0.240 2.070 0.360 ;
        RECT 7.540 0.360 7.830 0.420 ;
        RECT 7.540 0.240 7.600 0.360 ;
        RECT 7.770 0.240 7.830 0.360 ;
        RECT 0.000 -0.240 8.640 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.140 2.150 5.430 2.440 ;
        RECT 5.210 1.500 5.350 2.150 ;
        RECT 5.140 1.210 5.430 1.500 ;
    END
  END Y
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.960 5.910 2.040 ;
        RECT 5.620 1.820 6.310 1.960 ;
        RECT 5.620 1.750 5.910 1.820 ;
        RECT 1.300 1.020 1.590 1.090 ;
        RECT 4.180 1.020 4.470 1.090 ;
        RECT 1.300 0.880 4.470 1.020 ;
        RECT 1.300 0.800 1.590 0.880 ;
        RECT 4.180 0.800 4.470 0.880 ;
        RECT 4.250 0.610 4.390 0.800 ;
        RECT 6.170 0.610 6.310 1.820 ;
        RECT 4.250 0.470 6.310 0.610 ;
    END
  END S
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.060 1.750 7.350 2.040 ;
        RECT 7.130 1.090 7.270 1.750 ;
        RECT 7.060 0.800 7.350 1.090 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.210 3.030 1.500 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 3.060 2.090 3.140 ;
        RECT 1.760 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.090 3.060 ;
        RECT 1.760 2.810 2.090 2.890 ;
        RECT 7.520 3.060 7.850 3.140 ;
        RECT 7.520 2.890 7.600 3.060 ;
        RECT 7.770 2.890 7.850 3.060 ;
        RECT 7.520 2.810 7.850 2.890 ;
        RECT 0.560 2.380 0.890 2.460 ;
        RECT 0.560 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.890 2.380 ;
        RECT 0.560 2.130 0.890 2.210 ;
        RECT 5.120 2.380 5.450 2.460 ;
        RECT 5.120 2.210 5.200 2.380 ;
        RECT 5.370 2.210 5.450 2.380 ;
        RECT 5.120 2.130 5.450 2.210 ;
        RECT 1.280 1.980 1.610 2.060 ;
        RECT 1.280 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 2.720 1.980 3.050 2.060 ;
        RECT 2.720 1.810 2.800 1.980 ;
        RECT 2.970 1.810 3.050 1.980 ;
        RECT 2.720 1.730 3.050 1.810 ;
        RECT 4.160 1.980 4.490 2.060 ;
        RECT 4.160 1.810 4.240 1.980 ;
        RECT 4.410 1.810 4.490 1.980 ;
        RECT 5.620 1.980 5.930 2.060 ;
        RECT 5.620 1.960 5.680 1.980 ;
        RECT 4.160 1.730 4.490 1.810 ;
        RECT 5.600 1.810 5.680 1.960 ;
        RECT 5.850 1.810 5.930 1.980 ;
        RECT 5.600 1.730 5.930 1.810 ;
        RECT 7.040 1.980 7.370 2.060 ;
        RECT 7.040 1.810 7.120 1.980 ;
        RECT 7.290 1.810 7.370 1.980 ;
        RECT 7.040 1.730 7.370 1.810 ;
        RECT 1.360 1.110 1.530 1.730 ;
        RECT 2.800 1.440 2.970 1.730 ;
        RECT 2.800 1.110 2.970 1.270 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.860 1.360 1.030 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.280 0.780 1.610 0.860 ;
        RECT 2.720 1.030 3.050 1.110 ;
        RECT 2.720 0.860 2.800 1.030 ;
        RECT 2.970 0.860 3.050 1.030 ;
        RECT 2.720 0.780 3.050 0.860 ;
        RECT 4.160 1.030 4.490 1.110 ;
        RECT 4.160 0.860 4.240 1.030 ;
        RECT 4.410 0.860 4.490 1.030 ;
        RECT 4.160 0.780 4.490 0.860 ;
        RECT 5.200 0.710 5.370 1.270 ;
        RECT 5.600 1.030 5.930 1.110 ;
        RECT 5.600 0.880 5.680 1.030 ;
        RECT 5.620 0.860 5.680 0.880 ;
        RECT 5.850 0.860 5.930 1.030 ;
        RECT 5.620 0.780 5.930 0.860 ;
        RECT 7.040 1.030 7.370 1.110 ;
        RECT 7.040 0.860 7.120 1.030 ;
        RECT 7.290 0.860 7.370 1.030 ;
        RECT 7.040 0.780 7.370 0.860 ;
        RECT 0.560 0.630 0.890 0.710 ;
        RECT 0.560 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.890 0.630 ;
        RECT 0.560 0.380 0.890 0.460 ;
        RECT 5.120 0.630 5.450 0.710 ;
        RECT 5.120 0.460 5.200 0.630 ;
        RECT 5.370 0.460 5.450 0.630 ;
        RECT 1.760 0.360 2.090 0.440 ;
        RECT 5.120 0.380 5.450 0.460 ;
        RECT 1.760 0.190 1.840 0.360 ;
        RECT 2.010 0.190 2.090 0.360 ;
        RECT 1.760 0.110 2.090 0.190 ;
        RECT 7.520 0.360 7.850 0.440 ;
        RECT 7.520 0.190 7.600 0.360 ;
        RECT 7.770 0.190 7.850 0.360 ;
        RECT 7.520 0.110 7.850 0.190 ;
      LAYER met1 ;
        RECT 0.580 2.380 0.870 2.440 ;
        RECT 0.580 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.870 2.380 ;
        RECT 0.580 2.150 0.870 2.210 ;
        RECT 0.650 1.960 0.790 2.150 ;
        RECT 4.180 1.980 4.470 2.040 ;
        RECT 4.180 1.960 4.240 1.980 ;
        RECT 0.650 1.820 4.240 1.960 ;
        RECT 0.650 0.690 0.790 1.820 ;
        RECT 4.180 1.810 4.240 1.820 ;
        RECT 4.410 1.960 4.470 1.980 ;
        RECT 4.410 1.820 4.870 1.960 ;
        RECT 4.410 1.810 4.470 1.820 ;
        RECT 4.180 1.750 4.470 1.810 ;
        RECT 4.730 1.020 4.870 1.820 ;
        RECT 5.620 1.030 5.910 1.090 ;
        RECT 5.620 1.020 5.680 1.030 ;
        RECT 4.730 0.880 5.680 1.020 ;
        RECT 5.620 0.860 5.680 0.880 ;
        RECT 5.850 0.860 5.910 1.030 ;
        RECT 5.620 0.800 5.910 0.860 ;
        RECT 0.580 0.630 0.870 0.690 ;
        RECT 0.580 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.870 0.630 ;
        RECT 0.580 0.400 0.870 0.460 ;
  END
END MUX2X1
END LIBRARY

