magic
tech sky130A
timestamp 1624067079
<< nwell >>
rect 0 179 576 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 226 67 255 73
rect 226 66 232 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 50 232 66
rect 249 66 255 67
rect 466 67 495 73
rect 466 66 472 67
rect 249 50 281 66
rect 152 24 281 50
rect 296 49 425 66
rect 296 32 328 49
rect 345 32 425 49
rect 296 24 425 32
rect 440 50 472 66
rect 489 66 495 67
rect 489 50 519 66
rect 440 24 519 50
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 301 281 309
rect 152 284 184 301
rect 201 284 281 301
rect 152 225 281 284
rect 296 225 425 309
rect 440 243 519 309
rect 440 226 472 243
rect 489 226 519 243
rect 440 225 519 226
rect 58 220 87 225
rect 466 220 495 225
<< ndiffc >>
rect 64 50 81 67
rect 232 50 249 67
rect 328 32 345 49
rect 472 50 489 67
<< pdiffc >>
rect 64 226 81 243
rect 184 284 201 301
rect 472 226 489 243
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
<< locali >>
rect 176 301 209 309
rect 176 284 184 301
rect 201 284 209 301
rect 176 276 209 284
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 464 243 497 251
rect 464 226 472 243
rect 489 226 497 243
rect 464 218 497 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 447 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 92 449 108
rect 441 91 447 92
rect 416 83 447 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 56 42 89 50
rect 224 67 255 75
rect 224 50 232 67
rect 249 66 255 67
rect 464 67 497 75
rect 249 50 257 66
rect 224 42 257 50
rect 320 49 353 57
rect 320 32 328 49
rect 345 32 353 49
rect 464 50 472 67
rect 489 50 497 67
rect 464 42 497 50
rect 320 27 353 32
rect 320 24 328 27
rect 345 24 353 27
<< viali >>
rect 184 284 201 301
rect 64 226 81 243
rect 472 226 489 243
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 64 50 81 67
rect 232 50 249 67
rect 472 50 489 67
rect 328 10 345 27
<< metal1 >>
rect 0 309 576 357
rect 178 301 207 309
rect 178 284 184 301
rect 201 284 207 301
rect 178 278 207 284
rect 58 243 87 249
rect 58 226 64 243
rect 81 241 87 243
rect 466 243 495 249
rect 466 241 472 243
rect 81 227 472 241
rect 81 226 87 227
rect 58 220 87 226
rect 466 226 472 227
rect 489 226 495 243
rect 466 220 495 226
rect 65 73 79 220
rect 130 201 159 207
rect 130 184 136 201
rect 153 184 159 201
rect 130 178 159 184
rect 274 201 303 207
rect 274 184 280 201
rect 297 184 303 201
rect 274 178 303 184
rect 418 201 447 207
rect 418 184 424 201
rect 441 184 447 201
rect 418 178 447 184
rect 137 114 151 178
rect 281 114 295 178
rect 425 114 439 178
rect 130 108 159 114
rect 130 91 136 108
rect 153 91 159 108
rect 130 85 159 91
rect 274 108 303 114
rect 274 91 280 108
rect 297 91 303 108
rect 274 85 303 91
rect 418 108 447 114
rect 418 91 424 108
rect 441 91 447 108
rect 418 85 447 91
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 58 44 87 50
rect 226 67 255 73
rect 226 50 232 67
rect 249 66 255 67
rect 466 67 495 73
rect 466 66 472 67
rect 249 52 472 66
rect 249 50 255 52
rect 226 44 255 50
rect 466 50 472 52
rect 489 50 495 67
rect 466 44 495 50
rect 322 27 351 33
rect 322 24 328 27
rect 0 10 328 24
rect 345 24 351 27
rect 345 10 576 24
rect 0 -24 576 10
<< labels >>
rlabel metal1 0 309 576 357 0 VDD
port 1 se
rlabel metal1 0 -24 576 24 0 GND
port 2 se
rlabel metal1 58 44 87 73 0 Y
port 3 se
rlabel metal1 65 73 79 220 0 Y
port 4 se
rlabel metal1 58 220 87 227 0 Y
port 5 se
rlabel metal1 466 220 495 227 0 Y
port 6 se
rlabel metal1 58 227 495 241 0 Y
port 7 se
rlabel metal1 58 241 87 249 0 Y
port 8 se
rlabel metal1 466 241 495 249 0 Y
port 9 se
rlabel metal1 274 85 303 114 0 A
port 10 se
rlabel metal1 281 114 295 178 0 A
port 11 se
rlabel metal1 274 178 303 207 0 A
port 12 se
rlabel metal1 418 85 447 114 0 B
port 13 se
rlabel metal1 425 114 439 178 0 B
port 14 se
rlabel metal1 418 178 447 207 0 B
port 15 se
rlabel metal1 130 85 159 114 0 C
port 16 se
rlabel metal1 137 114 151 178 0 C
port 17 se
rlabel metal1 130 178 159 207 0 C
port 18 se
<< properties >>
string FIXED_BBOX 0 0 576 333
<< end >>
