VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 15.840 3.570 ;
        RECT 1.780 3.010 2.070 3.090 ;
        RECT 1.780 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.070 3.010 ;
        RECT 1.780 2.780 2.070 2.840 ;
        RECT 4.660 3.010 4.950 3.090 ;
        RECT 4.660 2.840 4.720 3.010 ;
        RECT 4.890 2.840 4.950 3.010 ;
        RECT 4.660 2.780 4.950 2.840 ;
        RECT 7.780 3.010 8.070 3.090 ;
        RECT 7.780 2.840 7.840 3.010 ;
        RECT 8.010 2.840 8.070 3.010 ;
        RECT 7.780 2.780 8.070 2.840 ;
        RECT 11.860 3.010 12.150 3.090 ;
        RECT 11.860 2.840 11.920 3.010 ;
        RECT 12.090 2.840 12.150 3.010 ;
        RECT 11.860 2.780 12.150 2.840 ;
        RECT 13.540 3.010 13.830 3.090 ;
        RECT 13.540 2.840 13.600 3.010 ;
        RECT 13.770 2.840 13.830 3.010 ;
        RECT 13.540 2.780 13.830 2.840 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.490 2.070 0.550 ;
        RECT 1.780 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.070 0.490 ;
        RECT 13.540 0.490 13.830 0.550 ;
        RECT 1.780 0.240 2.070 0.320 ;
        RECT 6.100 0.270 6.390 0.330 ;
        RECT 6.100 0.240 6.160 0.270 ;
        RECT 6.330 0.240 6.390 0.270 ;
        RECT 7.780 0.270 8.070 0.330 ;
        RECT 7.780 0.240 7.840 0.270 ;
        RECT 8.010 0.240 8.070 0.270 ;
        RECT 13.540 0.320 13.600 0.490 ;
        RECT 13.770 0.320 13.830 0.490 ;
        RECT 13.540 0.240 13.830 0.320 ;
        RECT 0.000 -0.240 15.840 0.240 ;
    END
  END gnd
  PIN YC
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.200 0.870 2.490 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 0.580 0.440 0.870 0.730 ;
    END
  END YC
  PIN YS
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 14.740 2.200 15.030 2.490 ;
        RECT 14.810 0.730 14.950 2.200 ;
        RECT 14.740 0.440 15.030 0.730 ;
    END
  END YS
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.780 4.470 2.070 ;
        RECT 4.250 1.140 4.390 1.780 ;
        RECT 4.180 0.850 4.470 1.140 ;
        RECT 9.940 1.060 10.230 1.140 ;
        RECT 6.170 0.920 10.230 1.060 ;
        RECT 4.250 0.660 4.390 0.850 ;
        RECT 6.170 0.660 6.310 0.920 ;
        RECT 9.940 0.850 10.230 0.920 ;
        RECT 4.250 0.520 6.310 0.660 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.780 5.910 2.070 ;
        RECT 11.380 1.780 11.670 2.070 ;
        RECT 5.690 1.470 5.830 1.780 ;
        RECT 11.450 1.470 11.590 1.780 ;
        RECT 5.690 1.330 11.590 1.470 ;
        RECT 5.690 1.140 5.830 1.330 ;
        RECT 11.450 1.140 11.590 1.330 ;
        RECT 5.620 0.850 5.910 1.140 ;
        RECT 11.380 0.850 11.670 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 1.760 3.010 2.090 3.090 ;
        RECT 1.760 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.090 3.010 ;
        RECT 1.760 2.760 2.090 2.840 ;
        RECT 4.640 3.010 4.970 3.090 ;
        RECT 4.640 2.840 4.720 3.010 ;
        RECT 4.890 2.840 4.970 3.010 ;
        RECT 4.640 2.760 4.970 2.840 ;
        RECT 7.760 3.010 8.090 3.090 ;
        RECT 7.760 2.840 7.840 3.010 ;
        RECT 8.010 2.840 8.090 3.010 ;
        RECT 7.760 2.760 8.090 2.840 ;
        RECT 11.840 3.010 12.170 3.090 ;
        RECT 11.840 2.840 11.920 3.010 ;
        RECT 12.090 2.840 12.170 3.010 ;
        RECT 11.840 2.760 12.170 2.840 ;
        RECT 13.520 3.010 13.850 3.090 ;
        RECT 13.520 2.840 13.600 3.010 ;
        RECT 13.770 2.840 13.850 3.010 ;
        RECT 13.520 2.760 13.850 2.840 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 3.440 2.430 3.770 2.510 ;
        RECT 3.440 2.260 3.520 2.430 ;
        RECT 3.690 2.260 3.770 2.430 ;
        RECT 3.440 2.180 3.770 2.260 ;
        RECT 6.080 2.430 6.410 2.510 ;
        RECT 6.080 2.260 6.160 2.430 ;
        RECT 6.330 2.260 6.410 2.430 ;
        RECT 6.080 2.180 6.410 2.260 ;
        RECT 9.440 2.430 9.770 2.510 ;
        RECT 9.440 2.260 9.520 2.430 ;
        RECT 9.690 2.260 9.770 2.430 ;
        RECT 14.720 2.430 15.050 2.510 ;
        RECT 14.720 2.260 14.800 2.430 ;
        RECT 14.970 2.260 15.050 2.430 ;
        RECT 9.440 2.180 9.750 2.260 ;
        RECT 14.740 2.180 15.050 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 2.010 5.910 2.090 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 9.920 2.010 10.250 2.090 ;
        RECT 9.920 1.760 10.000 2.010 ;
        RECT 10.170 1.760 10.250 2.010 ;
        RECT 11.360 2.010 11.690 2.090 ;
        RECT 11.360 1.840 11.440 2.010 ;
        RECT 11.610 1.840 11.690 2.010 ;
        RECT 11.360 1.760 11.690 1.840 ;
        RECT 14.240 2.010 14.570 2.090 ;
        RECT 14.240 1.840 14.320 2.010 ;
        RECT 14.490 1.840 14.570 2.010 ;
        RECT 14.240 1.760 14.570 1.840 ;
        RECT 8.560 1.160 8.730 1.760 ;
        RECT 10.000 1.160 10.170 1.720 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.600 0.830 5.930 0.910 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 8.480 0.910 8.560 1.080 ;
        RECT 8.730 0.910 8.810 1.080 ;
        RECT 8.480 0.830 8.810 0.910 ;
        RECT 9.920 1.080 10.250 1.160 ;
        RECT 9.920 0.910 10.000 1.080 ;
        RECT 10.170 0.920 10.250 1.080 ;
        RECT 10.170 0.910 10.230 0.920 ;
        RECT 9.920 0.830 10.230 0.910 ;
        RECT 10.480 0.750 10.650 1.720 ;
        RECT 11.360 1.080 11.690 1.160 ;
        RECT 11.360 0.910 11.440 1.080 ;
        RECT 11.610 0.910 11.690 1.080 ;
        RECT 11.360 0.830 11.690 0.910 ;
        RECT 14.240 1.080 14.570 1.160 ;
        RECT 14.240 0.910 14.320 1.080 ;
        RECT 14.490 0.920 14.570 1.080 ;
        RECT 14.490 0.910 14.550 0.920 ;
        RECT 14.240 0.830 14.550 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 3.440 0.670 3.770 0.750 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 1.760 0.490 2.090 0.570 ;
        RECT 1.760 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.090 0.490 ;
        RECT 3.440 0.500 3.520 0.670 ;
        RECT 3.690 0.500 3.770 0.670 ;
        RECT 9.440 0.670 9.750 0.750 ;
        RECT 3.440 0.420 3.770 0.500 ;
        RECT 6.080 0.490 6.410 0.570 ;
        RECT 1.760 0.240 2.090 0.320 ;
        RECT 6.080 0.320 6.160 0.490 ;
        RECT 6.330 0.320 6.410 0.490 ;
        RECT 6.080 0.270 6.410 0.320 ;
        RECT 6.080 0.240 6.160 0.270 ;
        RECT 6.330 0.240 6.410 0.270 ;
        RECT 7.760 0.490 8.090 0.570 ;
        RECT 7.760 0.320 7.840 0.490 ;
        RECT 8.010 0.320 8.090 0.490 ;
        RECT 9.440 0.500 9.520 0.670 ;
        RECT 9.690 0.660 9.750 0.670 ;
        RECT 10.400 0.670 10.730 0.750 ;
        RECT 9.690 0.500 9.770 0.660 ;
        RECT 9.440 0.420 9.770 0.500 ;
        RECT 10.400 0.500 10.480 0.670 ;
        RECT 10.650 0.500 10.730 0.670 ;
        RECT 11.860 0.670 12.170 0.750 ;
        RECT 11.860 0.660 11.920 0.670 ;
        RECT 10.400 0.420 10.730 0.500 ;
        RECT 11.840 0.500 11.920 0.660 ;
        RECT 12.090 0.500 12.170 0.670 ;
        RECT 14.720 0.670 15.050 0.750 ;
        RECT 11.840 0.420 12.170 0.500 ;
        RECT 13.520 0.490 13.850 0.570 ;
        RECT 7.760 0.270 8.090 0.320 ;
        RECT 7.760 0.240 7.840 0.270 ;
        RECT 8.010 0.240 8.090 0.270 ;
        RECT 13.520 0.320 13.600 0.490 ;
        RECT 13.770 0.320 13.850 0.490 ;
        RECT 14.720 0.500 14.800 0.670 ;
        RECT 14.970 0.500 15.050 0.670 ;
        RECT 14.720 0.420 15.050 0.500 ;
        RECT 13.520 0.240 13.850 0.320 ;
      LAYER met1 ;
        RECT 3.460 2.430 3.750 2.490 ;
        RECT 3.460 2.260 3.520 2.430 ;
        RECT 3.690 2.410 3.750 2.430 ;
        RECT 6.100 2.430 6.390 2.490 ;
        RECT 6.100 2.410 6.160 2.430 ;
        RECT 3.690 2.270 6.160 2.410 ;
        RECT 3.690 2.260 3.750 2.270 ;
        RECT 3.460 2.200 3.750 2.260 ;
        RECT 6.100 2.260 6.160 2.270 ;
        RECT 6.330 2.410 6.390 2.430 ;
        RECT 9.460 2.430 9.750 2.490 ;
        RECT 6.330 2.270 8.710 2.410 ;
        RECT 6.330 2.260 6.390 2.270 ;
        RECT 6.100 2.200 6.390 2.260 ;
        RECT 1.300 2.010 1.590 2.070 ;
        RECT 1.300 1.840 1.360 2.010 ;
        RECT 1.530 2.000 1.590 2.010 ;
        RECT 3.530 2.000 3.670 2.200 ;
        RECT 8.570 2.070 8.710 2.270 ;
        RECT 9.460 2.260 9.520 2.430 ;
        RECT 9.690 2.410 9.750 2.430 ;
        RECT 9.690 2.270 14.470 2.410 ;
        RECT 9.690 2.260 9.750 2.270 ;
        RECT 9.460 2.200 9.750 2.260 ;
        RECT 1.530 1.860 3.670 2.000 ;
        RECT 1.530 1.840 1.590 1.860 ;
        RECT 1.300 1.780 1.590 1.840 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 1.080 1.590 1.140 ;
        RECT 1.300 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.590 1.080 ;
        RECT 1.300 0.850 1.590 0.910 ;
        RECT 3.530 0.730 3.670 1.860 ;
        RECT 8.500 2.010 8.790 2.070 ;
        RECT 8.500 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.790 2.010 ;
        RECT 8.500 1.780 8.790 1.840 ;
        RECT 9.940 2.010 10.230 2.070 ;
        RECT 9.940 1.720 10.000 2.010 ;
        RECT 10.170 1.720 10.230 2.010 ;
        RECT 10.490 1.950 10.630 2.270 ;
        RECT 14.330 2.070 14.470 2.270 ;
        RECT 14.260 2.010 14.550 2.070 ;
        RECT 9.940 1.660 10.230 1.720 ;
        RECT 10.420 1.890 10.710 1.950 ;
        RECT 10.420 1.720 10.480 1.890 ;
        RECT 10.650 1.720 10.710 1.890 ;
        RECT 14.260 1.840 14.320 2.010 ;
        RECT 14.490 1.840 14.550 2.010 ;
        RECT 14.260 1.780 14.550 1.840 ;
        RECT 10.420 1.660 10.710 1.720 ;
        RECT 14.330 1.140 14.470 1.780 ;
        RECT 14.260 1.080 14.550 1.140 ;
        RECT 14.260 0.910 14.320 1.080 ;
        RECT 14.490 0.910 14.550 1.080 ;
        RECT 14.260 0.850 14.550 0.910 ;
        RECT 3.460 0.670 3.750 0.730 ;
        RECT 3.460 0.500 3.520 0.670 ;
        RECT 3.690 0.500 3.750 0.670 ;
        RECT 3.460 0.440 3.750 0.500 ;
        RECT 9.460 0.670 9.750 0.730 ;
        RECT 9.460 0.500 9.520 0.670 ;
        RECT 9.690 0.660 9.750 0.670 ;
        RECT 11.860 0.670 12.150 0.730 ;
        RECT 11.860 0.660 11.920 0.670 ;
        RECT 9.690 0.520 11.920 0.660 ;
        RECT 9.690 0.500 9.750 0.520 ;
        RECT 9.460 0.440 9.750 0.500 ;
        RECT 11.860 0.500 11.920 0.520 ;
        RECT 12.090 0.500 12.150 0.670 ;
        RECT 11.860 0.440 12.150 0.500 ;
  END
END HAX1
END LIBRARY

