VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO VANBERKEL1991
  CLASS CORE ;
  FOREIGN VANBERKEL1991 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 8.980 2.970 9.270 3.090 ;
        RECT 8.980 2.800 9.040 2.970 ;
        RECT 9.210 2.800 9.270 2.970 ;
        RECT 8.980 2.740 9.270 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 11.520 3.570 ;
        RECT 4.640 2.970 4.970 3.090 ;
        RECT 4.640 2.800 4.720 2.970 ;
        RECT 4.890 2.800 4.970 2.970 ;
        RECT 4.640 2.720 4.970 2.800 ;
        RECT 8.960 2.970 9.290 3.090 ;
        RECT 8.960 2.800 9.040 2.970 ;
        RECT 9.210 2.800 9.290 2.970 ;
        RECT 8.960 2.720 9.290 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.640 0.670 4.970 0.750 ;
        RECT 4.640 0.500 4.720 0.670 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
        RECT 8.960 0.670 9.290 0.750 ;
        RECT 8.960 0.500 9.040 0.670 ;
        RECT 9.210 0.500 9.290 0.670 ;
        RECT 8.960 0.420 9.290 0.500 ;
        RECT 4.720 0.240 4.890 0.420 ;
        RECT 9.040 0.240 9.210 0.420 ;
        RECT 0.000 -0.240 11.520 0.240 ;
    END
  END VGND
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.060 2.410 7.350 2.490 ;
        RECT 10.420 2.410 10.710 2.490 ;
        RECT 7.060 2.270 10.710 2.410 ;
        RECT 7.060 2.200 7.350 2.270 ;
        RECT 10.420 2.200 10.710 2.270 ;
        RECT 10.490 0.730 10.630 2.200 ;
        RECT 10.420 0.440 10.710 0.730 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.060 3.030 1.140 ;
        RECT 8.500 1.060 8.790 1.140 ;
        RECT 2.740 0.920 8.790 1.060 ;
        RECT 2.740 0.850 3.030 0.920 ;
        RECT 8.500 0.850 8.790 0.920 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
        RECT 1.370 0.660 1.510 0.850 ;
        RECT 3.220 0.660 3.510 0.730 ;
        RECT 1.370 0.520 3.510 0.660 ;
        RECT 3.220 0.440 3.510 0.520 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.800 2.830 1.130 2.910 ;
        RECT 0.800 2.660 0.880 2.830 ;
        RECT 1.050 2.660 1.130 2.830 ;
        RECT 0.800 2.580 1.130 2.660 ;
        RECT 7.520 2.830 7.850 2.910 ;
        RECT 7.520 2.660 7.600 2.830 ;
        RECT 7.770 2.660 7.850 2.830 ;
        RECT 7.520 2.580 7.850 2.660 ;
        RECT 1.760 2.430 2.090 2.510 ;
        RECT 1.760 2.260 1.840 2.430 ;
        RECT 2.010 2.260 2.090 2.430 ;
        RECT 1.780 2.180 2.090 2.260 ;
        RECT 3.680 2.430 4.010 2.510 ;
        RECT 3.680 2.260 3.760 2.430 ;
        RECT 3.930 2.260 4.010 2.430 ;
        RECT 6.320 2.430 6.650 2.510 ;
        RECT 6.320 2.260 6.400 2.430 ;
        RECT 6.570 2.260 6.650 2.430 ;
        RECT 10.400 2.430 10.730 2.510 ;
        RECT 10.400 2.260 10.480 2.430 ;
        RECT 10.650 2.260 10.730 2.430 ;
        RECT 3.680 2.180 3.990 2.260 ;
        RECT 6.320 2.180 6.650 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.840 1.890 2.010 2.180 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.920 1.610 1.080 ;
        RECT 1.530 0.910 1.590 0.920 ;
        RECT 1.280 0.830 1.590 0.910 ;
        RECT 1.840 0.750 2.010 1.720 ;
        RECT 2.320 1.480 2.490 2.120 ;
        RECT 7.120 2.090 7.290 2.260 ;
        RECT 10.420 2.180 10.730 2.260 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 8.480 2.010 8.810 2.090 ;
        RECT 8.480 1.840 8.560 2.010 ;
        RECT 8.730 1.840 8.810 2.010 ;
        RECT 8.480 1.760 8.810 1.840 ;
        RECT 9.920 2.010 10.250 2.090 ;
        RECT 9.920 1.840 10.000 2.010 ;
        RECT 10.170 1.840 10.250 2.010 ;
        RECT 9.920 1.760 10.250 1.840 ;
        RECT 2.800 1.160 2.970 1.760 ;
        RECT 4.240 1.210 4.410 1.760 ;
        RECT 3.280 1.160 4.410 1.210 ;
        RECT 7.120 1.160 7.290 1.760 ;
        RECT 8.560 1.160 8.730 1.760 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 3.280 1.080 4.490 1.160 ;
        RECT 3.280 1.040 4.240 1.080 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 1.760 0.670 2.090 0.750 ;
        RECT 3.280 0.670 3.450 1.040 ;
        RECT 4.160 0.910 4.240 1.040 ;
        RECT 4.410 0.920 4.490 1.080 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 4.410 0.910 4.470 0.920 ;
        RECT 4.160 0.830 4.470 0.910 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.370 1.080 ;
        RECT 8.480 1.080 8.810 1.160 ;
        RECT 8.480 0.920 8.560 1.080 ;
        RECT 7.040 0.830 7.370 0.910 ;
        RECT 8.500 0.910 8.560 0.920 ;
        RECT 8.730 0.920 8.810 1.080 ;
        RECT 9.920 1.080 10.250 1.160 ;
        RECT 8.730 0.910 8.790 0.920 ;
        RECT 8.500 0.830 8.790 0.910 ;
        RECT 9.920 0.910 10.000 1.080 ;
        RECT 10.170 0.920 10.250 1.080 ;
        RECT 10.170 0.910 10.230 0.920 ;
        RECT 9.920 0.830 10.230 0.910 ;
        RECT 3.680 0.670 3.990 0.750 ;
        RECT 1.760 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.090 0.670 ;
        RECT 1.760 0.420 2.090 0.500 ;
        RECT 3.680 0.500 3.760 0.670 ;
        RECT 3.930 0.660 3.990 0.670 ;
        RECT 6.320 0.670 6.650 0.750 ;
        RECT 3.930 0.500 4.010 0.660 ;
        RECT 3.680 0.420 4.010 0.500 ;
        RECT 6.320 0.500 6.400 0.670 ;
        RECT 6.570 0.500 6.650 0.670 ;
        RECT 6.320 0.420 6.650 0.500 ;
        RECT 8.000 0.670 8.330 0.750 ;
        RECT 8.000 0.500 8.080 0.670 ;
        RECT 8.250 0.500 8.330 0.670 ;
        RECT 8.000 0.420 8.330 0.500 ;
        RECT 10.400 0.670 10.730 0.750 ;
        RECT 10.400 0.500 10.480 0.670 ;
        RECT 10.650 0.500 10.730 0.670 ;
        RECT 10.400 0.420 10.730 0.500 ;
      LAYER met1 ;
        RECT 0.820 2.830 1.110 2.890 ;
        RECT 0.820 2.660 0.880 2.830 ;
        RECT 1.050 2.820 1.110 2.830 ;
        RECT 7.540 2.830 7.830 2.890 ;
        RECT 7.540 2.820 7.600 2.830 ;
        RECT 1.050 2.680 7.600 2.820 ;
        RECT 1.050 2.660 1.110 2.680 ;
        RECT 0.820 2.600 1.110 2.660 ;
        RECT 7.540 2.660 7.600 2.680 ;
        RECT 7.770 2.660 7.830 2.830 ;
        RECT 7.540 2.600 7.830 2.660 ;
        RECT 3.700 2.430 3.990 2.490 ;
        RECT 0.650 2.350 2.470 2.410 ;
        RECT 0.650 2.290 2.550 2.350 ;
        RECT 0.650 2.270 2.320 2.290 ;
        RECT 0.650 0.730 0.790 2.270 ;
        RECT 2.260 2.120 2.320 2.270 ;
        RECT 2.490 2.120 2.550 2.290 ;
        RECT 3.700 2.260 3.760 2.430 ;
        RECT 3.930 2.410 3.990 2.430 ;
        RECT 6.340 2.430 6.630 2.490 ;
        RECT 6.340 2.410 6.400 2.430 ;
        RECT 3.930 2.270 6.400 2.410 ;
        RECT 3.930 2.260 3.990 2.270 ;
        RECT 3.700 2.200 3.990 2.260 ;
        RECT 6.340 2.260 6.400 2.270 ;
        RECT 6.570 2.260 6.630 2.430 ;
        RECT 6.340 2.200 6.630 2.260 ;
        RECT 2.260 2.060 2.550 2.120 ;
        RECT 9.940 2.010 10.230 2.070 ;
        RECT 1.780 1.890 2.070 1.950 ;
        RECT 1.780 1.720 1.840 1.890 ;
        RECT 2.010 1.870 2.070 1.890 ;
        RECT 9.940 1.870 10.000 2.010 ;
        RECT 2.010 1.840 10.000 1.870 ;
        RECT 10.170 1.840 10.230 2.010 ;
        RECT 2.010 1.780 10.230 1.840 ;
        RECT 2.010 1.730 10.150 1.780 ;
        RECT 2.010 1.720 2.070 1.730 ;
        RECT 1.780 1.660 2.070 1.720 ;
        RECT 2.260 1.480 2.550 1.540 ;
        RECT 2.260 1.310 2.320 1.480 ;
        RECT 2.490 1.470 2.550 1.480 ;
        RECT 2.490 1.330 9.190 1.470 ;
        RECT 2.490 1.310 2.550 1.330 ;
        RECT 2.260 1.250 2.550 1.310 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 3.700 0.670 3.990 0.730 ;
        RECT 3.700 0.500 3.760 0.670 ;
        RECT 3.930 0.660 3.990 0.670 ;
        RECT 6.340 0.670 6.630 0.730 ;
        RECT 6.340 0.660 6.400 0.670 ;
        RECT 3.930 0.520 6.400 0.660 ;
        RECT 3.930 0.500 3.990 0.520 ;
        RECT 3.700 0.440 3.990 0.500 ;
        RECT 6.340 0.500 6.400 0.520 ;
        RECT 6.570 0.500 6.630 0.670 ;
        RECT 6.340 0.440 6.630 0.500 ;
        RECT 8.020 0.670 8.310 0.730 ;
        RECT 8.020 0.500 8.080 0.670 ;
        RECT 8.250 0.660 8.310 0.670 ;
        RECT 9.050 0.660 9.190 1.330 ;
        RECT 10.010 1.140 10.150 1.730 ;
        RECT 9.940 1.080 10.230 1.140 ;
        RECT 9.940 0.910 10.000 1.080 ;
        RECT 10.170 0.910 10.230 1.080 ;
        RECT 9.940 0.850 10.230 0.910 ;
        RECT 8.250 0.520 9.190 0.660 ;
        RECT 8.250 0.500 8.310 0.520 ;
        RECT 8.020 0.440 8.310 0.500 ;
  END
END VANBERKEL1991
END LIBRARY

