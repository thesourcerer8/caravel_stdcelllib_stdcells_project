VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MARTIN1989
  CLASS CORE ;
  FOREIGN MARTIN1989 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 7.200 3.570 ;
        RECT 0.580 2.970 0.870 3.090 ;
        RECT 0.580 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.870 2.970 ;
        RECT 0.580 2.740 0.870 2.800 ;
        RECT 4.660 2.970 4.950 3.090 ;
        RECT 4.660 2.800 4.720 2.970 ;
        RECT 4.890 2.800 4.950 2.970 ;
        RECT 4.660 2.740 4.950 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 7.200 3.570 ;
        RECT 0.560 2.970 0.890 3.090 ;
        RECT 0.560 2.800 0.640 2.970 ;
        RECT 0.810 2.800 0.890 2.970 ;
        RECT 0.560 2.720 0.890 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
        RECT 0.650 0.240 0.790 0.440 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.660 0.670 4.970 0.750 ;
        RECT 4.660 0.660 4.720 0.670 ;
        RECT 4.640 0.500 4.720 0.660 ;
        RECT 4.890 0.500 4.970 0.670 ;
        RECT 4.640 0.420 4.970 0.500 ;
        RECT 4.720 0.240 4.890 0.420 ;
        RECT 0.000 -0.240 7.200 0.240 ;
    END
  END VGND
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 6.100 2.200 6.390 2.490 ;
        RECT 4.180 0.850 4.470 1.140 ;
        RECT 4.250 0.660 4.390 0.850 ;
        RECT 6.170 0.730 6.310 2.200 ;
        RECT 6.100 0.660 6.390 0.730 ;
        RECT 4.250 0.520 6.390 0.660 ;
        RECT 6.100 0.440 6.390 0.520 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.780 3.030 2.070 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 2.740 0.850 3.030 1.140 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 4.640 2.970 4.970 3.050 ;
        RECT 4.640 2.800 4.720 2.970 ;
        RECT 4.890 2.800 4.970 2.970 ;
        RECT 4.640 2.720 4.970 2.800 ;
        RECT 3.200 2.430 3.530 2.510 ;
        RECT 3.200 2.260 3.280 2.430 ;
        RECT 3.450 2.260 3.530 2.430 ;
        RECT 6.080 2.430 6.410 2.510 ;
        RECT 6.080 2.260 6.160 2.430 ;
        RECT 6.330 2.260 6.410 2.430 ;
        RECT 3.220 2.180 3.530 2.260 ;
        RECT 6.100 2.180 6.410 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 2.010 5.930 2.090 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 4.240 1.160 4.410 1.760 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.920 3.050 1.080 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 2.970 0.910 3.030 0.920 ;
        RECT 2.720 0.830 3.030 0.910 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.910 5.680 1.080 ;
        RECT 5.850 0.920 5.930 1.080 ;
        RECT 5.850 0.910 5.910 0.920 ;
        RECT 5.600 0.830 5.910 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 3.200 0.670 3.530 0.750 ;
        RECT 3.200 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
        RECT 6.080 0.670 6.410 0.750 ;
        RECT 6.080 0.500 6.160 0.670 ;
        RECT 6.330 0.500 6.410 0.670 ;
        RECT 6.080 0.420 6.410 0.500 ;
      LAYER met1 ;
        RECT 3.220 2.430 3.510 2.490 ;
        RECT 3.220 2.260 3.280 2.430 ;
        RECT 3.450 2.260 3.510 2.430 ;
        RECT 3.220 2.200 3.510 2.260 ;
        RECT 3.290 2.000 3.430 2.200 ;
        RECT 5.620 2.010 5.910 2.070 ;
        RECT 5.620 2.000 5.680 2.010 ;
        RECT 3.290 1.860 5.680 2.000 ;
        RECT 3.290 0.730 3.430 1.860 ;
        RECT 5.620 1.840 5.680 1.860 ;
        RECT 5.850 1.840 5.910 2.010 ;
        RECT 5.620 1.780 5.910 1.840 ;
        RECT 5.690 1.140 5.830 1.780 ;
        RECT 5.620 1.080 5.910 1.140 ;
        RECT 5.620 0.910 5.680 1.080 ;
        RECT 5.850 0.910 5.910 1.080 ;
        RECT 5.620 0.850 5.910 0.910 ;
        RECT 3.220 0.670 3.510 0.730 ;
        RECT 3.220 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.510 0.670 ;
        RECT 3.220 0.440 3.510 0.500 ;
  END
END MARTIN1989
END LIBRARY

