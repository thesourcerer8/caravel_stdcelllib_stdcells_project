VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.960 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.370 2.675 2.950 2.815 ;
        RECT 1.370 2.070 1.510 2.675 ;
        RECT 2.810 2.070 2.950 2.675 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 2.810 1.540 2.950 1.780 ;
        RECT 2.735 1.250 3.025 1.540 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.795 1.155 2.965 1.480 ;
        RECT 2.715 0.825 3.045 1.155 ;
      LAYER mcon ;
        RECT 2.795 1.310 2.965 1.480 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.275 1.760 1.605 2.090 ;
      LAYER mcon ;
        RECT 1.355 1.840 1.525 2.010 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.715 1.760 3.045 2.090 ;
      LAYER mcon ;
        RECT 2.795 1.840 2.965 2.010 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 2.289000 ;
    PORT
      LAYER met1 ;
        RECT 0.575 0.240 0.865 0.570 ;
        RECT 3.215 0.240 3.505 0.570 ;
        RECT 6.095 0.240 6.385 0.570 ;
        RECT 8.975 0.240 9.265 0.570 ;
        RECT 11.855 0.240 12.145 0.570 ;
        RECT 0.000 -0.240 12.960 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.555 0.240 0.885 0.590 ;
        RECT 3.195 0.240 3.525 0.590 ;
        RECT 6.075 0.240 6.405 0.590 ;
        RECT 8.955 0.240 9.285 0.590 ;
        RECT 11.835 0.240 12.165 0.590 ;
        RECT 0.155 0.085 12.805 0.240 ;
        RECT 0.000 -0.085 12.960 0.085 ;
      LAYER mcon ;
        RECT 0.635 0.340 0.805 0.510 ;
        RECT 3.275 0.340 3.445 0.510 ;
        RECT 6.155 0.340 6.325 0.510 ;
        RECT 9.035 0.340 9.205 0.510 ;
        RECT 11.915 0.340 12.085 0.510 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 12.960 3.570 ;
        RECT 0.575 2.760 0.865 3.090 ;
        RECT 3.215 2.760 3.505 3.090 ;
        RECT 6.095 2.760 6.385 3.090 ;
        RECT 8.975 2.760 9.265 3.090 ;
        RECT 11.855 2.760 12.145 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 4.578000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 12.960 3.415 ;
        RECT 0.155 3.090 12.805 3.245 ;
        RECT 0.555 2.740 0.885 3.090 ;
        RECT 3.195 2.740 3.525 3.090 ;
        RECT 6.075 2.740 6.405 3.090 ;
        RECT 8.955 2.740 9.285 3.090 ;
        RECT 11.835 2.740 12.165 3.090 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 0.635 2.820 0.805 2.990 ;
        RECT 3.275 2.820 3.445 2.990 ;
        RECT 6.155 2.820 6.325 2.990 ;
        RECT 9.035 2.820 9.205 2.990 ;
        RECT 11.915 2.820 12.085 2.990 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 10.415 0.440 10.705 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 12.960 3.330 ;
      LAYER li1 ;
        RECT 1.755 2.260 2.085 2.505 ;
        RECT 4.635 2.260 4.965 2.505 ;
        RECT 1.775 2.175 2.085 2.260 ;
        RECT 4.655 2.175 4.965 2.260 ;
        RECT 5.675 2.090 5.845 2.830 ;
        RECT 7.515 2.175 7.845 2.505 ;
        RECT 8.555 2.090 8.725 2.830 ;
        RECT 10.395 2.260 10.725 2.505 ;
        RECT 10.415 2.175 10.725 2.260 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 7.035 2.005 7.345 2.090 ;
        RECT 7.035 1.760 7.365 2.005 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 5.675 1.445 5.845 1.760 ;
        RECT 8.555 1.445 8.725 1.760 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 4.155 0.920 4.485 1.155 ;
        RECT 4.155 0.825 4.465 0.920 ;
        RECT 5.595 0.825 5.925 1.155 ;
        RECT 7.035 0.920 7.365 1.155 ;
        RECT 7.035 0.825 7.345 0.920 ;
        RECT 8.475 0.825 8.805 1.155 ;
        RECT 9.915 0.920 10.245 1.155 ;
        RECT 9.915 0.825 10.225 0.920 ;
        RECT 10.475 0.750 10.645 2.175 ;
        RECT 11.355 1.760 11.685 2.090 ;
        RECT 11.355 0.825 11.685 1.155 ;
        RECT 1.775 0.655 2.085 0.750 ;
        RECT 1.755 0.420 2.085 0.655 ;
        RECT 4.635 0.420 4.965 0.750 ;
        RECT 7.515 0.420 7.845 0.750 ;
        RECT 10.395 0.420 10.725 0.750 ;
      LAYER mcon ;
        RECT 5.675 2.660 5.845 2.830 ;
        RECT 1.835 2.255 2.005 2.425 ;
        RECT 4.715 2.255 4.885 2.425 ;
        RECT 8.555 2.660 8.725 2.830 ;
        RECT 7.595 2.255 7.765 2.425 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 7.115 1.840 7.285 2.010 ;
        RECT 9.995 1.840 10.165 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 7.115 0.905 7.285 1.075 ;
        RECT 8.555 0.905 8.725 1.075 ;
        RECT 9.995 0.905 10.165 1.075 ;
        RECT 11.435 1.840 11.605 2.010 ;
        RECT 11.435 0.905 11.605 1.075 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 4.715 0.500 4.885 0.670 ;
        RECT 7.595 0.500 7.765 0.670 ;
        RECT 10.475 0.500 10.645 0.670 ;
      LAYER met1 ;
        RECT 5.615 2.815 5.905 2.890 ;
        RECT 8.495 2.815 8.785 2.890 ;
        RECT 4.250 2.675 5.905 2.815 ;
        RECT 1.775 2.195 2.065 2.485 ;
        RECT 1.850 1.060 1.990 2.195 ;
        RECT 4.250 2.070 4.390 2.675 ;
        RECT 5.615 2.600 5.905 2.675 ;
        RECT 7.130 2.675 8.785 2.815 ;
        RECT 4.655 2.195 4.945 2.485 ;
        RECT 4.175 1.780 4.465 2.070 ;
        RECT 4.730 1.995 4.870 2.195 ;
        RECT 7.130 2.070 7.270 2.675 ;
        RECT 8.495 2.600 8.785 2.675 ;
        RECT 7.535 2.195 7.825 2.485 ;
        RECT 7.055 1.995 7.345 2.070 ;
        RECT 4.730 1.855 7.345 1.995 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 1.850 0.920 4.465 1.060 ;
        RECT 1.850 0.730 1.990 0.920 ;
        RECT 4.175 0.845 4.465 0.920 ;
        RECT 4.730 0.730 4.870 1.855 ;
        RECT 7.055 1.780 7.345 1.855 ;
        RECT 7.610 1.995 7.750 2.195 ;
        RECT 9.935 1.995 10.225 2.070 ;
        RECT 11.375 1.995 11.665 2.070 ;
        RECT 7.610 1.855 11.665 1.995 ;
        RECT 5.615 1.385 5.905 1.675 ;
        RECT 5.690 1.135 5.830 1.385 ;
        RECT 7.130 1.135 7.270 1.780 ;
        RECT 5.615 0.845 5.905 1.135 ;
        RECT 7.055 0.845 7.345 1.135 ;
        RECT 7.610 0.730 7.750 1.855 ;
        RECT 9.935 1.780 10.225 1.855 ;
        RECT 11.375 1.780 11.665 1.855 ;
        RECT 8.495 1.385 8.785 1.675 ;
        RECT 8.570 1.135 8.710 1.385 ;
        RECT 10.010 1.135 10.150 1.780 ;
        RECT 11.450 1.135 11.590 1.780 ;
        RECT 8.495 0.845 8.785 1.135 ;
        RECT 9.935 0.845 10.225 1.135 ;
        RECT 11.375 0.845 11.665 1.135 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 4.655 0.440 4.945 0.730 ;
        RECT 7.535 0.440 7.825 0.730 ;
  END
END CLKBUF1
END LIBRARY

