MACRO AOI21X1
 CLASS CORE ;
 FOREIGN AOI21X1 0 0 ;
 SIZE 5.76 BY 3.33 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;
       LAYER met1 ;
        RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER li1 ;
        RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.57500000 0.44000000 0.86500000 0.51500000 ;
        RECT 4.65500000 0.44000000 4.94500000 0.51500000 ;
        RECT 0.57500000 0.51500000 4.94500000 0.65500000 ;
        RECT 0.57500000 0.65500000 0.86500000 0.73000000 ;
        RECT 4.65500000 0.65500000 4.94500000 0.73000000 ;
        RECT 0.65000000 0.73000000 0.79000000 2.19500000 ;
        RECT 0.57500000 2.19500000 0.86500000 2.48500000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
        RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
        RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
    END
  END C

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
        RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
        RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 4.17500000 0.84500000 4.46500000 1.13500000 ;
        RECT 4.25000000 1.13500000 4.39000000 1.78000000 ;
        RECT 4.17500000 1.78000000 4.46500000 2.07000000 ;
    END
  END B

 OBS
    LAYER polycont ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;

    LAYER pdiffc ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 2.31500000 2.25500000 2.48500000 2.42500000 ;
     RECT 4.71500000 2.25500000 4.88500000 2.42500000 ;
     RECT 3.27500000 2.82000000 3.44500000 2.99000000 ;

    LAYER ndiffc ;
     RECT 1.83500000 0.34000000 2.00500000 0.51000000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 4.71500000 0.50000000 4.88500000 0.67000000 ;

    LAYER li1 ;
     RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
     RECT 1.75500000 0.24000000 2.08500000 0.59000000 ;
     RECT 0.55500000 0.42000000 0.88500000 0.75000000 ;
     RECT 4.63500000 0.42000000 4.96500000 0.75000000 ;
     RECT 1.27500000 0.82500000 1.60500000 1.15500000 ;
     RECT 2.71500000 0.82500000 3.04500000 1.15500000 ;
     RECT 4.15500000 0.82500000 4.48500000 1.15500000 ;
     RECT 1.27500000 1.76000000 1.60500000 2.09000000 ;
     RECT 2.71500000 1.76000000 3.04500000 2.09000000 ;
     RECT 4.15500000 1.76000000 4.48500000 2.09000000 ;
     RECT 0.55500000 2.17500000 0.88500000 2.50500000 ;
     RECT 2.23500000 2.17500000 2.56500000 2.50500000 ;
     RECT 4.63500000 2.17500000 4.96500000 2.50500000 ;
     RECT 3.19500000 2.74000000 3.52500000 3.07000000 ;
     RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;

    LAYER viali ;
     RECT 0.15500000 -0.08500000 0.32500000 0.08500000 ;
     RECT 0.63500000 -0.08500000 0.80500000 0.08500000 ;
     RECT 1.11500000 -0.08500000 1.28500000 0.08500000 ;
     RECT 1.59500000 -0.08500000 1.76500000 0.08500000 ;
     RECT 2.07500000 -0.08500000 2.24500000 0.08500000 ;
     RECT 2.55500000 -0.08500000 2.72500000 0.08500000 ;
     RECT 3.03500000 -0.08500000 3.20500000 0.08500000 ;
     RECT 3.51500000 -0.08500000 3.68500000 0.08500000 ;
     RECT 3.99500000 -0.08500000 4.16500000 0.08500000 ;
     RECT 4.47500000 -0.08500000 4.64500000 0.08500000 ;
     RECT 4.95500000 -0.08500000 5.12500000 0.08500000 ;
     RECT 5.43500000 -0.08500000 5.60500000 0.08500000 ;
     RECT 0.63500000 0.50000000 0.80500000 0.67000000 ;
     RECT 4.71500000 0.50000000 4.88500000 0.67000000 ;
     RECT 1.35500000 0.90500000 1.52500000 1.07500000 ;
     RECT 2.79500000 0.90500000 2.96500000 1.07500000 ;
     RECT 4.23500000 0.90500000 4.40500000 1.07500000 ;
     RECT 1.35500000 1.84000000 1.52500000 2.01000000 ;
     RECT 2.79500000 1.84000000 2.96500000 2.01000000 ;
     RECT 4.23500000 1.84000000 4.40500000 2.01000000 ;
     RECT 0.63500000 2.25500000 0.80500000 2.42500000 ;
     RECT 2.31500000 2.25500000 2.48500000 2.42500000 ;
     RECT 4.71500000 2.25500000 4.88500000 2.42500000 ;
     RECT 3.27500000 2.82000000 3.44500000 2.99000000 ;
     RECT 0.15500000 3.24500000 0.32500000 3.41500000 ;
     RECT 0.63500000 3.24500000 0.80500000 3.41500000 ;
     RECT 1.11500000 3.24500000 1.28500000 3.41500000 ;
     RECT 1.59500000 3.24500000 1.76500000 3.41500000 ;
     RECT 2.07500000 3.24500000 2.24500000 3.41500000 ;
     RECT 2.55500000 3.24500000 2.72500000 3.41500000 ;
     RECT 3.03500000 3.24500000 3.20500000 3.41500000 ;
     RECT 3.51500000 3.24500000 3.68500000 3.41500000 ;
     RECT 3.99500000 3.24500000 4.16500000 3.41500000 ;
     RECT 4.47500000 3.24500000 4.64500000 3.41500000 ;
     RECT 4.95500000 3.24500000 5.12500000 3.41500000 ;
     RECT 5.43500000 3.24500000 5.60500000 3.41500000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 5.76000000 0.24000000 ;
     RECT 1.29500000 0.84500000 1.58500000 1.13500000 ;
     RECT 1.37000000 1.13500000 1.51000000 1.78000000 ;
     RECT 1.29500000 1.78000000 1.58500000 2.07000000 ;
     RECT 2.73500000 0.84500000 3.02500000 1.13500000 ;
     RECT 2.81000000 1.13500000 2.95000000 1.78000000 ;
     RECT 2.73500000 1.78000000 3.02500000 2.07000000 ;
     RECT 4.17500000 0.84500000 4.46500000 1.13500000 ;
     RECT 4.25000000 1.13500000 4.39000000 1.78000000 ;
     RECT 4.17500000 1.78000000 4.46500000 2.07000000 ;
     RECT 0.57500000 0.44000000 0.86500000 0.51500000 ;
     RECT 4.65500000 0.44000000 4.94500000 0.51500000 ;
     RECT 0.57500000 0.51500000 4.94500000 0.65500000 ;
     RECT 0.57500000 0.65500000 0.86500000 0.73000000 ;
     RECT 4.65500000 0.65500000 4.94500000 0.73000000 ;
     RECT 0.65000000 0.73000000 0.79000000 2.19500000 ;
     RECT 0.57500000 2.19500000 0.86500000 2.48500000 ;
     RECT 2.25500000 2.19500000 2.54500000 2.27000000 ;
     RECT 4.65500000 2.19500000 4.94500000 2.27000000 ;
     RECT 2.25500000 2.27000000 4.94500000 2.41000000 ;
     RECT 2.25500000 2.41000000 2.54500000 2.48500000 ;
     RECT 4.65500000 2.41000000 4.94500000 2.48500000 ;
     RECT 3.21500000 2.76000000 3.50500000 3.09000000 ;
     RECT 0.00000000 3.09000000 5.76000000 3.57000000 ;

 END
END AOI21X1
