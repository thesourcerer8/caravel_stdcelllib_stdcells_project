VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 15.840 3.570 ;
        RECT 1.780 3.060 2.070 3.090 ;
        RECT 1.780 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.070 3.060 ;
        RECT 1.780 2.830 2.070 2.890 ;
        RECT 4.660 3.060 4.950 3.090 ;
        RECT 4.660 2.890 4.720 3.060 ;
        RECT 4.890 2.890 4.950 3.060 ;
        RECT 7.780 3.020 7.840 3.090 ;
        RECT 8.010 3.020 8.070 3.090 ;
        RECT 7.780 2.960 8.070 3.020 ;
        RECT 11.860 3.060 12.150 3.090 ;
        RECT 4.660 2.830 4.950 2.890 ;
        RECT 11.860 2.890 11.920 3.060 ;
        RECT 12.090 2.890 12.150 3.060 ;
        RECT 11.860 2.830 12.150 2.890 ;
        RECT 13.540 3.060 13.830 3.090 ;
        RECT 13.540 2.890 13.600 3.060 ;
        RECT 13.770 2.890 13.830 3.060 ;
        RECT 13.540 2.830 13.830 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.360 2.070 0.420 ;
        RECT 1.780 0.240 1.840 0.360 ;
        RECT 2.010 0.240 2.070 0.360 ;
        RECT 6.100 0.240 6.390 0.280 ;
        RECT 7.780 0.240 8.070 0.280 ;
        RECT 13.540 0.240 13.830 0.280 ;
        RECT 0.000 -0.240 15.840 0.240 ;
    END
  END gnd
  PIN YS
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 14.740 2.150 15.030 2.440 ;
        RECT 14.810 0.690 14.950 2.150 ;
        RECT 14.740 0.400 15.030 0.690 ;
    END
  END YS
  PIN YC
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.150 0.870 2.440 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
    END
  END YC
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 1.750 5.910 2.040 ;
        RECT 5.690 1.090 5.830 1.750 ;
        RECT 5.620 0.800 5.910 1.090 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.750 4.470 2.040 ;
        RECT 9.940 1.750 10.230 2.040 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 10.010 1.090 10.150 1.750 ;
        RECT 4.180 0.800 4.470 1.090 ;
        RECT 9.940 0.800 10.230 1.090 ;
        RECT 4.250 0.610 4.390 0.800 ;
        RECT 10.010 0.610 10.150 0.800 ;
        RECT 4.250 0.470 10.150 0.610 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 1.760 3.060 2.090 3.140 ;
        RECT 1.760 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.090 3.060 ;
        RECT 1.760 2.810 2.090 2.890 ;
        RECT 4.640 3.060 4.970 3.140 ;
        RECT 4.640 2.890 4.720 3.060 ;
        RECT 4.890 2.890 4.970 3.060 ;
        RECT 4.640 2.810 4.970 2.890 ;
        RECT 7.760 2.890 7.840 3.140 ;
        RECT 8.010 2.890 8.090 3.140 ;
        RECT 7.760 2.810 8.090 2.890 ;
        RECT 11.840 3.060 12.170 3.140 ;
        RECT 11.840 2.890 11.920 3.060 ;
        RECT 12.090 2.890 12.170 3.060 ;
        RECT 11.840 2.810 12.170 2.890 ;
        RECT 13.520 3.060 13.850 3.140 ;
        RECT 13.520 2.890 13.600 3.060 ;
        RECT 13.770 2.890 13.850 3.060 ;
        RECT 13.520 2.810 13.850 2.890 ;
        RECT 0.560 2.380 0.890 2.460 ;
        RECT 0.560 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.890 2.380 ;
        RECT 0.560 2.130 0.890 2.210 ;
        RECT 3.440 2.380 3.770 2.460 ;
        RECT 3.440 2.210 3.520 2.380 ;
        RECT 3.690 2.210 3.770 2.380 ;
        RECT 3.440 2.130 3.770 2.210 ;
        RECT 5.680 2.060 5.850 2.620 ;
        RECT 6.080 2.380 6.410 2.460 ;
        RECT 6.080 2.210 6.160 2.380 ;
        RECT 6.330 2.210 6.410 2.380 ;
        RECT 6.080 2.130 6.410 2.210 ;
        RECT 9.440 2.380 9.770 2.460 ;
        RECT 9.440 2.210 9.520 2.380 ;
        RECT 9.690 2.230 9.770 2.380 ;
        RECT 14.720 2.380 15.050 2.460 ;
        RECT 14.720 2.230 14.800 2.380 ;
        RECT 9.690 2.210 9.750 2.230 ;
        RECT 9.440 2.130 9.750 2.210 ;
        RECT 14.740 2.210 14.800 2.230 ;
        RECT 14.970 2.210 15.050 2.380 ;
        RECT 14.740 2.130 15.050 2.210 ;
        RECT 1.280 1.980 1.610 2.060 ;
        RECT 1.280 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 4.160 1.980 4.490 2.060 ;
        RECT 4.160 1.810 4.240 1.980 ;
        RECT 4.410 1.810 4.490 1.980 ;
        RECT 4.160 1.730 4.490 1.810 ;
        RECT 5.600 1.980 5.910 2.060 ;
        RECT 5.600 1.810 5.680 1.980 ;
        RECT 5.850 1.960 5.910 1.980 ;
        RECT 8.480 1.980 8.810 2.060 ;
        RECT 5.850 1.810 5.930 1.960 ;
        RECT 5.600 1.730 5.930 1.810 ;
        RECT 8.480 1.810 8.560 1.980 ;
        RECT 8.730 1.810 8.810 1.980 ;
        RECT 8.480 1.730 8.810 1.810 ;
        RECT 9.920 1.980 10.250 2.060 ;
        RECT 9.920 1.810 10.000 1.980 ;
        RECT 10.170 1.810 10.250 1.980 ;
        RECT 9.920 1.730 10.250 1.810 ;
        RECT 11.360 1.980 11.690 2.060 ;
        RECT 11.360 1.810 11.440 1.980 ;
        RECT 11.610 1.810 11.690 1.980 ;
        RECT 11.360 1.730 11.690 1.810 ;
        RECT 14.240 1.980 14.570 2.060 ;
        RECT 14.240 1.810 14.320 1.980 ;
        RECT 14.490 1.810 14.570 1.980 ;
        RECT 14.240 1.730 14.570 1.810 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.860 1.360 1.030 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.280 0.780 1.610 0.860 ;
        RECT 4.160 1.030 4.490 1.110 ;
        RECT 4.160 0.860 4.240 1.030 ;
        RECT 4.410 0.860 4.490 1.030 ;
        RECT 4.160 0.780 4.490 0.860 ;
        RECT 5.600 1.030 5.930 1.110 ;
        RECT 5.600 0.860 5.680 1.030 ;
        RECT 5.850 0.860 5.930 1.030 ;
        RECT 5.600 0.780 5.930 0.860 ;
        RECT 8.480 1.030 8.810 1.110 ;
        RECT 8.480 0.860 8.560 1.030 ;
        RECT 8.730 0.860 8.810 1.030 ;
        RECT 8.480 0.780 8.810 0.860 ;
        RECT 9.920 1.030 10.250 1.110 ;
        RECT 9.920 0.860 10.000 1.030 ;
        RECT 10.170 0.860 10.250 1.030 ;
        RECT 9.920 0.780 10.250 0.860 ;
        RECT 11.360 1.030 11.690 1.110 ;
        RECT 11.360 0.860 11.440 1.030 ;
        RECT 11.610 0.860 11.690 1.030 ;
        RECT 11.360 0.780 11.690 0.860 ;
        RECT 14.240 1.030 14.570 1.110 ;
        RECT 14.240 0.860 14.320 1.030 ;
        RECT 14.490 0.880 14.570 1.030 ;
        RECT 14.490 0.860 14.550 0.880 ;
        RECT 14.240 0.780 14.550 0.860 ;
        RECT 0.560 0.630 0.890 0.710 ;
        RECT 0.560 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.890 0.630 ;
        RECT 0.560 0.380 0.890 0.460 ;
        RECT 3.440 0.630 3.770 0.710 ;
        RECT 3.440 0.460 3.520 0.630 ;
        RECT 3.690 0.460 3.770 0.630 ;
        RECT 10.420 0.630 10.730 0.710 ;
        RECT 10.420 0.610 10.480 0.630 ;
        RECT 1.760 0.360 2.090 0.440 ;
        RECT 3.440 0.380 3.770 0.460 ;
        RECT 10.400 0.460 10.480 0.610 ;
        RECT 10.650 0.460 10.730 0.630 ;
        RECT 1.760 0.190 1.840 0.360 ;
        RECT 2.010 0.190 2.090 0.360 ;
        RECT 1.760 0.110 2.090 0.190 ;
        RECT 6.080 0.360 6.410 0.440 ;
        RECT 6.080 0.110 6.160 0.360 ;
        RECT 6.330 0.110 6.410 0.360 ;
        RECT 7.760 0.360 8.090 0.440 ;
        RECT 7.760 0.110 7.840 0.360 ;
        RECT 8.010 0.110 8.090 0.360 ;
        RECT 9.440 0.360 9.770 0.440 ;
        RECT 10.400 0.390 10.730 0.460 ;
        RECT 14.720 0.630 15.050 0.710 ;
        RECT 14.720 0.460 14.800 0.630 ;
        RECT 14.970 0.460 15.050 0.630 ;
        RECT 9.440 0.190 9.520 0.360 ;
        RECT 9.690 0.220 9.770 0.360 ;
        RECT 11.840 0.360 12.170 0.440 ;
        RECT 11.840 0.220 11.920 0.360 ;
        RECT 9.690 0.190 11.920 0.220 ;
        RECT 12.090 0.190 12.170 0.360 ;
        RECT 9.440 0.110 12.170 0.190 ;
        RECT 13.520 0.360 13.850 0.440 ;
        RECT 14.720 0.380 15.050 0.460 ;
        RECT 13.520 0.110 13.600 0.360 ;
        RECT 13.770 0.110 13.850 0.360 ;
        RECT 9.520 0.050 12.090 0.110 ;
      LAYER met1 ;
        RECT 5.620 2.790 5.910 2.850 ;
        RECT 5.620 2.620 5.680 2.790 ;
        RECT 5.850 2.770 5.910 2.790 ;
        RECT 5.850 2.630 11.590 2.770 ;
        RECT 5.850 2.620 5.910 2.630 ;
        RECT 5.620 2.560 5.910 2.620 ;
        RECT 3.460 2.380 3.750 2.440 ;
        RECT 3.460 2.210 3.520 2.380 ;
        RECT 3.690 2.370 3.750 2.380 ;
        RECT 6.100 2.380 6.390 2.440 ;
        RECT 6.100 2.370 6.160 2.380 ;
        RECT 3.690 2.230 6.160 2.370 ;
        RECT 3.690 2.210 3.750 2.230 ;
        RECT 3.460 2.150 3.750 2.210 ;
        RECT 6.100 2.210 6.160 2.230 ;
        RECT 6.330 2.370 6.390 2.380 ;
        RECT 9.460 2.380 9.750 2.440 ;
        RECT 6.330 2.230 8.710 2.370 ;
        RECT 6.330 2.210 6.390 2.230 ;
        RECT 6.100 2.150 6.390 2.210 ;
        RECT 1.300 1.980 1.590 2.040 ;
        RECT 1.300 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.590 1.980 ;
        RECT 1.300 1.750 1.590 1.810 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 1.030 1.590 1.090 ;
        RECT 1.300 0.860 1.360 1.030 ;
        RECT 1.530 1.020 1.590 1.030 ;
        RECT 3.530 1.020 3.670 2.150 ;
        RECT 8.570 2.040 8.710 2.230 ;
        RECT 9.460 2.210 9.520 2.380 ;
        RECT 9.690 2.370 9.750 2.380 ;
        RECT 9.690 2.230 10.630 2.370 ;
        RECT 9.690 2.210 9.750 2.230 ;
        RECT 9.460 2.150 9.750 2.210 ;
        RECT 8.500 1.980 8.790 2.040 ;
        RECT 8.500 1.810 8.560 1.980 ;
        RECT 8.730 1.810 8.790 1.980 ;
        RECT 8.500 1.750 8.790 1.810 ;
        RECT 8.570 1.090 8.710 1.750 ;
        RECT 1.530 0.880 3.670 1.020 ;
        RECT 1.530 0.860 1.590 0.880 ;
        RECT 1.300 0.800 1.590 0.860 ;
        RECT 3.530 0.690 3.670 0.880 ;
        RECT 8.500 1.030 8.790 1.090 ;
        RECT 8.500 0.860 8.560 1.030 ;
        RECT 8.730 0.860 8.790 1.030 ;
        RECT 8.500 0.800 8.790 0.860 ;
        RECT 10.490 0.690 10.630 2.230 ;
        RECT 11.450 2.040 11.590 2.630 ;
        RECT 11.380 1.980 11.670 2.040 ;
        RECT 11.380 1.810 11.440 1.980 ;
        RECT 11.610 1.810 11.670 1.980 ;
        RECT 11.380 1.750 11.670 1.810 ;
        RECT 14.260 1.980 14.550 2.040 ;
        RECT 14.260 1.810 14.320 1.980 ;
        RECT 14.490 1.810 14.550 1.980 ;
        RECT 14.260 1.750 14.550 1.810 ;
        RECT 11.450 1.090 11.590 1.750 ;
        RECT 14.330 1.090 14.470 1.750 ;
        RECT 11.380 1.030 11.670 1.090 ;
        RECT 11.380 0.860 11.440 1.030 ;
        RECT 11.610 0.860 11.670 1.030 ;
        RECT 11.380 0.800 11.670 0.860 ;
        RECT 14.260 1.030 14.550 1.090 ;
        RECT 14.260 0.860 14.320 1.030 ;
        RECT 14.490 0.860 14.550 1.030 ;
        RECT 14.260 0.800 14.550 0.860 ;
        RECT 3.460 0.630 3.750 0.690 ;
        RECT 3.460 0.460 3.520 0.630 ;
        RECT 3.690 0.460 3.750 0.630 ;
        RECT 3.460 0.400 3.750 0.460 ;
        RECT 10.420 0.630 10.710 0.690 ;
        RECT 10.420 0.460 10.480 0.630 ;
        RECT 10.650 0.610 10.710 0.630 ;
        RECT 14.330 0.610 14.470 0.800 ;
        RECT 10.650 0.470 14.470 0.610 ;
        RECT 10.650 0.460 10.710 0.470 ;
        RECT 10.420 0.400 10.710 0.460 ;
  END
END HAX1
END LIBRARY

