VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.840 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 5.615 1.780 5.905 2.070 ;
        RECT 11.375 1.780 11.665 2.070 ;
        RECT 5.690 1.135 5.830 1.780 ;
        RECT 11.450 1.135 11.590 1.780 ;
        RECT 5.615 1.060 5.905 1.135 ;
        RECT 11.375 1.060 11.665 1.135 ;
        RECT 5.615 0.920 11.665 1.060 ;
        RECT 5.615 0.845 5.905 0.920 ;
        RECT 11.375 0.845 11.665 0.920 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 4.175 2.815 4.465 2.890 ;
        RECT 4.175 2.675 10.150 2.815 ;
        RECT 4.175 2.600 4.465 2.675 ;
        RECT 10.010 2.070 10.150 2.675 ;
        RECT 4.175 1.780 4.465 2.070 ;
        RECT 9.935 1.780 10.225 2.070 ;
        RECT 4.250 1.135 4.390 1.780 ;
        RECT 4.175 0.845 4.465 1.135 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 1.408400 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 6.095 0.440 6.385 0.730 ;
        RECT 7.775 0.440 8.065 0.730 ;
        RECT 13.535 0.440 13.825 0.730 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 6.170 0.240 6.310 0.440 ;
        RECT 7.850 0.240 7.990 0.440 ;
        RECT 13.610 0.240 13.750 0.440 ;
        RECT 0.000 -0.240 15.840 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 15.840 3.570 ;
        RECT 1.775 2.735 2.065 3.090 ;
        RECT 11.855 2.735 12.145 3.090 ;
        RECT 13.535 2.735 13.825 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 3.074400 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 15.840 3.415 ;
        RECT 0.155 3.215 15.685 3.245 ;
        RECT 0.155 3.090 11.665 3.215 ;
        RECT 12.335 3.090 15.685 3.215 ;
        RECT 1.755 2.715 2.085 3.090 ;
        RECT 4.635 2.715 4.965 3.090 ;
        RECT 7.755 2.715 8.085 3.090 ;
        RECT 13.515 2.715 13.845 3.090 ;
      LAYER mcon ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 3.035 3.245 3.205 3.415 ;
        RECT 3.515 3.245 3.685 3.415 ;
        RECT 3.995 3.245 4.165 3.415 ;
        RECT 4.475 3.245 4.645 3.415 ;
        RECT 4.955 3.245 5.125 3.415 ;
        RECT 5.435 3.245 5.605 3.415 ;
        RECT 5.915 3.245 6.085 3.415 ;
        RECT 6.395 3.245 6.565 3.415 ;
        RECT 6.875 3.245 7.045 3.415 ;
        RECT 7.355 3.245 7.525 3.415 ;
        RECT 7.835 3.245 8.005 3.415 ;
        RECT 8.315 3.245 8.485 3.415 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 9.275 3.245 9.445 3.415 ;
        RECT 9.755 3.245 9.925 3.415 ;
        RECT 10.235 3.245 10.405 3.415 ;
        RECT 10.715 3.245 10.885 3.415 ;
        RECT 11.195 3.245 11.365 3.415 ;
        RECT 11.675 3.245 11.845 3.415 ;
        RECT 12.155 3.245 12.325 3.415 ;
        RECT 12.635 3.245 12.805 3.415 ;
        RECT 13.115 3.245 13.285 3.415 ;
        RECT 13.595 3.245 13.765 3.415 ;
        RECT 14.075 3.245 14.245 3.415 ;
        RECT 14.555 3.245 14.725 3.415 ;
        RECT 15.035 3.245 15.205 3.415 ;
        RECT 1.835 2.795 2.005 2.965 ;
        RECT 13.595 2.795 13.765 2.965 ;
    END
  END VPWR
  PIN YC
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 0.650 0.730 0.790 2.195 ;
        RECT 0.575 0.440 0.865 0.730 ;
    END
  END YC
  PIN YS
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 14.735 2.195 15.025 2.485 ;
        RECT 14.810 0.730 14.950 2.195 ;
        RECT 14.735 0.440 15.025 0.730 ;
    END
  END YS
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 15.840 3.330 ;
      LAYER li1 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 3.435 2.175 3.765 2.505 ;
        RECT 4.235 2.090 4.405 2.830 ;
        RECT 11.835 2.715 12.165 3.045 ;
        RECT 6.075 2.260 6.405 2.505 ;
        RECT 6.095 2.175 6.405 2.260 ;
        RECT 9.435 2.260 9.765 2.505 ;
        RECT 14.715 2.260 15.045 2.505 ;
        RECT 9.435 2.175 9.745 2.260 ;
        RECT 14.735 2.175 15.045 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 4.155 1.760 4.485 2.090 ;
        RECT 5.595 1.760 5.925 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 9.915 1.760 10.245 2.090 ;
        RECT 11.355 1.760 11.685 2.090 ;
        RECT 14.235 1.760 14.565 2.090 ;
        RECT 8.555 1.155 8.725 1.760 ;
        RECT 9.995 1.155 10.165 1.760 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 4.155 0.825 4.485 1.155 ;
        RECT 5.595 0.825 5.925 1.155 ;
        RECT 8.475 0.825 8.805 1.155 ;
        RECT 9.915 0.920 10.245 1.155 ;
        RECT 9.935 0.825 10.225 0.920 ;
        RECT 10.475 0.750 10.645 1.480 ;
        RECT 11.355 0.920 11.685 1.155 ;
        RECT 14.235 0.920 14.565 1.155 ;
        RECT 11.355 0.825 11.665 0.920 ;
        RECT 14.235 0.825 14.545 0.920 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.435 0.420 3.765 0.750 ;
        RECT 6.095 0.655 6.405 0.750 ;
        RECT 6.075 0.420 6.405 0.655 ;
        RECT 7.755 0.420 8.085 0.750 ;
        RECT 9.435 0.420 9.765 0.750 ;
        RECT 10.395 0.420 10.725 0.750 ;
        RECT 11.835 0.420 12.165 0.750 ;
        RECT 13.515 0.420 13.845 0.750 ;
        RECT 14.715 0.420 15.045 0.750 ;
        RECT 0.155 0.085 15.685 0.240 ;
        RECT 0.000 -0.085 15.840 0.085 ;
      LAYER mcon ;
        RECT 4.235 2.660 4.405 2.830 ;
        RECT 11.915 2.795 12.085 2.965 ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 3.515 2.255 3.685 2.425 ;
        RECT 6.155 2.255 6.325 2.425 ;
        RECT 9.515 2.255 9.685 2.425 ;
        RECT 14.795 2.255 14.965 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 4.235 1.840 4.405 2.010 ;
        RECT 5.675 1.840 5.845 2.010 ;
        RECT 8.555 1.840 8.725 2.010 ;
        RECT 9.995 1.840 10.165 2.010 ;
        RECT 11.435 1.840 11.605 2.010 ;
        RECT 14.315 1.840 14.485 2.010 ;
        RECT 10.475 1.310 10.645 1.480 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 11.435 0.905 11.605 1.075 ;
        RECT 14.315 0.905 14.485 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.515 0.500 3.685 0.670 ;
        RECT 6.155 0.500 6.325 0.670 ;
        RECT 7.835 0.500 8.005 0.670 ;
        RECT 9.515 0.500 9.685 0.670 ;
        RECT 11.915 0.500 12.085 0.670 ;
        RECT 13.595 0.500 13.765 0.670 ;
        RECT 14.795 0.500 14.965 0.670 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
        RECT 3.035 -0.085 3.205 0.085 ;
        RECT 3.515 -0.085 3.685 0.085 ;
        RECT 3.995 -0.085 4.165 0.085 ;
        RECT 4.475 -0.085 4.645 0.085 ;
        RECT 4.955 -0.085 5.125 0.085 ;
        RECT 5.435 -0.085 5.605 0.085 ;
        RECT 5.915 -0.085 6.085 0.085 ;
        RECT 6.395 -0.085 6.565 0.085 ;
        RECT 6.875 -0.085 7.045 0.085 ;
        RECT 7.355 -0.085 7.525 0.085 ;
        RECT 7.835 -0.085 8.005 0.085 ;
        RECT 8.315 -0.085 8.485 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.275 -0.085 9.445 0.085 ;
        RECT 9.755 -0.085 9.925 0.085 ;
        RECT 10.235 -0.085 10.405 0.085 ;
        RECT 10.715 -0.085 10.885 0.085 ;
        RECT 11.195 -0.085 11.365 0.085 ;
        RECT 11.675 -0.085 11.845 0.085 ;
        RECT 12.155 -0.085 12.325 0.085 ;
        RECT 12.635 -0.085 12.805 0.085 ;
        RECT 13.115 -0.085 13.285 0.085 ;
        RECT 13.595 -0.085 13.765 0.085 ;
        RECT 14.075 -0.085 14.245 0.085 ;
        RECT 14.555 -0.085 14.725 0.085 ;
        RECT 15.035 -0.085 15.205 0.085 ;
      LAYER met1 ;
        RECT 3.455 2.410 3.745 2.485 ;
        RECT 6.095 2.410 6.385 2.485 ;
        RECT 3.455 2.270 8.710 2.410 ;
        RECT 3.455 2.195 3.745 2.270 ;
        RECT 6.095 2.195 6.385 2.270 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 1.060 1.585 1.135 ;
        RECT 3.530 1.060 3.670 2.195 ;
        RECT 8.570 2.070 8.710 2.270 ;
        RECT 9.455 2.195 9.745 2.485 ;
        RECT 10.490 2.270 14.470 2.410 ;
        RECT 8.495 1.780 8.785 2.070 ;
        RECT 9.530 1.465 9.670 2.195 ;
        RECT 10.490 1.540 10.630 2.270 ;
        RECT 14.330 2.070 14.470 2.270 ;
        RECT 14.255 1.780 14.545 2.070 ;
        RECT 10.415 1.465 10.705 1.540 ;
        RECT 9.530 1.325 10.705 1.465 ;
        RECT 10.415 1.250 10.705 1.325 ;
        RECT 14.330 1.135 14.470 1.780 ;
        RECT 1.295 0.920 3.670 1.060 ;
        RECT 1.295 0.845 1.585 0.920 ;
        RECT 3.530 0.730 3.670 0.920 ;
        RECT 14.255 0.845 14.545 1.135 ;
        RECT 3.455 0.440 3.745 0.730 ;
        RECT 9.455 0.655 9.745 0.730 ;
        RECT 11.855 0.655 12.145 0.730 ;
        RECT 9.455 0.515 12.145 0.655 ;
        RECT 9.455 0.440 9.745 0.515 ;
        RECT 11.855 0.440 12.145 0.515 ;
  END
END HAX1
END LIBRARY

