VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OAI21X1
  CLASS CORE ;
  FOREIGN OAI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.760 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 5.760 3.570 ;
        RECT 1.780 3.060 2.070 3.090 ;
        RECT 1.780 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.070 3.060 ;
        RECT 1.780 2.830 2.070 2.890 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.220 0.240 3.510 0.280 ;
        RECT 0.000 -0.240 5.760 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.370 0.870 2.440 ;
        RECT 4.660 2.370 4.950 2.440 ;
        RECT 0.580 2.230 4.950 2.370 ;
        RECT 0.580 2.150 0.870 2.230 ;
        RECT 4.660 2.150 4.950 2.230 ;
        RECT 0.650 0.690 0.790 2.150 ;
        RECT 0.580 0.400 0.870 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.750 3.030 2.040 ;
        RECT 2.810 1.090 2.950 1.750 ;
        RECT 2.740 0.800 3.030 1.090 ;
    END
  END A
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.750 1.590 2.040 ;
        RECT 1.370 1.090 1.510 1.750 ;
        RECT 1.300 0.800 1.590 1.090 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 4.180 1.750 4.470 2.040 ;
        RECT 4.250 1.090 4.390 1.750 ;
        RECT 4.180 0.800 4.470 1.090 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 1.760 3.060 2.090 3.140 ;
        RECT 1.760 2.890 1.840 3.060 ;
        RECT 2.010 2.890 2.090 3.060 ;
        RECT 1.760 2.810 2.090 2.890 ;
        RECT 0.560 2.380 0.890 2.460 ;
        RECT 0.560 2.210 0.640 2.380 ;
        RECT 0.810 2.210 0.890 2.380 ;
        RECT 0.560 2.130 0.890 2.210 ;
        RECT 4.640 2.380 4.970 2.460 ;
        RECT 4.640 2.210 4.720 2.380 ;
        RECT 4.890 2.210 4.970 2.380 ;
        RECT 4.640 2.130 4.970 2.210 ;
        RECT 1.280 1.980 1.610 2.060 ;
        RECT 1.280 1.810 1.360 1.980 ;
        RECT 1.530 1.810 1.610 1.980 ;
        RECT 1.280 1.730 1.610 1.810 ;
        RECT 2.720 1.980 3.050 2.060 ;
        RECT 2.720 1.810 2.800 1.980 ;
        RECT 2.970 1.810 3.050 1.980 ;
        RECT 2.720 1.730 3.050 1.810 ;
        RECT 4.160 1.980 4.470 2.060 ;
        RECT 4.160 1.810 4.240 1.980 ;
        RECT 4.410 1.960 4.470 1.980 ;
        RECT 4.410 1.810 4.490 1.960 ;
        RECT 4.160 1.730 4.490 1.810 ;
        RECT 1.280 1.030 1.610 1.110 ;
        RECT 1.280 0.860 1.360 1.030 ;
        RECT 1.530 0.860 1.610 1.030 ;
        RECT 1.280 0.780 1.610 0.860 ;
        RECT 2.720 1.030 3.050 1.110 ;
        RECT 2.720 0.860 2.800 1.030 ;
        RECT 2.970 0.860 3.050 1.030 ;
        RECT 2.720 0.780 3.050 0.860 ;
        RECT 4.160 1.030 4.490 1.110 ;
        RECT 4.160 0.860 4.240 1.030 ;
        RECT 4.410 0.880 4.490 1.030 ;
        RECT 4.410 0.860 4.470 0.880 ;
        RECT 4.160 0.780 4.470 0.860 ;
        RECT 0.560 0.630 0.890 0.710 ;
        RECT 0.560 0.460 0.640 0.630 ;
        RECT 0.810 0.460 0.890 0.630 ;
        RECT 0.560 0.380 0.890 0.460 ;
        RECT 2.240 0.630 2.550 0.710 ;
        RECT 2.240 0.460 2.320 0.630 ;
        RECT 2.490 0.610 2.550 0.630 ;
        RECT 4.640 0.630 4.970 0.710 ;
        RECT 2.490 0.460 2.570 0.610 ;
        RECT 2.240 0.380 2.570 0.460 ;
        RECT 4.640 0.460 4.720 0.630 ;
        RECT 4.890 0.460 4.970 0.630 ;
        RECT 3.200 0.360 3.530 0.440 ;
        RECT 4.640 0.380 4.970 0.460 ;
        RECT 3.200 0.110 3.280 0.360 ;
        RECT 3.450 0.110 3.530 0.360 ;
      LAYER met1 ;
        RECT 2.260 0.630 2.550 0.690 ;
        RECT 2.260 0.460 2.320 0.630 ;
        RECT 2.490 0.610 2.550 0.630 ;
        RECT 4.660 0.630 4.950 0.690 ;
        RECT 4.660 0.610 4.720 0.630 ;
        RECT 2.490 0.470 4.720 0.610 ;
        RECT 2.490 0.460 2.550 0.470 ;
        RECT 2.260 0.400 2.550 0.460 ;
        RECT 4.660 0.460 4.720 0.470 ;
        RECT 4.890 0.460 4.950 0.630 ;
        RECT 4.660 0.400 4.950 0.460 ;
  END
END OAI21X1
END LIBRARY

