VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 1.780 2.990 2.070 3.090 ;
        RECT 1.780 2.820 1.840 2.990 ;
        RECT 2.010 2.820 2.070 2.990 ;
        RECT 1.780 2.760 2.070 2.820 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 1.760 2.990 2.090 3.090 ;
        RECT 1.760 2.820 1.840 2.990 ;
        RECT 2.010 2.820 2.090 2.990 ;
        RECT 1.760 2.740 2.090 2.820 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.510 2.070 0.570 ;
        RECT 1.780 0.340 1.840 0.510 ;
        RECT 2.010 0.340 2.070 0.510 ;
        RECT 1.780 0.240 2.070 0.340 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.760 0.510 2.090 0.590 ;
        RECT 1.760 0.340 1.840 0.510 ;
        RECT 2.010 0.340 2.090 0.510 ;
        RECT 1.760 0.260 2.090 0.340 ;
        RECT 1.590 0.240 2.260 0.260 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.410 0.870 2.490 ;
        RECT 3.220 2.410 3.510 2.490 ;
        RECT 0.580 2.270 3.510 2.410 ;
        RECT 0.580 2.200 0.870 2.270 ;
        RECT 3.220 2.200 3.510 2.270 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 3.290 0.730 3.430 2.200 ;
        RECT 0.580 0.440 0.870 0.730 ;
        RECT 3.220 0.440 3.510 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 2.000 1.590 2.070 ;
        RECT 2.740 2.000 3.030 2.070 ;
        RECT 1.300 1.860 3.030 2.000 ;
        RECT 1.300 1.780 1.590 1.860 ;
        RECT 2.740 1.780 3.030 1.860 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 2.810 1.140 2.950 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
        RECT 2.740 0.850 3.030 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 3.200 2.430 3.530 2.510 ;
        RECT 3.200 2.260 3.280 2.430 ;
        RECT 3.450 2.260 3.530 2.430 ;
        RECT 3.200 2.180 3.530 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.030 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.920 3.050 1.080 ;
        RECT 2.970 0.910 3.030 0.920 ;
        RECT 2.720 0.830 3.030 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 3.200 0.670 3.530 0.750 ;
        RECT 3.200 0.500 3.280 0.670 ;
        RECT 3.450 0.500 3.530 0.670 ;
        RECT 3.200 0.420 3.530 0.500 ;
  END
END INVX4
END LIBRARY

