VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.275 1.760 1.605 2.090 ;
      LAYER mcon ;
        RECT 1.355 1.840 1.525 2.010 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 0.331800 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.240 2.065 0.570 ;
        RECT 0.000 -0.240 2.880 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.755 0.240 2.085 0.590 ;
        RECT 0.155 0.085 2.725 0.240 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 1.835 0.340 2.005 0.510 ;
        RECT 0.155 -0.085 0.325 0.085 ;
        RECT 0.635 -0.085 0.805 0.085 ;
        RECT 1.115 -0.085 1.285 0.085 ;
        RECT 1.595 -0.085 1.765 0.085 ;
        RECT 2.075 -0.085 2.245 0.085 ;
        RECT 2.555 -0.085 2.725 0.085 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 2.880 3.570 ;
        RECT 1.775 2.760 2.065 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 0.663600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 2.880 3.415 ;
        RECT 0.155 3.090 2.725 3.245 ;
        RECT 1.755 2.740 2.085 3.090 ;
      LAYER mcon ;
        RECT 0.155 3.245 0.325 3.415 ;
        RECT 0.635 3.245 0.805 3.415 ;
        RECT 1.115 3.245 1.285 3.415 ;
        RECT 1.595 3.245 1.765 3.415 ;
        RECT 2.075 3.245 2.245 3.415 ;
        RECT 2.555 3.245 2.725 3.415 ;
        RECT 1.835 2.820 2.005 2.990 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 0.650 0.730 0.790 2.195 ;
        RECT 0.575 0.440 0.865 0.730 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.555 2.175 0.885 2.505 ;
      LAYER mcon ;
        RECT 0.635 2.255 0.805 2.425 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 2.880 3.330 ;
      LAYER li1 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
      LAYER mcon ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
  END
END INVX2
END LIBRARY

