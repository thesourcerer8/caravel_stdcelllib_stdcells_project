magic
tech sky130A
magscale 1 2
timestamp 1624917760
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 2592 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
rect 1425 48 1455 132
rect 1713 48 1743 132
rect 2001 48 2031 132
rect 2289 48 2319 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
rect 1425 450 1455 618
rect 1713 450 1743 618
rect 2001 450 2031 618
rect 2289 450 2319 618
<< ndiff >>
rect 355 134 413 146
rect 355 132 367 134
rect 115 102 273 132
rect 115 68 127 102
rect 161 68 273 102
rect 115 48 273 68
rect 303 100 367 132
rect 401 132 413 134
rect 931 134 989 146
rect 931 132 943 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 102 849 132
rect 591 68 655 102
rect 689 68 849 102
rect 591 48 849 68
rect 879 100 943 132
rect 977 132 989 134
rect 1507 134 1565 146
rect 1507 132 1519 134
rect 977 100 1137 132
rect 879 48 1137 100
rect 1167 102 1425 132
rect 1167 68 1231 102
rect 1265 68 1425 102
rect 1167 48 1425 68
rect 1455 100 1519 132
rect 1553 132 1565 134
rect 2083 134 2141 146
rect 2083 132 2095 134
rect 1553 100 1713 132
rect 1455 48 1713 100
rect 1743 102 2001 132
rect 1743 68 1807 102
rect 1841 68 2001 102
rect 1743 48 2001 68
rect 2031 100 2095 132
rect 2129 132 2141 134
rect 2129 100 2289 132
rect 2031 48 2289 100
rect 2319 102 2477 132
rect 2319 68 2383 102
rect 2417 68 2477 102
rect 2319 48 2477 68
<< pdiff >>
rect 115 598 273 618
rect 115 564 127 598
rect 161 564 273 598
rect 115 450 273 564
rect 303 485 561 618
rect 303 451 367 485
rect 401 451 561 485
rect 303 450 561 451
rect 591 598 849 618
rect 591 564 655 598
rect 689 564 849 598
rect 591 450 849 564
rect 879 485 1137 618
rect 879 451 943 485
rect 977 451 1137 485
rect 879 450 1137 451
rect 1167 598 1425 618
rect 1167 564 1231 598
rect 1265 564 1425 598
rect 1167 450 1425 564
rect 1455 485 1713 618
rect 1455 451 1519 485
rect 1553 451 1713 485
rect 1455 450 1713 451
rect 1743 598 2001 618
rect 1743 564 1807 598
rect 1841 564 2001 598
rect 1743 450 2001 564
rect 2031 485 2289 618
rect 2031 451 2095 485
rect 2129 451 2289 485
rect 2031 450 2289 451
rect 2319 598 2477 618
rect 2319 564 2383 598
rect 2417 564 2477 598
rect 2319 450 2477 564
rect 355 439 413 450
rect 931 439 989 450
rect 1507 439 1565 450
rect 2083 439 2141 450
<< ndiffc >>
rect 127 68 161 102
rect 367 100 401 134
rect 655 68 689 102
rect 943 100 977 134
rect 1231 68 1265 102
rect 1519 100 1553 134
rect 1807 68 1841 102
rect 2095 100 2129 134
rect 2383 68 2417 102
<< pdiffc >>
rect 127 564 161 598
rect 367 451 401 485
rect 655 564 689 598
rect 943 451 977 485
rect 1231 564 1265 598
rect 1519 451 1553 485
rect 1807 564 1841 598
rect 2095 451 2129 485
rect 2383 564 2417 598
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 1425 618 1455 644
rect 1713 618 1743 644
rect 2001 618 2031 644
rect 2289 618 2319 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 1425 418 1455 450
rect 1713 418 1743 450
rect 2001 418 2031 450
rect 2289 418 2319 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1473 418
rect 1407 368 1423 402
rect 1457 368 1473 402
rect 1407 352 1473 368
rect 1695 402 1761 418
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 181 1473 215
rect 1407 165 1473 181
rect 1695 215 1761 231
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 181 2049 215
rect 1983 165 2049 181
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 181 2337 215
rect 2271 165 2337 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 1425 132 1455 165
rect 1713 132 1743 165
rect 2001 132 2031 165
rect 2289 132 2319 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
rect 1425 22 1455 48
rect 1713 22 1743 48
rect 2001 22 2031 48
rect 2289 22 2319 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 1423 368 1457 402
rect 1711 368 1745 402
rect 1999 368 2033 402
rect 2287 368 2321 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 2287 181 2321 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 31 618 2561 649
rect 111 598 177 618
rect 111 564 127 598
rect 161 564 177 598
rect 111 548 177 564
rect 639 598 705 618
rect 639 564 655 598
rect 689 564 705 598
rect 1215 598 1281 618
rect 639 548 705 564
rect 1215 564 1231 598
rect 1265 564 1281 598
rect 1791 598 1857 618
rect 1215 548 1281 564
rect 351 485 417 501
rect 351 452 367 485
rect 355 451 367 452
rect 401 451 417 485
rect 927 485 993 501
rect 927 452 943 485
rect 355 435 417 451
rect 931 451 943 452
rect 977 451 993 485
rect 931 435 993 451
rect 1135 418 1169 532
rect 1791 564 1807 598
rect 1841 564 1857 598
rect 1791 548 1857 564
rect 2367 598 2433 618
rect 2367 564 2383 598
rect 2417 564 2433 598
rect 2367 548 2433 564
rect 1503 485 1569 501
rect 1503 451 1519 485
rect 1553 451 1569 485
rect 1503 435 1569 451
rect 1711 418 1745 532
rect 2079 485 2145 501
rect 2079 452 2095 485
rect 2083 451 2095 452
rect 2129 451 2145 485
rect 2083 435 2145 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 1407 402 1469 418
rect 1407 368 1423 402
rect 1457 401 1469 402
rect 1695 402 1761 418
rect 1457 368 1473 401
rect 1407 352 1473 368
rect 1695 368 1711 402
rect 1745 368 1761 402
rect 1695 352 1761 368
rect 1983 402 2049 418
rect 1983 368 1999 402
rect 2033 368 2049 402
rect 1983 352 2049 368
rect 1135 323 1169 352
rect 1711 323 1745 352
rect 559 231 593 262
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 184 897 215
rect 1119 215 1185 231
rect 881 181 893 184
rect 831 165 893 181
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 1407 215 1473 231
rect 1407 181 1423 215
rect 1457 184 1473 215
rect 1695 215 1761 231
rect 1457 181 1469 184
rect 1407 165 1469 181
rect 1695 181 1711 215
rect 1745 181 1761 215
rect 1695 165 1761 181
rect 1983 215 2049 231
rect 1983 181 1999 215
rect 2033 184 2049 215
rect 2033 181 2045 184
rect 1983 165 2045 181
rect 2095 150 2129 435
rect 2271 402 2337 418
rect 2271 368 2287 402
rect 2321 368 2337 402
rect 2271 352 2337 368
rect 2271 215 2337 231
rect 2271 181 2287 215
rect 2321 181 2337 215
rect 2271 165 2337 181
rect 355 134 417 150
rect 355 131 367 134
rect 111 102 177 118
rect 111 68 127 102
rect 161 68 177 102
rect 351 100 367 131
rect 401 100 417 134
rect 927 134 993 150
rect 351 84 417 100
rect 639 102 705 118
rect 111 48 177 68
rect 639 68 655 102
rect 689 68 705 102
rect 927 100 943 134
rect 977 100 993 134
rect 1503 134 1569 150
rect 927 84 993 100
rect 1215 102 1281 118
rect 639 48 705 68
rect 1215 68 1231 102
rect 1265 68 1281 102
rect 1503 100 1519 134
rect 1553 100 1569 134
rect 2079 134 2145 150
rect 1503 84 1569 100
rect 1791 102 1857 118
rect 1215 48 1281 68
rect 1791 68 1807 102
rect 1841 68 1857 102
rect 2079 100 2095 134
rect 2129 100 2145 134
rect 2079 84 2145 100
rect 2367 102 2433 118
rect 1791 48 1857 68
rect 2367 68 2383 102
rect 2417 68 2433 102
rect 2367 48 2433 68
rect 31 17 2561 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 127 564 161 598
rect 655 564 689 598
rect 1135 532 1169 566
rect 1231 564 1265 598
rect 367 451 401 485
rect 943 451 977 485
rect 1711 532 1745 566
rect 1807 564 1841 598
rect 2383 564 2417 598
rect 1519 451 1553 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1423 368 1457 402
rect 1999 368 2033 402
rect 559 262 593 296
rect 1135 289 1169 323
rect 1711 289 1745 323
rect 271 181 305 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 1423 181 1457 215
rect 1711 181 1745 215
rect 1999 181 2033 215
rect 2287 368 2321 402
rect 2287 181 2321 215
rect 127 68 161 102
rect 367 100 401 134
rect 655 68 689 102
rect 943 100 977 134
rect 1231 68 1265 102
rect 1519 100 1553 134
rect 1807 68 1841 102
rect 2095 100 2129 134
rect 2383 68 2417 102
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 714
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 618 2592 649
rect 115 598 173 618
rect 115 564 127 598
rect 161 564 173 598
rect 115 552 173 564
rect 643 598 701 618
rect 643 564 655 598
rect 689 564 701 598
rect 1219 598 1277 618
rect 274 535 590 563
rect 643 552 701 564
rect 1123 566 1181 578
rect 1123 563 1135 566
rect 274 414 302 535
rect 355 485 413 497
rect 355 451 367 485
rect 401 451 413 485
rect 355 439 413 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 274 227 302 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 370 212 398 439
rect 562 414 590 535
rect 850 535 1135 563
rect 850 414 878 535
rect 1123 532 1135 535
rect 1169 532 1181 566
rect 1219 564 1231 598
rect 1265 564 1277 598
rect 1795 598 1853 618
rect 1219 552 1277 564
rect 1699 566 1757 578
rect 1699 563 1711 566
rect 1123 520 1181 532
rect 1426 535 1711 563
rect 931 485 989 497
rect 931 451 943 485
rect 977 451 989 485
rect 931 439 989 451
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 946 399 974 439
rect 1426 414 1454 535
rect 1699 532 1711 535
rect 1745 532 1757 566
rect 1795 564 1807 598
rect 1841 564 1853 598
rect 1795 552 1853 564
rect 2371 598 2429 618
rect 2371 564 2383 598
rect 2417 564 2429 598
rect 2371 552 2429 564
rect 1699 520 1757 532
rect 1507 485 1565 497
rect 1507 451 1519 485
rect 1553 451 1565 485
rect 1507 439 1565 451
rect 1411 402 1469 414
rect 1411 399 1423 402
rect 946 371 1423 399
rect 562 308 590 356
rect 547 296 605 308
rect 547 262 559 296
rect 593 262 605 296
rect 547 250 605 262
rect 850 227 878 356
rect 835 215 893 227
rect 835 212 847 215
rect 370 184 847 212
rect 370 146 398 184
rect 835 181 847 184
rect 881 181 893 215
rect 835 169 893 181
rect 946 146 974 371
rect 1411 368 1423 371
rect 1457 368 1469 402
rect 1411 356 1469 368
rect 1522 399 1550 439
rect 1987 402 2045 414
rect 1987 399 1999 402
rect 1522 371 1999 399
rect 1123 323 1181 335
rect 1123 289 1135 323
rect 1169 289 1181 323
rect 1123 277 1181 289
rect 1138 227 1166 277
rect 1426 227 1454 356
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 1411 215 1469 227
rect 1411 181 1423 215
rect 1457 181 1469 215
rect 1411 169 1469 181
rect 1522 146 1550 371
rect 1987 368 1999 371
rect 2033 399 2045 402
rect 2275 402 2333 414
rect 2275 399 2287 402
rect 2033 371 2287 399
rect 2033 368 2045 371
rect 1987 356 2045 368
rect 2275 368 2287 371
rect 2321 368 2333 402
rect 2275 356 2333 368
rect 1699 323 1757 335
rect 1699 289 1711 323
rect 1745 289 1757 323
rect 1699 277 1757 289
rect 1714 227 1742 277
rect 2002 227 2030 356
rect 2290 227 2318 356
rect 1699 215 1757 227
rect 1699 181 1711 215
rect 1745 181 1757 215
rect 1699 169 1757 181
rect 1987 215 2045 227
rect 1987 181 1999 215
rect 2033 181 2045 215
rect 1987 169 2045 181
rect 2275 215 2333 227
rect 2275 181 2287 215
rect 2321 181 2333 215
rect 2275 169 2333 181
rect 355 134 413 146
rect 115 102 173 114
rect 115 68 127 102
rect 161 68 173 102
rect 355 100 367 134
rect 401 100 413 134
rect 931 134 989 146
rect 355 88 413 100
rect 643 102 701 114
rect 115 48 173 68
rect 643 68 655 102
rect 689 68 701 102
rect 931 100 943 134
rect 977 100 989 134
rect 1507 134 1565 146
rect 931 88 989 100
rect 1219 102 1277 114
rect 643 48 701 68
rect 1219 68 1231 102
rect 1265 68 1277 102
rect 1507 100 1519 134
rect 1553 100 1565 134
rect 2083 134 2141 146
rect 1507 88 1565 100
rect 1795 102 1853 114
rect 1219 48 1277 68
rect 1795 68 1807 102
rect 1841 68 1853 102
rect 2083 100 2095 134
rect 2129 100 2141 134
rect 2083 88 2141 100
rect 2371 102 2429 114
rect 1795 48 1853 68
rect 2371 68 2383 102
rect 2417 68 2429 102
rect 2371 48 2429 68
rect 0 17 2592 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -48 2592 -17
<< labels >>
rlabel metal1 0 618 2592 714 0 VPWR
port 2 se
rlabel metal1 0 618 2592 714 0 VPWR
port 2 se
rlabel metal1 0 -48 2592 48 0 VGND
port 1 se
rlabel metal1 0 -48 2592 48 0 VGND
port 1 se
rlabel metal1 2083 88 2141 146 0 Y
port 3 se
rlabel metal1 259 169 317 227 0 A
port 0 se
rlabel metal1 547 250 605 308 0 A
port 0 se
rlabel metal1 274 227 302 356 0 A
port 0 se
rlabel metal1 562 308 590 356 0 A
port 0 se
rlabel metal1 259 356 317 414 0 A
port 0 se
rlabel metal1 547 356 605 414 0 A
port 0 se
rlabel metal1 274 414 302 535 0 A
port 0 se
rlabel metal1 562 414 590 535 0 A
port 0 se
rlabel metal1 274 535 590 563 0 A
port 0 se
rlabel locali 0 -17 2592 17 4 VGND
port 1 se ground default abutment
rlabel locali 31 17 2561 48 4 VGND
port 1 se ground default abutment
rlabel locali 0 649 2592 683 4 VPWR
port 2 se power default abutment
rlabel locali 31 618 2561 649 4 VGND
port 1 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 2592 666
<< end >>
