VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.385 1.585 1.675 ;
        RECT 1.370 1.135 1.510 1.385 ;
        RECT 1.295 0.845 1.585 1.135 ;
    END
  END A
  PIN VGND
    ANTENNADIFFAREA 0.562100 ;
    PORT
      LAYER met1 ;
        RECT 1.775 0.440 2.065 0.730 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 0.000 -0.240 4.320 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 4.320 3.570 ;
        RECT 1.775 2.735 2.065 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 4.320 3.415 ;
        RECT 0.155 3.090 4.165 3.245 ;
        RECT 1.755 2.715 2.085 3.090 ;
      LAYER mcon ;
        RECT 1.835 3.245 2.005 3.415 ;
        RECT 1.835 2.795 2.005 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.031650 ;
    PORT
      LAYER met1 ;
        RECT 3.215 2.195 3.505 2.485 ;
        RECT 3.290 0.730 3.430 2.195 ;
        RECT 3.215 0.440 3.505 0.730 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 4.320 3.330 ;
      LAYER li1 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 3.195 2.260 3.525 2.505 ;
        RECT 3.215 2.175 3.525 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 1.355 1.445 1.525 1.760 ;
        RECT 1.275 0.920 1.605 1.155 ;
        RECT 2.715 0.920 3.045 1.155 ;
        RECT 1.275 0.825 1.585 0.920 ;
        RECT 2.715 0.825 3.025 0.920 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.755 0.420 2.085 0.750 ;
        RECT 3.195 0.420 3.525 0.750 ;
        RECT 0.155 0.085 4.165 0.240 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 3.275 2.255 3.445 2.425 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 1.835 0.500 2.005 0.670 ;
        RECT 3.275 0.500 3.445 0.670 ;
        RECT 1.835 -0.085 2.005 0.085 ;
      LAYER met1 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 0.650 1.995 0.790 2.195 ;
        RECT 2.735 1.995 3.025 2.070 ;
        RECT 0.650 1.855 3.025 1.995 ;
        RECT 0.650 0.730 0.790 1.855 ;
        RECT 2.735 1.780 3.025 1.855 ;
        RECT 2.810 1.135 2.950 1.780 ;
        RECT 2.735 0.845 3.025 1.135 ;
        RECT 0.575 0.440 0.865 0.730 ;
  END
END BUFX2
END LIBRARY

