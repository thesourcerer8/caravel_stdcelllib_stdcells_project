MACRO LATCH
 CLASS CORE ;
 FOREIGN LATCH 0 0 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE CORE ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.09000000 10.08000000 3.57000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 10.08000000 0.24000000 ;
    END
  END GND

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 8.97500000 0.39500000 9.26500000 0.68500000 ;
        RECT 7.05500000 1.74500000 7.34500000 2.03500000 ;
        RECT 9.05000000 0.68500000 9.19000000 2.15000000 ;
        RECT 7.13000000 2.03500000 7.27000000 2.22500000 ;
        RECT 8.97500000 2.15000000 9.26500000 2.22500000 ;
        RECT 7.13000000 2.22500000 9.26500000 2.36500000 ;
        RECT 8.97500000 2.36500000 9.26500000 2.44000000 ;
    END
  END Q

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.73500000 1.20500000 3.02500000 1.49500000 ;
    END
  END D

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.29500000 0.80000000 1.58500000 0.87500000 ;
        RECT 4.17500000 0.80000000 4.46500000 0.87500000 ;
        RECT 1.29500000 0.87500000 4.46500000 1.01500000 ;
        RECT 1.29500000 1.01500000 1.58500000 1.09000000 ;
        RECT 4.17500000 1.01500000 4.46500000 1.09000000 ;
    END
  END CLK


END LATCH
