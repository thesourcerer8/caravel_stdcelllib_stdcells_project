magic
tech sky130A
timestamp 1621277951
<< end >>
