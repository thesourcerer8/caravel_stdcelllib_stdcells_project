magic
tech sky130A
timestamp 1623602962
<< nwell >>
rect 0 179 432 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
<< ndiff >>
rect 58 66 87 69
rect 322 66 351 69
rect 58 63 137 66
rect 58 46 64 63
rect 81 46 137 63
rect 58 24 137 46
rect 152 36 281 66
rect 152 24 184 36
rect 178 19 184 24
rect 201 24 281 36
rect 296 63 375 66
rect 296 46 328 63
rect 345 46 375 63
rect 296 24 375 46
rect 201 19 207 24
rect 178 13 207 19
<< pdiff >>
rect 178 309 207 312
rect 58 238 137 309
rect 58 221 64 238
rect 81 225 137 238
rect 152 306 281 309
rect 152 289 184 306
rect 201 289 281 306
rect 152 225 281 289
rect 296 238 375 309
rect 296 225 328 238
rect 81 221 87 225
rect 58 215 87 221
rect 322 221 328 225
rect 345 225 375 238
rect 345 221 351 225
rect 322 215 351 221
<< ndiffc >>
rect 64 46 81 63
rect 184 19 201 36
rect 328 46 345 63
<< pdiffc >>
rect 64 221 81 238
rect 184 289 201 306
rect 328 221 345 238
<< poly >>
rect 137 309 152 330
rect 281 309 296 330
rect 137 206 152 225
rect 281 206 296 225
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 305 206
rect 272 181 280 198
rect 297 181 305 198
rect 272 173 305 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 86 305 103
rect 272 78 305 86
rect 137 66 152 78
rect 281 66 296 78
rect 137 11 152 24
rect 281 11 296 24
<< polycont >>
rect 136 181 153 198
rect 280 181 297 198
rect 136 86 153 103
rect 280 86 297 103
<< locali >>
rect 176 306 209 314
rect 176 289 184 306
rect 201 289 209 306
rect 176 281 209 289
rect 56 238 89 246
rect 56 221 64 238
rect 81 221 89 238
rect 56 213 89 221
rect 320 238 353 246
rect 320 221 328 238
rect 345 221 353 238
rect 320 213 353 221
rect 128 198 161 206
rect 128 181 136 198
rect 153 181 161 198
rect 128 173 161 181
rect 272 198 303 206
rect 272 181 280 198
rect 297 196 303 198
rect 297 181 305 196
rect 272 173 305 181
rect 128 103 161 111
rect 128 86 136 103
rect 153 86 161 103
rect 128 78 161 86
rect 272 103 305 111
rect 272 86 280 103
rect 297 88 305 103
rect 297 86 303 88
rect 272 78 303 86
rect 56 63 89 71
rect 56 46 64 63
rect 81 46 89 63
rect 56 38 89 46
rect 320 63 353 71
rect 320 46 328 63
rect 345 46 353 63
rect 176 36 209 44
rect 320 38 353 46
rect 176 19 184 36
rect 201 19 209 36
rect 176 11 209 19
<< viali >>
rect 184 289 201 306
rect 64 221 81 238
rect 328 221 345 238
rect 136 181 153 198
rect 280 181 297 198
rect 136 86 153 103
rect 280 86 297 103
rect 64 46 81 63
rect 328 46 345 63
rect 184 19 201 36
<< metal1 >>
rect 0 309 432 357
rect 178 306 207 309
rect 178 289 184 306
rect 201 289 207 306
rect 178 283 207 289
rect 58 238 87 244
rect 58 221 64 238
rect 81 237 87 238
rect 322 238 351 244
rect 322 237 328 238
rect 81 223 328 237
rect 81 221 87 223
rect 58 215 87 221
rect 322 221 328 223
rect 345 221 351 238
rect 322 215 351 221
rect 65 69 79 215
rect 130 198 159 204
rect 130 181 136 198
rect 153 181 159 198
rect 130 175 159 181
rect 274 198 303 204
rect 274 181 280 198
rect 297 181 303 198
rect 274 175 303 181
rect 137 109 151 175
rect 281 109 295 175
rect 130 103 159 109
rect 130 86 136 103
rect 153 102 159 103
rect 274 103 303 109
rect 274 102 280 103
rect 153 88 280 102
rect 153 86 159 88
rect 130 80 159 86
rect 274 86 280 88
rect 297 86 303 103
rect 274 80 303 86
rect 329 69 343 215
rect 58 63 87 69
rect 58 46 64 63
rect 81 46 87 63
rect 58 40 87 46
rect 322 63 351 69
rect 322 46 328 63
rect 345 46 351 63
rect 178 36 207 42
rect 322 40 351 46
rect 178 24 184 36
rect 0 19 184 24
rect 201 24 207 36
rect 201 19 432 24
rect 0 -24 432 19
<< labels >>
rlabel metal1 0 309 432 357 0 VDD
port 1 se
rlabel metal1 0 -24 432 24 0 GND
port 2 se
rlabel metal1 58 40 87 69 0 Y
port 3 se
rlabel metal1 322 40 351 69 0 Y
port 4 se
rlabel metal1 65 69 79 215 0 Y
port 5 se
rlabel metal1 329 69 343 215 0 Y
port 6 se
rlabel metal1 58 215 87 223 0 Y
port 7 se
rlabel metal1 322 215 351 223 0 Y
port 8 se
rlabel metal1 58 223 351 237 0 Y
port 9 se
rlabel metal1 58 237 87 244 0 Y
port 10 se
rlabel metal1 322 237 351 244 0 Y
port 11 se
rlabel metal1 130 80 159 88 0 A
port 12 se
rlabel metal1 274 80 303 88 0 A
port 13 se
rlabel metal1 130 88 303 102 0 A
port 14 se
rlabel metal1 130 102 159 109 0 A
port 15 se
rlabel metal1 274 102 303 109 0 A
port 16 se
rlabel metal1 137 109 151 175 0 A
port 17 se
rlabel metal1 281 109 295 175 0 A
port 18 se
rlabel metal1 130 175 159 204 0 A
port 19 se
rlabel metal1 274 175 303 204 0 A
port 20 se
<< properties >>
string FIXED_BBOX 0 0 432 333
<< end >>
