VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 2.880 3.570 ;
        RECT 1.780 2.970 2.070 3.090 ;
        RECT 1.780 2.800 1.840 2.970 ;
        RECT 2.010 2.800 2.070 2.970 ;
        RECT 1.780 2.740 2.070 2.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.090 2.880 3.570 ;
        RECT 1.760 2.970 2.090 3.090 ;
        RECT 1.760 2.800 1.840 2.970 ;
        RECT 2.010 2.800 2.090 2.970 ;
        RECT 1.760 2.720 2.090 2.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.670 2.070 0.730 ;
        RECT 1.780 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.070 0.670 ;
        RECT 1.780 0.440 2.070 0.500 ;
        RECT 1.850 0.240 1.990 0.440 ;
        RECT 0.000 -0.240 2.880 0.240 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.240 2.880 0.240 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.580 2.200 0.870 2.490 ;
        RECT 0.650 0.730 0.790 2.200 ;
        RECT 0.580 0.440 0.870 0.730 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.300 1.780 1.590 2.070 ;
        RECT 1.370 1.140 1.510 1.780 ;
        RECT 1.300 0.850 1.590 1.140 ;
    END
  END A
  OBS
      LAYER li1 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.920 1.610 1.080 ;
        RECT 1.530 0.910 1.590 0.920 ;
        RECT 1.280 0.830 1.590 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 1.760 0.670 2.090 0.750 ;
        RECT 1.760 0.500 1.840 0.670 ;
        RECT 2.010 0.500 2.090 0.670 ;
        RECT 1.760 0.420 2.090 0.500 ;
  END
END INVX2
END LIBRARY

