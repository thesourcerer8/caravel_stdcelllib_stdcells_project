magic
tech sky130A
magscale 1 2
timestamp 1636809598
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1440 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
<< ndiff >>
rect 163 134 221 146
rect 163 132 175 134
rect 115 100 175 132
rect 209 132 221 134
rect 355 134 413 146
rect 355 132 367 134
rect 209 100 273 132
rect 115 48 273 100
rect 303 100 367 132
rect 401 132 413 134
rect 739 134 797 146
rect 739 132 751 134
rect 401 100 561 132
rect 303 48 561 100
rect 591 100 751 132
rect 785 132 797 134
rect 1027 134 1085 146
rect 1027 132 1039 134
rect 785 100 849 132
rect 591 48 849 100
rect 879 100 1039 132
rect 1073 132 1085 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 1073 100 1137 132
rect 879 48 1137 100
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1265 100 1325 132
rect 1167 48 1325 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 175 485
rect 209 451 273 485
rect 115 450 273 451
rect 303 450 561 618
rect 591 593 849 618
rect 591 559 655 593
rect 689 559 849 593
rect 591 450 849 559
rect 879 450 1137 618
rect 1167 485 1325 618
rect 1167 451 1231 485
rect 1265 451 1325 485
rect 1167 450 1325 451
rect 163 439 221 450
rect 1219 439 1277 450
<< ndiffc >>
rect 175 100 209 134
rect 367 100 401 134
rect 751 100 785 134
rect 1039 100 1073 134
rect 1231 100 1265 134
<< pdiffc >>
rect 175 451 209 485
rect 655 559 689 593
rect 1231 451 1265 485
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
<< locali >>
rect 0 649 655 683
rect 689 649 1440 683
rect 31 618 1409 649
rect 639 593 705 618
rect 639 559 655 593
rect 689 559 705 593
rect 639 543 705 559
rect 159 485 225 501
rect 159 451 175 485
rect 209 452 225 485
rect 1215 485 1281 501
rect 209 451 221 452
rect 159 435 221 451
rect 1215 451 1231 485
rect 1265 451 1281 485
rect 1215 435 1281 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1181 418
rect 1119 368 1135 402
rect 1169 401 1181 402
rect 1169 368 1185 401
rect 1119 352 1185 368
rect 255 215 321 231
rect 255 184 271 215
rect 259 181 271 184
rect 305 181 321 215
rect 259 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 831 215 897 231
rect 1119 215 1185 231
rect 831 184 847 215
rect 543 165 609 181
rect 835 181 847 184
rect 881 181 897 215
rect 835 165 897 181
rect 1039 150 1073 181
rect 1119 181 1135 215
rect 1169 184 1185 215
rect 1169 181 1181 184
rect 1119 165 1181 181
rect 159 134 225 150
rect 159 100 175 134
rect 209 100 225 134
rect 355 134 417 150
rect 355 131 367 134
rect 159 84 225 100
rect 351 100 367 131
rect 401 100 417 134
rect 351 84 417 100
rect 735 134 801 150
rect 735 100 751 134
rect 785 100 801 134
rect 735 84 801 100
rect 1023 134 1085 150
rect 1023 100 1039 134
rect 1073 131 1085 134
rect 1215 134 1281 150
rect 1073 100 1089 131
rect 1023 84 1089 100
rect 1215 100 1231 134
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 367 48 401 84
rect 31 17 1409 48
rect 0 -17 367 17
rect 401 -17 1440 17
<< viali >>
rect 655 649 689 683
rect 655 559 689 593
rect 175 451 209 485
rect 1231 451 1265 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1039 181 1073 215
rect 1135 181 1169 215
rect 175 100 209 134
rect 751 100 785 134
rect 1231 100 1265 134
rect 367 -17 401 17
<< metal1 >>
rect 0 683 1440 714
rect 0 649 655 683
rect 689 649 1440 683
rect 0 618 1440 649
rect 643 593 701 618
rect 643 559 655 593
rect 689 559 701 593
rect 643 547 701 559
rect 163 485 221 497
rect 163 451 175 485
rect 209 482 221 485
rect 1219 485 1277 497
rect 1219 482 1231 485
rect 209 454 1231 482
rect 209 451 221 454
rect 163 439 221 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 274 227 302 356
rect 562 227 590 356
rect 850 227 878 356
rect 1042 227 1070 454
rect 1219 451 1231 454
rect 1265 451 1277 485
rect 1219 439 1277 451
rect 1123 402 1181 414
rect 1123 368 1135 402
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 1138 227 1166 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 835 215 893 227
rect 835 181 847 215
rect 881 181 893 215
rect 835 169 893 181
rect 1027 215 1085 227
rect 1027 181 1039 215
rect 1073 181 1085 215
rect 1027 169 1085 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 163 134 221 146
rect 163 100 175 134
rect 209 131 221 134
rect 739 134 797 146
rect 739 131 751 134
rect 209 103 751 131
rect 209 100 221 103
rect 163 88 221 100
rect 739 100 751 103
rect 785 131 797 134
rect 1219 134 1277 146
rect 1219 131 1231 134
rect 785 103 1231 131
rect 785 100 797 103
rect 739 88 797 100
rect 1219 100 1231 103
rect 1265 100 1277 134
rect 1219 88 1277 100
rect 0 17 1440 48
rect 0 -17 367 17
rect 401 -17 1440 17
rect 0 -48 1440 -17
<< labels >>
rlabel metal1 0 618 1440 714 0 VPWR
port 5 se
rlabel metal1 0 618 1440 714 0 VPWR
port 5 se
rlabel metal1 0 -48 1440 48 0 VGND
port 4 se
rlabel metal1 0 -48 1440 48 0 VGND
port 4 se
rlabel metal1 1027 169 1085 227 0 Y
port 6 se
rlabel metal1 163 439 221 454 0 Y
port 6 se
rlabel metal1 1042 227 1070 454 0 Y
port 6 se
rlabel metal1 1219 439 1277 454 0 Y
port 6 se
rlabel metal1 163 454 1277 482 0 Y
port 6 se
rlabel metal1 163 482 221 497 0 Y
port 6 se
rlabel metal1 1219 482 1277 497 0 Y
port 6 se
rlabel metal1 835 169 893 227 0 C
port 2 se
rlabel metal1 850 227 878 356 0 C
port 2 se
rlabel metal1 835 356 893 414 0 C
port 2 se
rlabel metal1 259 169 317 227 0 B
port 1 se
rlabel metal1 274 227 302 356 0 B
port 1 se
rlabel metal1 259 356 317 414 0 B
port 1 se
rlabel metal1 1123 169 1181 227 0 D
port 3 se
rlabel metal1 1138 227 1166 356 0 D
port 3 se
rlabel metal1 1123 356 1181 414 0 D
port 3 se
rlabel metal1 547 169 605 227 0 A
port 0 se
rlabel metal1 562 227 590 356 0 A
port 0 se
rlabel metal1 547 356 605 414 0 A
port 0 se
rlabel locali 0 -17 1440 17 4 VGND
port 4 se ground default abutment
rlabel locali 31 17 1409 48 4 VGND
port 4 se ground default abutment
rlabel locali 0 649 1440 683 4 VPWR
port 5 se power default abutment
rlabel locali 31 618 1409 649 4 VGND
port 4 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1440 666
<< end >>
