magic
tech sky130A
timestamp 1624066365
<< nwell >>
rect 0 179 864 333
<< nmos >>
rect 137 24 152 66
rect 281 24 296 66
rect 425 24 440 66
rect 569 24 584 66
rect 713 24 728 66
<< pmos >>
rect 137 225 152 309
rect 281 225 296 309
rect 425 225 440 309
rect 569 225 584 309
rect 713 225 728 309
<< ndiff >>
rect 58 67 87 73
rect 58 50 64 67
rect 81 66 87 67
rect 514 67 543 73
rect 514 66 520 67
rect 81 50 137 66
rect 58 24 137 50
rect 152 49 281 66
rect 152 32 184 49
rect 201 32 281 49
rect 152 24 281 32
rect 296 24 425 66
rect 440 50 520 66
rect 537 66 543 67
rect 537 50 569 66
rect 440 24 569 50
rect 584 24 713 66
rect 728 49 807 66
rect 728 32 760 49
rect 777 32 807 49
rect 728 24 807 32
<< pdiff >>
rect 58 243 137 309
rect 58 226 64 243
rect 81 226 137 243
rect 58 225 137 226
rect 152 301 281 309
rect 152 284 184 301
rect 201 284 281 301
rect 152 225 281 284
rect 296 225 425 309
rect 440 243 569 309
rect 440 226 520 243
rect 537 226 569 243
rect 440 225 569 226
rect 584 225 713 309
rect 728 301 807 309
rect 728 284 760 301
rect 777 284 807 301
rect 728 225 807 284
rect 58 220 87 225
rect 514 220 543 225
<< ndiffc >>
rect 64 50 81 67
rect 184 32 201 49
rect 520 50 537 67
rect 760 32 777 49
<< pdiffc >>
rect 64 226 81 243
rect 184 284 201 301
rect 520 226 537 243
rect 760 284 777 301
<< poly >>
rect 137 309 152 322
rect 281 309 296 322
rect 425 309 440 322
rect 569 309 584 322
rect 713 309 728 322
rect 137 209 152 225
rect 281 209 296 225
rect 425 209 440 225
rect 569 209 584 225
rect 713 209 728 225
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 201 593 209
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 560 108 593 116
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 137 66 152 83
rect 281 66 296 83
rect 425 66 440 83
rect 569 66 584 83
rect 713 66 728 83
rect 137 11 152 24
rect 281 11 296 24
rect 425 11 440 24
rect 569 11 584 24
rect 713 11 728 24
<< polycont >>
rect 136 184 153 201
rect 280 184 297 201
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 136 91 153 108
rect 280 91 297 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
<< locali >>
rect 176 301 209 309
rect 176 284 184 301
rect 201 284 209 301
rect 176 276 209 284
rect 752 301 785 309
rect 752 284 760 301
rect 777 284 785 301
rect 752 276 785 284
rect 56 243 89 251
rect 56 226 64 243
rect 81 226 89 243
rect 56 218 89 226
rect 512 243 545 251
rect 512 226 520 243
rect 537 226 545 243
rect 512 218 545 226
rect 128 201 161 209
rect 128 184 136 201
rect 153 184 161 201
rect 128 176 161 184
rect 272 201 305 209
rect 272 184 280 201
rect 297 184 305 201
rect 272 176 305 184
rect 416 201 449 209
rect 562 201 593 209
rect 416 184 424 201
rect 441 184 449 201
rect 416 176 449 184
rect 560 184 568 201
rect 585 184 593 201
rect 560 176 593 184
rect 704 201 737 209
rect 704 184 712 201
rect 729 184 737 201
rect 704 176 737 184
rect 136 116 153 176
rect 280 148 297 176
rect 280 116 297 131
rect 128 108 161 116
rect 128 91 136 108
rect 153 91 161 108
rect 128 83 161 91
rect 272 108 305 116
rect 272 91 280 108
rect 297 91 305 108
rect 272 83 305 91
rect 416 108 449 116
rect 416 91 424 108
rect 441 91 449 108
rect 416 83 449 91
rect 520 75 537 131
rect 560 108 593 116
rect 560 92 568 108
rect 562 91 568 92
rect 585 91 593 108
rect 562 83 593 91
rect 704 108 737 116
rect 704 91 712 108
rect 729 91 737 108
rect 704 83 737 91
rect 56 67 89 75
rect 56 50 64 67
rect 81 50 89 67
rect 512 67 545 75
rect 56 42 89 50
rect 176 49 209 57
rect 176 32 184 49
rect 201 32 209 49
rect 512 50 520 67
rect 537 50 545 67
rect 512 42 545 50
rect 752 49 785 57
rect 176 24 209 32
rect 752 32 760 49
rect 777 32 785 49
rect 752 24 785 32
<< viali >>
rect 184 284 201 301
rect 760 284 777 301
rect 64 226 81 243
rect 520 226 537 243
rect 424 184 441 201
rect 568 184 585 201
rect 712 184 729 201
rect 280 131 297 148
rect 520 131 537 148
rect 136 91 153 108
rect 424 91 441 108
rect 568 91 585 108
rect 712 91 729 108
rect 64 50 81 67
rect 184 32 201 49
rect 760 32 777 49
<< metal1 >>
rect 0 309 864 357
rect 178 301 207 309
rect 178 284 184 301
rect 201 284 207 301
rect 178 278 207 284
rect 754 301 783 309
rect 754 284 760 301
rect 777 284 783 301
rect 754 278 783 284
rect 58 243 87 249
rect 58 226 64 243
rect 81 226 87 243
rect 58 220 87 226
rect 514 243 543 249
rect 514 226 520 243
rect 537 226 543 243
rect 514 220 543 226
rect 65 200 79 220
rect 418 201 447 207
rect 418 200 424 201
rect 65 186 424 200
rect 65 73 79 186
rect 418 184 424 186
rect 441 200 447 201
rect 441 186 487 200
rect 441 184 447 186
rect 418 178 447 184
rect 274 148 303 154
rect 274 131 280 148
rect 297 131 303 148
rect 274 125 303 131
rect 130 108 159 114
rect 130 91 136 108
rect 153 106 159 108
rect 418 108 447 114
rect 418 106 424 108
rect 153 92 424 106
rect 153 91 159 92
rect 130 85 159 91
rect 418 91 424 92
rect 441 91 447 108
rect 473 106 487 186
rect 521 154 535 220
rect 562 201 591 207
rect 562 184 568 201
rect 585 200 591 201
rect 706 201 735 207
rect 585 186 631 200
rect 585 184 591 186
rect 562 178 591 184
rect 514 148 543 154
rect 514 131 520 148
rect 537 131 543 148
rect 514 125 543 131
rect 562 108 591 114
rect 562 106 568 108
rect 473 92 568 106
rect 418 85 447 91
rect 562 91 568 92
rect 585 91 591 108
rect 562 85 591 91
rect 58 67 87 73
rect 58 50 64 67
rect 81 50 87 67
rect 425 66 439 85
rect 617 66 631 186
rect 706 184 712 201
rect 729 184 735 201
rect 706 178 735 184
rect 713 114 727 178
rect 706 108 735 114
rect 706 91 712 108
rect 729 91 735 108
rect 706 85 735 91
rect 58 44 87 50
rect 178 49 207 55
rect 425 52 631 66
rect 178 32 184 49
rect 201 32 207 49
rect 178 24 207 32
rect 754 49 783 55
rect 754 32 760 49
rect 777 32 783 49
rect 754 24 783 32
rect 0 -24 864 24
<< labels >>
rlabel metal1 0 309 864 357 0 VDD
port 1 se
rlabel metal1 0 -24 864 24 0 GND
port 2 se
rlabel metal1 514 125 543 154 0 Y
port 3 se
rlabel metal1 521 154 535 220 0 Y
port 4 se
rlabel metal1 514 220 543 249 0 Y
port 5 se
rlabel metal1 425 52 631 66 0 S
port 6 se
rlabel metal1 425 66 439 85 0 S
port 7 se
rlabel metal1 130 85 159 92 0 S
port 8 se
rlabel metal1 418 85 447 92 0 S
port 9 se
rlabel metal1 130 92 447 106 0 S
port 10 se
rlabel metal1 130 106 159 114 0 S
port 11 se
rlabel metal1 418 106 447 114 0 S
port 12 se
rlabel metal1 562 178 591 186 0 S
port 13 se
rlabel metal1 617 66 631 186 0 S
port 14 se
rlabel metal1 562 186 631 200 0 S
port 15 se
rlabel metal1 562 200 591 207 0 S
port 16 se
rlabel metal1 274 125 303 154 0 A
port 17 se
rlabel metal1 706 85 735 114 0 B
port 18 se
rlabel metal1 713 114 727 178 0 B
port 19 se
rlabel metal1 706 178 735 207 0 B
port 20 se
<< properties >>
string FIXED_BBOX 0 0 864 333
<< end >>
