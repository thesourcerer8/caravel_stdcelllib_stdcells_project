magic
tech sky130A
magscale 1 2
timestamp 1636962369
<< checkpaint >>
rect -1260 -1374 11260 2038
<< nwell >>
rect 0 358 1440 666
<< nmos >>
rect 273 48 303 132
rect 561 48 591 132
rect 849 48 879 132
rect 1137 48 1167 132
<< pmos >>
rect 273 450 303 618
rect 561 450 591 618
rect 849 450 879 618
rect 1137 450 1167 618
<< ndiff >>
rect 163 134 221 146
rect 163 132 175 134
rect 115 100 175 132
rect 209 132 221 134
rect 643 134 701 146
rect 643 132 655 134
rect 209 100 273 132
rect 115 48 273 100
rect 303 48 561 132
rect 591 100 655 132
rect 689 132 701 134
rect 1219 134 1277 146
rect 1219 132 1231 134
rect 689 100 849 132
rect 591 48 849 100
rect 879 48 1137 132
rect 1167 100 1231 132
rect 1265 132 1277 134
rect 1265 100 1325 132
rect 1167 48 1325 100
<< pdiff >>
rect 115 485 273 618
rect 115 451 175 485
rect 209 451 273 485
rect 115 450 273 451
rect 303 593 561 618
rect 303 559 367 593
rect 401 559 561 593
rect 303 450 561 559
rect 591 485 849 618
rect 591 451 655 485
rect 689 451 849 485
rect 591 450 849 451
rect 879 485 1137 618
rect 879 451 1039 485
rect 1073 451 1137 485
rect 879 450 1137 451
rect 1167 566 1325 618
rect 1167 532 1231 566
rect 1265 532 1325 566
rect 1167 450 1325 532
rect 163 439 221 450
rect 643 439 701 450
rect 1027 439 1085 450
<< ndiffc >>
rect 175 100 209 134
rect 655 100 689 134
rect 1231 100 1265 134
<< pdiffc >>
rect 175 451 209 485
rect 367 559 401 593
rect 655 451 689 485
rect 1039 451 1073 485
rect 1231 532 1265 566
<< poly >>
rect 273 618 303 644
rect 561 618 591 644
rect 849 618 879 644
rect 1137 618 1167 644
rect 273 418 303 450
rect 561 418 591 450
rect 849 418 879 450
rect 1137 418 1167 450
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 255 215 321 231
rect 255 181 271 215
rect 305 181 321 215
rect 255 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 181 1185 215
rect 1119 165 1185 181
rect 273 132 303 165
rect 561 132 591 165
rect 849 132 879 165
rect 1137 132 1167 165
rect 273 22 303 48
rect 561 22 591 48
rect 849 22 879 48
rect 1137 22 1167 48
<< polycont >>
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
<< locali >>
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1440 683
rect 31 618 1409 649
rect 351 593 417 618
rect 351 559 367 593
rect 401 559 417 593
rect 351 543 417 559
rect 1215 566 1281 582
rect 1215 532 1231 566
rect 1265 532 1281 566
rect 1215 516 1281 532
rect 159 485 225 501
rect 159 451 175 485
rect 209 452 225 485
rect 639 485 705 501
rect 639 452 655 485
rect 209 451 221 452
rect 159 435 221 451
rect 643 451 655 452
rect 689 451 705 485
rect 643 435 705 451
rect 1023 485 1089 501
rect 1023 451 1039 485
rect 1073 452 1089 485
rect 1073 451 1085 452
rect 1023 435 1085 451
rect 255 402 321 418
rect 255 368 271 402
rect 305 368 321 402
rect 255 352 321 368
rect 543 402 609 418
rect 543 368 559 402
rect 593 368 609 402
rect 543 352 609 368
rect 831 402 897 418
rect 831 368 847 402
rect 881 368 897 402
rect 831 352 897 368
rect 1119 402 1185 418
rect 1119 368 1135 402
rect 1169 368 1185 402
rect 1119 352 1185 368
rect 255 215 321 231
rect 255 184 271 215
rect 259 181 271 184
rect 305 181 321 215
rect 259 165 321 181
rect 543 215 609 231
rect 543 181 559 215
rect 593 181 609 215
rect 543 165 609 181
rect 831 215 897 231
rect 831 181 847 215
rect 881 181 897 215
rect 831 165 897 181
rect 1119 215 1185 231
rect 1119 181 1135 215
rect 1169 184 1185 215
rect 1169 181 1181 184
rect 1119 165 1181 181
rect 159 134 225 150
rect 159 100 175 134
rect 209 100 225 134
rect 643 134 705 150
rect 643 131 655 134
rect 159 84 225 100
rect 639 100 655 131
rect 689 100 705 134
rect 639 84 705 100
rect 1215 134 1281 150
rect 1215 100 1231 134
rect 1265 100 1281 134
rect 1215 84 1281 100
rect 655 48 689 84
rect 31 17 1409 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1440 17
<< viali >>
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 367 559 401 593
rect 1231 532 1265 566
rect 175 451 209 485
rect 655 451 689 485
rect 1039 451 1073 485
rect 271 368 305 402
rect 559 368 593 402
rect 847 368 881 402
rect 1135 368 1169 402
rect 271 181 305 215
rect 559 181 593 215
rect 847 181 881 215
rect 1135 181 1169 215
rect 175 100 209 134
rect 1231 100 1265 134
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1440 714
rect 0 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1440 683
rect 0 618 1440 649
rect 355 593 413 618
rect 355 559 367 593
rect 401 559 413 593
rect 1219 566 1277 578
rect 1219 563 1231 566
rect 355 547 413 559
rect 658 535 1231 563
rect 658 497 686 535
rect 1219 532 1231 535
rect 1265 532 1277 566
rect 1219 520 1277 532
rect 163 485 221 497
rect 163 451 175 485
rect 209 482 221 485
rect 643 485 701 497
rect 643 482 655 485
rect 209 454 655 482
rect 209 451 221 454
rect 163 439 221 451
rect 643 451 655 454
rect 689 451 701 485
rect 643 439 701 451
rect 1027 485 1085 497
rect 1027 451 1039 485
rect 1073 482 1085 485
rect 1073 454 1262 482
rect 1073 451 1085 454
rect 1027 439 1085 451
rect 259 402 317 414
rect 259 368 271 402
rect 305 368 317 402
rect 259 356 317 368
rect 547 402 605 414
rect 547 368 559 402
rect 593 368 605 402
rect 547 356 605 368
rect 835 402 893 414
rect 835 368 847 402
rect 881 368 893 402
rect 835 356 893 368
rect 1123 402 1181 414
rect 1123 368 1135 402
rect 1169 368 1181 402
rect 1123 356 1181 368
rect 274 227 302 356
rect 562 227 590 356
rect 850 227 878 356
rect 1138 227 1166 356
rect 259 215 317 227
rect 259 181 271 215
rect 305 181 317 215
rect 259 169 317 181
rect 547 215 605 227
rect 547 181 559 215
rect 593 181 605 215
rect 547 169 605 181
rect 835 215 893 227
rect 835 181 847 215
rect 881 181 893 215
rect 835 169 893 181
rect 1123 215 1181 227
rect 1123 181 1135 215
rect 1169 181 1181 215
rect 1123 169 1181 181
rect 1234 146 1262 454
rect 163 134 221 146
rect 163 100 175 134
rect 209 131 221 134
rect 1219 134 1277 146
rect 1219 131 1231 134
rect 209 103 1231 131
rect 209 100 221 103
rect 163 88 221 100
rect 1219 100 1231 103
rect 1265 100 1277 134
rect 1219 88 1277 100
rect 0 17 1440 48
rect 0 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1440 17
rect 0 -48 1440 -17
<< labels >>
rlabel metal1 0 618 1440 714 0 VPWR
port 5 se
rlabel metal1 0 618 1440 714 0 VPWR
port 5 se
rlabel metal1 0 -48 1440 48 0 VGND
port 4 se
rlabel metal1 0 -48 1440 48 0 VGND
port 4 se
rlabel metal1 163 88 221 103 0 Y
port 6 se
rlabel metal1 1219 88 1277 103 0 Y
port 6 se
rlabel metal1 163 103 1277 131 0 Y
port 6 se
rlabel metal1 163 131 221 146 0 Y
port 6 se
rlabel metal1 1219 131 1277 146 0 Y
port 6 se
rlabel metal1 1027 439 1085 454 0 Y
port 6 se
rlabel metal1 1234 146 1262 454 0 Y
port 6 se
rlabel metal1 1027 454 1262 482 0 Y
port 6 se
rlabel metal1 1027 482 1085 497 0 Y
port 6 se
rlabel metal1 259 169 317 227 0 B
port 1 se
rlabel metal1 274 227 302 356 0 B
port 1 se
rlabel metal1 259 356 317 414 0 B
port 1 se
rlabel metal1 547 169 605 227 0 A
port 0 se
rlabel metal1 562 227 590 356 0 A
port 0 se
rlabel metal1 547 356 605 414 0 A
port 0 se
rlabel metal1 1123 169 1181 227 0 D
port 3 se
rlabel metal1 1138 227 1166 356 0 D
port 3 se
rlabel metal1 1123 356 1181 414 0 D
port 3 se
rlabel metal1 835 169 893 227 0 C
port 2 se
rlabel metal1 850 227 878 356 0 C
port 2 se
rlabel metal1 835 356 893 414 0 C
port 2 se
rlabel locali 0 -17 1440 17 4 VGND
port 4 se ground default abutment
rlabel locali 31 17 1409 48 4 VGND
port 4 se ground default abutment
rlabel locali 0 649 1440 683 4 VPWR
port 5 se power default abutment
rlabel locali 31 618 1409 649 4 VGND
port 4 se power default abutment
<< properties >>
string FIXED_BBOX 0 0 1440 666
<< end >>
