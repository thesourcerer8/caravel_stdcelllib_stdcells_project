VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.330 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 1.295 1.780 1.585 2.070 ;
        RECT 5.615 1.995 5.905 2.070 ;
        RECT 4.250 1.855 5.905 1.995 ;
        RECT 1.370 1.135 1.510 1.780 ;
        RECT 4.250 1.135 4.390 1.855 ;
        RECT 5.615 1.780 5.905 1.855 ;
        RECT 1.295 1.060 1.585 1.135 ;
        RECT 4.175 1.060 4.465 1.135 ;
        RECT 1.295 0.920 4.465 1.060 ;
        RECT 1.295 0.845 1.585 0.920 ;
        RECT 4.175 0.845 4.465 0.920 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met1 ;
        RECT 2.810 2.270 8.710 2.410 ;
        RECT 2.810 2.070 2.950 2.270 ;
        RECT 8.570 2.070 8.710 2.270 ;
        RECT 2.735 1.780 3.025 2.070 ;
        RECT 8.495 1.780 8.785 2.070 ;
        RECT 8.570 1.135 8.710 1.780 ;
        RECT 8.495 0.845 8.785 1.135 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA 1.124200 ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.080 0.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 10.080 3.570 ;
        RECT 1.775 2.735 2.065 3.090 ;
        RECT 7.535 2.735 7.825 3.090 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA 1.083600 ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.245 10.080 3.415 ;
        RECT 0.155 3.215 9.925 3.245 ;
        RECT 0.155 3.090 7.345 3.215 ;
        RECT 8.015 3.090 9.925 3.215 ;
        RECT 1.755 2.715 2.085 3.090 ;
      LAYER mcon ;
        RECT 1.835 3.245 2.005 3.415 ;
        RECT 1.835 2.795 2.005 2.965 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA 1.661650 ;
    PORT
      LAYER met1 ;
        RECT 4.655 2.600 4.945 2.890 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT 0.000 1.790 10.080 3.330 ;
      LAYER li1 ;
        RECT 4.635 2.580 4.965 2.910 ;
        RECT 7.515 2.715 7.845 3.045 ;
        RECT 0.555 2.175 0.885 2.505 ;
        RECT 5.135 2.410 5.445 2.505 ;
        RECT 5.115 2.175 5.445 2.410 ;
        RECT 8.955 2.260 9.285 2.505 ;
        RECT 8.975 2.175 9.285 2.260 ;
        RECT 1.275 1.760 1.605 2.090 ;
        RECT 2.715 1.760 3.045 2.090 ;
        RECT 4.155 2.010 4.485 2.090 ;
        RECT 4.155 1.840 4.885 2.010 ;
        RECT 4.155 1.760 4.485 1.840 ;
        RECT 2.795 1.155 2.965 1.760 ;
        RECT 1.275 0.825 1.605 1.155 ;
        RECT 2.715 0.825 3.045 1.155 ;
        RECT 4.155 0.825 4.485 1.155 ;
        RECT 0.555 0.420 0.885 0.750 ;
        RECT 1.775 0.655 2.085 0.750 ;
        RECT 1.755 0.420 2.085 0.655 ;
        RECT 4.715 0.500 4.885 1.840 ;
        RECT 5.195 0.750 5.365 2.175 ;
        RECT 5.615 2.005 5.925 2.090 ;
        RECT 5.595 1.760 5.925 2.005 ;
        RECT 7.035 1.760 7.365 2.090 ;
        RECT 8.475 1.760 8.805 2.090 ;
        RECT 5.595 0.920 5.925 1.155 ;
        RECT 5.615 0.825 5.925 0.920 ;
        RECT 7.035 0.825 7.365 1.155 ;
        RECT 8.475 0.920 8.805 1.155 ;
        RECT 8.475 0.825 8.785 0.920 ;
        RECT 5.115 0.420 5.445 0.750 ;
        RECT 7.535 0.655 7.845 0.750 ;
        RECT 7.515 0.420 7.845 0.655 ;
        RECT 8.955 0.420 9.285 0.750 ;
        RECT 1.835 0.240 2.005 0.420 ;
        RECT 7.595 0.240 7.765 0.420 ;
        RECT 0.155 0.085 9.925 0.240 ;
        RECT 0.000 -0.085 10.080 0.085 ;
      LAYER mcon ;
        RECT 4.715 2.660 4.885 2.830 ;
        RECT 7.595 2.795 7.765 2.965 ;
        RECT 0.635 2.255 0.805 2.425 ;
        RECT 9.035 2.255 9.205 2.425 ;
        RECT 1.355 1.840 1.525 2.010 ;
        RECT 2.795 1.840 2.965 2.010 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 4.235 0.905 4.405 1.075 ;
        RECT 0.635 0.500 0.805 0.670 ;
        RECT 5.675 1.840 5.845 2.010 ;
        RECT 7.115 1.840 7.285 2.010 ;
        RECT 8.555 1.840 8.725 2.010 ;
        RECT 5.675 0.905 5.845 1.075 ;
        RECT 7.115 0.905 7.285 1.075 ;
        RECT 8.555 0.905 8.725 1.075 ;
        RECT 9.035 0.500 9.205 0.670 ;
        RECT 7.595 -0.085 7.765 0.085 ;
      LAYER met1 ;
        RECT 0.575 2.195 0.865 2.485 ;
        RECT 8.975 2.195 9.265 2.485 ;
        RECT 0.650 0.730 0.790 2.195 ;
        RECT 7.055 1.780 7.345 2.070 ;
        RECT 7.130 1.135 7.270 1.780 ;
        RECT 5.615 0.845 5.905 1.135 ;
        RECT 7.055 0.845 7.345 1.135 ;
        RECT 0.575 0.655 0.865 0.730 ;
        RECT 4.655 0.655 4.945 0.730 ;
        RECT 5.690 0.655 5.830 0.845 ;
        RECT 0.575 0.515 5.830 0.655 ;
        RECT 7.130 0.655 7.270 0.845 ;
        RECT 9.050 0.730 9.190 2.195 ;
        RECT 8.975 0.655 9.265 0.730 ;
        RECT 7.130 0.515 9.265 0.655 ;
        RECT 0.575 0.440 0.865 0.515 ;
        RECT 4.655 0.440 4.945 0.515 ;
        RECT 8.975 0.440 9.265 0.515 ;
  END
END XOR2X1
END LIBRARY

