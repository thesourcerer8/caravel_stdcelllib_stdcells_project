magic
tech sky130A
timestamp 1621277831
<< end >>
