VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MUX2X1
  CLASS CORE ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 3.330 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.090 8.640 3.570 ;
        RECT 1.780 3.010 2.070 3.090 ;
        RECT 1.780 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.070 3.010 ;
        RECT 1.780 2.780 2.070 2.840 ;
        RECT 7.540 3.010 7.830 3.090 ;
        RECT 7.540 2.840 7.600 3.010 ;
        RECT 7.770 2.840 7.830 3.010 ;
        RECT 7.540 2.780 7.830 2.840 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.780 0.490 2.070 0.550 ;
        RECT 1.780 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.070 0.490 ;
        RECT 1.780 0.240 2.070 0.320 ;
        RECT 7.540 0.490 7.830 0.550 ;
        RECT 7.540 0.320 7.600 0.490 ;
        RECT 7.770 0.320 7.830 0.490 ;
        RECT 7.540 0.240 7.830 0.320 ;
        RECT 0.000 -0.240 8.640 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.140 2.200 5.430 2.490 ;
        RECT 5.210 1.540 5.350 2.200 ;
        RECT 5.140 1.250 5.430 1.540 ;
    END
  END Y
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.620 2.000 5.910 2.070 ;
        RECT 5.620 1.860 6.310 2.000 ;
        RECT 5.620 1.780 5.910 1.860 ;
        RECT 1.300 1.060 1.590 1.140 ;
        RECT 4.180 1.060 4.470 1.140 ;
        RECT 1.300 0.920 4.470 1.060 ;
        RECT 1.300 0.850 1.590 0.920 ;
        RECT 4.180 0.850 4.470 0.920 ;
        RECT 4.250 0.660 4.390 0.850 ;
        RECT 6.170 0.660 6.310 1.860 ;
        RECT 4.250 0.520 6.310 0.660 ;
    END
  END S
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.740 1.250 3.030 1.540 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.060 1.780 7.350 2.070 ;
        RECT 7.130 1.140 7.270 1.780 ;
        RECT 7.060 0.850 7.350 1.140 ;
    END
  END B
  OBS
      LAYER li1 ;
        RECT 1.760 3.010 2.090 3.090 ;
        RECT 1.760 2.840 1.840 3.010 ;
        RECT 2.010 2.840 2.090 3.010 ;
        RECT 1.760 2.760 2.090 2.840 ;
        RECT 7.520 3.010 7.850 3.090 ;
        RECT 7.520 2.840 7.600 3.010 ;
        RECT 7.770 2.840 7.850 3.010 ;
        RECT 7.520 2.760 7.850 2.840 ;
        RECT 0.560 2.430 0.890 2.510 ;
        RECT 0.560 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.890 2.430 ;
        RECT 0.560 2.180 0.890 2.260 ;
        RECT 5.120 2.430 5.450 2.510 ;
        RECT 5.120 2.260 5.200 2.430 ;
        RECT 5.370 2.260 5.450 2.430 ;
        RECT 5.120 2.180 5.450 2.260 ;
        RECT 1.280 2.010 1.610 2.090 ;
        RECT 1.280 1.840 1.360 2.010 ;
        RECT 1.530 1.840 1.610 2.010 ;
        RECT 1.280 1.760 1.610 1.840 ;
        RECT 2.720 2.010 3.050 2.090 ;
        RECT 2.720 1.840 2.800 2.010 ;
        RECT 2.970 1.840 3.050 2.010 ;
        RECT 2.720 1.760 3.050 1.840 ;
        RECT 4.160 2.010 4.490 2.090 ;
        RECT 5.620 2.010 5.930 2.090 ;
        RECT 4.160 1.840 4.240 2.010 ;
        RECT 4.410 1.840 4.490 2.010 ;
        RECT 4.160 1.760 4.490 1.840 ;
        RECT 5.600 1.840 5.680 2.010 ;
        RECT 5.850 1.840 5.930 2.010 ;
        RECT 5.600 1.760 5.930 1.840 ;
        RECT 7.040 2.010 7.370 2.090 ;
        RECT 7.040 1.840 7.120 2.010 ;
        RECT 7.290 1.840 7.370 2.010 ;
        RECT 7.040 1.760 7.370 1.840 ;
        RECT 1.360 1.160 1.530 1.760 ;
        RECT 2.800 1.480 2.970 1.760 ;
        RECT 2.800 1.160 2.970 1.310 ;
        RECT 1.280 1.080 1.610 1.160 ;
        RECT 1.280 0.910 1.360 1.080 ;
        RECT 1.530 0.910 1.610 1.080 ;
        RECT 1.280 0.830 1.610 0.910 ;
        RECT 2.720 1.080 3.050 1.160 ;
        RECT 2.720 0.910 2.800 1.080 ;
        RECT 2.970 0.910 3.050 1.080 ;
        RECT 2.720 0.830 3.050 0.910 ;
        RECT 4.160 1.080 4.490 1.160 ;
        RECT 4.160 0.910 4.240 1.080 ;
        RECT 4.410 0.910 4.490 1.080 ;
        RECT 4.160 0.830 4.490 0.910 ;
        RECT 5.200 0.750 5.370 1.310 ;
        RECT 5.600 1.080 5.930 1.160 ;
        RECT 5.600 0.920 5.680 1.080 ;
        RECT 5.620 0.910 5.680 0.920 ;
        RECT 5.850 0.910 5.930 1.080 ;
        RECT 5.620 0.830 5.930 0.910 ;
        RECT 7.040 1.080 7.370 1.160 ;
        RECT 7.040 0.910 7.120 1.080 ;
        RECT 7.290 0.910 7.370 1.080 ;
        RECT 7.040 0.830 7.370 0.910 ;
        RECT 0.560 0.670 0.890 0.750 ;
        RECT 0.560 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.890 0.670 ;
        RECT 5.120 0.670 5.450 0.750 ;
        RECT 0.560 0.420 0.890 0.500 ;
        RECT 1.760 0.490 2.090 0.570 ;
        RECT 1.760 0.320 1.840 0.490 ;
        RECT 2.010 0.320 2.090 0.490 ;
        RECT 5.120 0.500 5.200 0.670 ;
        RECT 5.370 0.500 5.450 0.670 ;
        RECT 5.120 0.420 5.450 0.500 ;
        RECT 7.520 0.490 7.850 0.570 ;
        RECT 1.760 0.240 2.090 0.320 ;
        RECT 7.520 0.320 7.600 0.490 ;
        RECT 7.770 0.320 7.850 0.490 ;
        RECT 7.520 0.240 7.850 0.320 ;
      LAYER met1 ;
        RECT 0.580 2.430 0.870 2.490 ;
        RECT 0.580 2.260 0.640 2.430 ;
        RECT 0.810 2.260 0.870 2.430 ;
        RECT 0.580 2.200 0.870 2.260 ;
        RECT 0.650 2.000 0.790 2.200 ;
        RECT 4.180 2.010 4.470 2.070 ;
        RECT 4.180 2.000 4.240 2.010 ;
        RECT 0.650 1.860 4.240 2.000 ;
        RECT 0.650 0.730 0.790 1.860 ;
        RECT 4.180 1.840 4.240 1.860 ;
        RECT 4.410 2.000 4.470 2.010 ;
        RECT 4.410 1.860 4.870 2.000 ;
        RECT 4.410 1.840 4.470 1.860 ;
        RECT 4.180 1.780 4.470 1.840 ;
        RECT 4.730 1.060 4.870 1.860 ;
        RECT 5.620 1.080 5.910 1.140 ;
        RECT 5.620 1.060 5.680 1.080 ;
        RECT 4.730 0.920 5.680 1.060 ;
        RECT 5.620 0.910 5.680 0.920 ;
        RECT 5.850 0.910 5.910 1.080 ;
        RECT 5.620 0.850 5.910 0.910 ;
        RECT 0.580 0.670 0.870 0.730 ;
        RECT 0.580 0.500 0.640 0.670 ;
        RECT 0.810 0.500 0.870 0.670 ;
        RECT 0.580 0.440 0.870 0.500 ;
  END
END MUX2X1
END LIBRARY

